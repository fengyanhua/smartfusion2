`timescale 1 ns/100 ps
// Version: 
// File used only for Simulation


module sdf_IOPAD_TRI(
       PAD,
       D,
       E
    );
output PAD;
input  D;
input  E;

    wire NET_OIN_VDD, NET_EIN_VDD;
    
    IOPAD_TRI_VDDI U_VCCI (.OIN_VDD(NET_OIN_VDD), .EIN_VDD(NET_EIN_VDD)
        , .PAD_P(PAD));
    IOPAD_VDD U_VCCA (.OIN_P(D), .EIN_P(E), .IOUT_VDD(), .OIN_VDD(
        NET_OIN_VDD), .EIN_VDD(NET_EIN_VDD), .IOUT_IN());
    
endmodule


module sdf_IOPAD_IN(
       PAD,
       Y
    );
input  PAD;
output Y;

    wire NET_IOUT_VDD, NET_IOUT_IN, ADLIB_GND;
    wire GND_power_net1;
    assign ADLIB_GND = GND_power_net1;
    
    IOPAD_IN_VDDI U_VCCI (.PAD_P(PAD), .IOUT_VDD(NET_IOUT_VDD));
    IOPAD_DELAY U_DELAY (.IOUT_IN(NET_IOUT_IN), .IOUT_P(Y));
    IOPAD_VDD U_VCCA (.OIN_P(ADLIB_GND), .EIN_P(ADLIB_GND), .IOUT_VDD(
        NET_IOUT_VDD), .OIN_VDD(), .EIN_VDD(), .IOUT_IN(NET_IOUT_IN));
    GND GND_power_inst1 (.Y(GND_power_net1));
    
endmodule


module hello_regs(
       GPIO_IN,
       GPIO_OUT_1,
       MMUART_0_RXD,
       MMUART_0_TXD,
       MSS_RESET_N_M2F
    );
input  [7:0] GPIO_IN;
output [7:0] GPIO_OUT_1;
input  MMUART_0_RXD;
output MMUART_0_TXD;
output MSS_RESET_N_M2F;

    wire \CoreAPB3_0_APBmslave5_PADDR[0] , 
        \CoreAPB3_0_APBmslave5_PADDR[1] , 
        \CoreAPB3_0_APBmslave5_PADDR[2] , 
        \CoreAPB3_0_APBmslave5_PADDR[3] , 
        \CoreAPB3_0_APBmslave5_PADDR[4] , 
        \CoreAPB3_0_APBmslave5_PADDR[5] , 
        \CoreAPB3_0_APBmslave5_PADDR[6] , 
        \CoreAPB3_0_APBmslave5_PADDR[7] , 
        \CoreAPB3_0_APBmslave5_PADDR[8] , 
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PADDR[16] , 
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PADDR[17] , 
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PADDR[18] , 
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PADDR[19] , 
        CoreAPB3_0_APBmslave5_PWRITE, CoreAPB3_0_APBmslave5_PENABLE, 
        hello_regs_MSS_0_FIC_0_APB_MASTER_PSELx, 
        \CoreAPB3_0_APBmslave5_PWDATA[0] , 
        \CoreAPB3_0_APBmslave5_PWDATA[1] , 
        \CoreAPB3_0_APBmslave5_PWDATA[2] , 
        \CoreAPB3_0_APBmslave5_PWDATA[3] , 
        \CoreAPB3_0_APBmslave5_PWDATA[4] , 
        \CoreAPB3_0_APBmslave5_PWDATA[5] , 
        \CoreAPB3_0_APBmslave5_PWDATA[6] , 
        \CoreAPB3_0_APBmslave5_PWDATA[7] , 
        \CoreAPB3_0_APBmslave5_PWDATA[8] , 
        \CoreAPB3_0_APBmslave5_PWDATA[9] , 
        \CoreAPB3_0_APBmslave5_PWDATA[10] , 
        \CoreAPB3_0_APBmslave5_PWDATA[11] , 
        \CoreAPB3_0_APBmslave5_PWDATA[12] , 
        \CoreAPB3_0_APBmslave5_PWDATA[13] , 
        \CoreAPB3_0_APBmslave5_PWDATA[14] , 
        \CoreAPB3_0_APBmslave5_PWDATA[15] , 
        \CoreAPB3_0_APBmslave5_PWDATA[16] , 
        \CoreAPB3_0_APBmslave5_PWDATA[17] , 
        \CoreAPB3_0_APBmslave5_PWDATA[18] , 
        \CoreAPB3_0_APBmslave5_PWDATA[19] , 
        \CoreAPB3_0_APBmslave5_PWDATA[20] , 
        \CoreAPB3_0_APBmslave5_PWDATA[21] , 
        \CoreAPB3_0_APBmslave5_PWDATA[22] , 
        \CoreAPB3_0_APBmslave5_PWDATA[23] , 
        \CoreAPB3_0_APBmslave5_PWDATA[24] , 
        \CoreAPB3_0_APBmslave5_PWDATA[25] , 
        \CoreAPB3_0_APBmslave5_PWDATA[26] , 
        \CoreAPB3_0_APBmslave5_PWDATA[27] , 
        \CoreAPB3_0_APBmslave5_PWDATA[28] , 
        \CoreAPB3_0_APBmslave5_PWDATA[29] , 
        \CoreAPB3_0_APBmslave5_PWDATA[30] , 
        \CoreAPB3_0_APBmslave5_PWDATA[31] , 
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[0] , 
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[1] , 
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[2] , 
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[3] , 
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[4] , 
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[5] , 
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[6] , 
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[7] , 
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[8] , 
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[9] , 
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[10] , 
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[11] , 
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[12] , 
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[13] , 
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[14] , 
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[15] , 
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[16] , 
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[17] , 
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[18] , 
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[19] , 
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[20] , 
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[21] , 
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[22] , 
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[23] , 
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[24] , 
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[25] , 
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[26] , 
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[27] , 
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[28] , 
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[29] , 
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[30] , 
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[31] , 
        \CoreAPB3_0_APBmslave5_PRDATA[0] , 
        \CoreAPB3_0_APBmslave5_PRDATA[1] , 
        \CoreAPB3_0_APBmslave5_PRDATA[2] , 
        \CoreAPB3_0_APBmslave5_PRDATA[3] , 
        \CoreAPB3_0_APBmslave5_PRDATA[4] , 
        \CoreAPB3_0_APBmslave5_PRDATA[5] , 
        \CoreAPB3_0_APBmslave5_PRDATA[6] , 
        \CoreAPB3_0_APBmslave5_PRDATA[7] , 
        CoreAPB3_0_APBmslave7_PREADY, \FCCC_0/GL1_INST/U0_YNn , 
        OSC_0_RCOSC_25_50MHZ_CCC_OUT_RCOSC_25_50MHZ_CCC, FCCC_0_LOCK, 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[0] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[1] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[2] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[3] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[4] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[5] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[6] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[7] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[8] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[9] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[10] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[11] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[12] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[13] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[14] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[15] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[16] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[17] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[18] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[19] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[20] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[21] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[22] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[23] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[24] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[25] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[26] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[27] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[28] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[29] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[30] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[31] , 
        \COREAPBLSRAM_0.PRDATA4 , \COREAPBLSRAM_0.PRDATA_reg[0] , 
        \COREAPBLSRAM_0.PRDATA_reg[1] , \COREAPBLSRAM_0.PRDATA_reg[2] , 
        \COREAPBLSRAM_0.PRDATA_reg[3] , \COREAPBLSRAM_0.PRDATA_reg[4] , 
        \COREAPBLSRAM_0.PRDATA_reg[5] , \COREAPBLSRAM_0.PRDATA_reg[6] , 
        \COREAPBLSRAM_0.PRDATA_reg[7] , \COREAPBLSRAM_0.PRDATA_reg[8] , 
        \COREAPBLSRAM_0.PRDATA_reg[9] , 
        \COREAPBLSRAM_0.PRDATA_reg[10] , 
        \COREAPBLSRAM_0.PRDATA_reg[11] , 
        \COREAPBLSRAM_0.PRDATA_reg[12] , 
        \COREAPBLSRAM_0.PRDATA_reg[13] , 
        \COREAPBLSRAM_0.PRDATA_reg[14] , 
        \COREAPBLSRAM_0.PRDATA_reg[15] , 
        \COREAPBLSRAM_0.PRDATA_reg[16] , 
        \COREAPBLSRAM_0.PRDATA_reg[17] , 
        \COREAPBLSRAM_0.PRDATA_reg[18] , 
        \COREAPBLSRAM_0.PRDATA_reg[19] , 
        \COREAPBLSRAM_0.PRDATA_reg[20] , 
        \COREAPBLSRAM_0.PRDATA_reg[21] , 
        \COREAPBLSRAM_0.PRDATA_reg[22] , 
        \COREAPBLSRAM_0.PRDATA_reg[23] , 
        \COREAPBLSRAM_0.PRDATA_reg[24] , 
        \COREAPBLSRAM_0.PRDATA_reg[25] , 
        \COREAPBLSRAM_0.PRDATA_reg[26] , 
        \COREAPBLSRAM_0.PRDATA_reg[27] , 
        \COREAPBLSRAM_0.PRDATA_reg[28] , 
        \COREAPBLSRAM_0.PRDATA_reg[29] , 
        \COREAPBLSRAM_0.PRDATA_reg[30] , 
        \COREAPBLSRAM_0.PRDATA_reg[31] , N_354, N_625, N_637, N_638, 
        N_639, \GPIO_OUT_1_c[0] , \GPIO_OUT_1_c[1] , \GPIO_OUT_1_c[2] , 
        \GPIO_OUT_1_c[3] , \GPIO_OUT_1_c[4] , \GPIO_OUT_1_c[5] , 
        \GPIO_OUT_1_c[6] , \GPIO_OUT_1_c[7] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST_RNIUO3B/U0_YNn , 
        \CoreAPB3_0.u_mux_p_to_b3.PRDATA_0_iv_0_a2_3_5[1] , 
        \COREAPBLSRAM_0.PRDATA4_0_a2_0 , N_537_i_0, 
        \CoreAPB3_0/u_mux_p_to_b3/N_636 , 
        \CoreAPB3_0/u_mux_p_to_b3/PRDATA_0_iv_0_1_0[7]_net_1 , 
        \CoreAPB3_0/u_mux_p_to_b3/PRDATA_0_iv_0_0[7]_net_1 , 
        \CoreAPB3_0/u_mux_p_to_b3/PRDATA_0_iv_0_1_0[2]_net_1 , 
        \CoreAPB3_0/u_mux_p_to_b3/PRDATA_0_iv_0_0[2]_net_1 , 
        \CoreAPB3_0/u_mux_p_to_b3/PRDATA_0_iv_0_1_0[5]_net_1 , 
        \CoreAPB3_0/u_mux_p_to_b3/PRDATA_0_iv_0_0[5]_net_1 , 
        \CoreAPB3_0/u_mux_p_to_b3/PRDATA_0_iv_0_1_0[6]_net_1 , 
        \CoreAPB3_0/u_mux_p_to_b3/PRDATA_0_iv_0_0[6]_net_1 , 
        \CoreAPB3_0/u_mux_p_to_b3/PRDATA_0_iv_0_1[3]_net_1 , 
        \CoreAPB3_0/u_mux_p_to_b3/PRDATA_0_iv_0_s_0_0[3]_net_1 , 
        \CoreAPB3_0/u_mux_p_to_b3/PRDATA_0_iv_0_1[4]_net_1 , 
        \CoreAPB3_0/u_mux_p_to_b3/PRDATA_m3_i_0_net_1 , 
        \CoreAPB3_0/u_mux_p_to_b3/PRDATA_0_iv_0_a2_3_5_4[1]_net_1 , 
        \CoreAPB3_0/u_mux_p_to_b3/PRDATA_0_iv_0_a2_3_5_3[1]_net_1 , 
        \CoreAPB3_0/u_mux_p_to_b3/PRDATA_N_8_0 , 
        \CoreAPB3_0/u_mux_p_to_b3/PRDATA_0_iv_0_a2_2_0[7]_net_1 , 
        \CoreAPB3_0/u_mux_p_to_b3/PRDATA_0_iv_0_a2_2_0[5]_net_1 , 
        \CoreAPB3_0/u_mux_p_to_b3/PRDATA_0_iv_0_a2_2_0[2]_net_1 , 
        \CoreAPB3_0/u_mux_p_to_b3/PRDATA_0_iv_0_a2_2_0[6]_net_1 , 
        \CoreAPB3_0/u_mux_p_to_b3/N_584 , 
        \CoreAPB3_0/u_mux_p_to_b3/N_585 , 
        \CoreAPB3_0/u_mux_p_to_b3/PRDATA_0_iv_0_0[0]_net_1 , 
        \CoreAPB3_0/u_mux_p_to_b3/PRDATA_0_iv_0_0[1]_net_1 , 
        \hello_regs_MSS_0/FPGA_RESET_N , 
        \hello_regs_MSS_0/MSS_ADLIB_INST_MMUART0_TXD_USBC_DIR_MGPIO27B_OUT , 
        \hello_regs_MSS_0/MSS_ADLIB_INST_MMUART0_TXD_USBC_DIR_MGPIO27B_OE , 
        \hello_regs_MSS_0/MMUART_0_RXD_PAD_Y , VCC, GND, 
        \FCCC_0/GL1_net , \reg_apb_wrp_0/rd_enable , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_121_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_25_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_9_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_80_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_27_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_11_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_81_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_57_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_112_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_104_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_16_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_88_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_97_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_72_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_7_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_124_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_28_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_12_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_13_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_82_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_58_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_113_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_105_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_17_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_89_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_98_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_73_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_5_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_126_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_30_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_14_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_2_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_123_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_83_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_59_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_114_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_106_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_18_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_90_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_99_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_74_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_64_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_48_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_32_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_43_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_4_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_125_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_29_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_56_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_115_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_107_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_19_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_91_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_96_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_75_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_66_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_50_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_34_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_41_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_6_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_127_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_31_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_15_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_116_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_108_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_20_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_92_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_101_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_76_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_68_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_52_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_36_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_47_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_65_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_49_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_33_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_40_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_84_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_109_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_21_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_93_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_102_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_77_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_69_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_54_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_38_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_45_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_67_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_51_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_35_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_42_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_85_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_61_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_22_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_94_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_103_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_78_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_70_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_3_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_120_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_24_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_8_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_53_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_37_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_44_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_86_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_62_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_117_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_95_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_100_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_79_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_71_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_1_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_122_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_26_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_10_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_55_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_39_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_46_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_87_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_63_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_118_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_110_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_60_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_119_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_111_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_23_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/N_7_i_0 , 
        \reg_apb_wrp_0/reg16x8_0/N_13_i_0 , 
        \reg_apb_wrp_0/reg16x8_0/N_15_i_0 , 
        \reg_apb_wrp_0/reg16x8_0/N_37_i_0 , 
        \reg_apb_wrp_0/reg16x8_0/N_41_i_0 , 
        \reg_apb_wrp_0/reg16x8_0/N_82_i_0 , 
        \reg_apb_wrp_0/reg16x8_0/N_22_i_0 , 
        \reg_apb_wrp_0/reg16x8_0/N_84_i_0 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_23_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_247_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_12_rs[7] , 
        \reg_apb_wrp_0/reg16x8_0/mem_12_[7]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_247_i , 
        \reg_apb_wrp_0/reg16x8_0/mem_12__1_sqmuxa , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_111_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_215_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_13_rs[7] , 
        \reg_apb_wrp_0/reg16x8_0/mem_13_[7]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_215_i , 
        \reg_apb_wrp_0/reg16x8_0/mem_13__1_sqmuxa , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_119_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_223_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_14_rs[7] , 
        \reg_apb_wrp_0/reg16x8_0/mem_14_[7]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_223_i , 
        \reg_apb_wrp_0/reg16x8_0/mem_14__1_sqmuxa , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_60_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_254_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_15_rs[7] , 
        \reg_apb_wrp_0/reg16x8_0/mem_15_[7]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_254_i , 
        \reg_apb_wrp_0/reg16x8_0/mem_15__1_sqmuxa , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_110_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_214_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_13_rs[6] , 
        \reg_apb_wrp_0/reg16x8_0/mem_13_[6]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_214_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_118_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_222_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_14_rs[6] , 
        \reg_apb_wrp_0/reg16x8_0/mem_14_[6]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_222_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_63_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_253_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_15_rs[6] , 
        \reg_apb_wrp_0/reg16x8_0/mem_15_[6]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_253_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_87_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_151_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_0_rs[7] , 
        \reg_apb_wrp_0/reg16x8_0/mem_0_[7]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_151_i , 
        \reg_apb_wrp_0/reg16x8_0/mem_0__1_sqmuxa , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_46_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_159_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_1_rs[7] , 
        \reg_apb_wrp_0/reg16x8_0/mem_1_[7]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_159_i , 
        \reg_apb_wrp_0/reg16x8_0/mem_1__1_sqmuxa , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_39_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_167_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_2_rs[7] , 
        \reg_apb_wrp_0/reg16x8_0/mem_2_[7]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_167_i , 
        \reg_apb_wrp_0/reg16x8_0/mem_2__1_sqmuxa , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_55_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_135_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_3_rs[7] , 
        \reg_apb_wrp_0/reg16x8_0/mem_3_[7]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_135_i , 
        \reg_apb_wrp_0/reg16x8_0/mem_3__1_sqmuxa , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_10_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_185_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_4_rs[7] , 
        \reg_apb_wrp_0/reg16x8_0/mem_4_[7]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_185_i , 
        \reg_apb_wrp_0/reg16x8_0/mem_4__1_sqmuxa , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_26_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_201_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_5_rs[7] , 
        \reg_apb_wrp_0/reg16x8_0/mem_5_[7]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_201_i , 
        \reg_apb_wrp_0/reg16x8_0/mem_5__1_sqmuxa , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_122_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_177_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_6_rs[7] , 
        \reg_apb_wrp_0/reg16x8_0/mem_6_[7]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_177_i , 
        \reg_apb_wrp_0/reg16x8_0/mem_6__1_sqmuxa , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_1_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_233_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_7_rs[7] , 
        \reg_apb_wrp_0/reg16x8_0/mem_7_[7]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_233_i , 
        \reg_apb_wrp_0/reg16x8_0/mem_7__1_sqmuxa , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_71_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_188_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_8_rs[7] , 
        \reg_apb_wrp_0/reg16x8_0/mem_8_[7]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_188_i , 
        \reg_apb_wrp_0/reg16x8_0/mem_8__1_sqmuxa , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_79_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_204_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_9_rs[7] , 
        \reg_apb_wrp_0/reg16x8_0/mem_9_[7]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_204_i , 
        \reg_apb_wrp_0/reg16x8_0/mem_9__1_sqmuxa , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_100_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_180_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_10_rs[7] , 
        \reg_apb_wrp_0/reg16x8_0/mem_10_[7]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_180_i , 
        \reg_apb_wrp_0/reg16x8_0/mem_10__1_sqmuxa , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_95_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_236_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_11_rs[7] , 
        \reg_apb_wrp_0/reg16x8_0/mem_11_[7]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_236_i , 
        \reg_apb_wrp_0/reg16x8_0/mem_11__1_sqmuxa , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_117_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_221_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_14_rs[5] , 
        \reg_apb_wrp_0/reg16x8_0/mem_14_[5]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_221_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_62_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_252_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_15_rs[5] , 
        \reg_apb_wrp_0/reg16x8_0/mem_15_[5]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_252_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_86_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_150_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_0_rs[6] , 
        \reg_apb_wrp_0/reg16x8_0/mem_0_[6]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_150_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_44_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_158_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_1_rs[6] , 
        \reg_apb_wrp_0/reg16x8_0/mem_1_[6]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_158_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_37_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_166_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_2_rs[6] , 
        \reg_apb_wrp_0/reg16x8_0/mem_2_[6]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_166_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_53_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_134_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_3_rs[6] , 
        \reg_apb_wrp_0/reg16x8_0/mem_3_[6]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_134_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_8_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_143_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_4_rs[6] , 
        \reg_apb_wrp_0/reg16x8_0/mem_4_[6]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_143_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_24_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_199_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_5_rs[6] , 
        \reg_apb_wrp_0/reg16x8_0/mem_5_[6]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_199_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_120_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_175_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_6_rs[6] , 
        \reg_apb_wrp_0/reg16x8_0/mem_6_[6]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_175_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_3_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_231_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_7_rs[6] , 
        \reg_apb_wrp_0/reg16x8_0/mem_7_[6]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_231_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_70_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_186_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_8_rs[6] , 
        \reg_apb_wrp_0/reg16x8_0/mem_8_[6]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_186_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_78_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_202_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_9_rs[6] , 
        \reg_apb_wrp_0/reg16x8_0/mem_9_[6]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_202_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_103_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_178_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_10_rs[6] , 
        \reg_apb_wrp_0/reg16x8_0/mem_10_[6]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_178_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_94_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_234_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_11_rs[6] , 
        \reg_apb_wrp_0/reg16x8_0/mem_11_[6]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_234_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_22_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_246_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_12_rs[6] , 
        \reg_apb_wrp_0/reg16x8_0/mem_12_[6]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_246_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_61_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_255_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_15_rs[4] , 
        \reg_apb_wrp_0/reg16x8_0/mem_15_[4]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_255_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_85_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_149_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_0_rs[5] , 
        \reg_apb_wrp_0/reg16x8_0/mem_0_[5]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_149_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_42_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_157_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_1_rs[5] , 
        \reg_apb_wrp_0/reg16x8_0/mem_1_[5]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_157_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_35_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_165_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_2_rs[5] , 
        \reg_apb_wrp_0/reg16x8_0/mem_2_[5]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_165_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_51_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_133_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_3_rs[5] , 
        \reg_apb_wrp_0/reg16x8_0/mem_3_[5]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_133_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_67_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_141_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_4_rs[5] , 
        \reg_apb_wrp_0/reg16x8_0/mem_4_[5]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_141_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_45_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_197_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_5_rs[5] , 
        \reg_apb_wrp_0/reg16x8_0/mem_5_[5]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_197_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_38_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_173_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_6_rs[5] , 
        \reg_apb_wrp_0/reg16x8_0/mem_6_[5]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_173_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_54_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_229_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_7_rs[5] , 
        \reg_apb_wrp_0/reg16x8_0/mem_7_[5]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_229_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_69_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_184_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_8_rs[5] , 
        \reg_apb_wrp_0/reg16x8_0/mem_8_[5]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_184_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_77_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_200_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_9_rs[5] , 
        \reg_apb_wrp_0/reg16x8_0/mem_9_[5]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_200_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_102_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_176_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_10_rs[5] , 
        \reg_apb_wrp_0/reg16x8_0/mem_10_[5]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_176_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_93_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_232_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_11_rs[5] , 
        \reg_apb_wrp_0/reg16x8_0/mem_11_[5]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_232_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_21_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_245_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_12_rs[5] , 
        \reg_apb_wrp_0/reg16x8_0/mem_12_[5]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_245_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_109_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_213_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_13_rs[5] , 
        \reg_apb_wrp_0/reg16x8_0/mem_13_[5]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_213_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_84_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_148_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_0_rs[4] , 
        \reg_apb_wrp_0/reg16x8_0/mem_0_[4]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_148_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_40_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_156_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_1_rs[4] , 
        \reg_apb_wrp_0/reg16x8_0/mem_1_[4]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_156_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_33_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_164_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_2_rs[4] , 
        \reg_apb_wrp_0/reg16x8_0/mem_2_[4]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_164_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_49_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_132_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_3_rs[4] , 
        \reg_apb_wrp_0/reg16x8_0/mem_3_[4]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_132_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_65_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_140_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_4_rs[4] , 
        \reg_apb_wrp_0/reg16x8_0/mem_4_[4]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_140_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_47_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_195_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_5_rs[4] , 
        \reg_apb_wrp_0/reg16x8_0/mem_5_[4]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_195_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_36_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_171_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_6_rs[4] , 
        \reg_apb_wrp_0/reg16x8_0/mem_6_[4]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_171_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_52_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_227_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_7_rs[4] , 
        \reg_apb_wrp_0/reg16x8_0/mem_7_[4]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_227_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_68_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_142_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_8_rs[4] , 
        \reg_apb_wrp_0/reg16x8_0/mem_8_[4]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_142_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_76_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_198_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_9_rs[4] , 
        \reg_apb_wrp_0/reg16x8_0/mem_9_[4]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_198_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_101_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_174_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_10_rs[4] , 
        \reg_apb_wrp_0/reg16x8_0/mem_10_[4]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_174_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_92_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_230_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_11_rs[4] , 
        \reg_apb_wrp_0/reg16x8_0/mem_11_[4]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_230_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_20_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_244_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_12_rs[4] , 
        \reg_apb_wrp_0/reg16x8_0/mem_12_[4]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_244_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_108_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_212_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_13_rs[4] , 
        \reg_apb_wrp_0/reg16x8_0/mem_13_[4]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_212_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_116_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_220_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_14_rs[4] , 
        \reg_apb_wrp_0/reg16x8_0/mem_14_[4]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_220_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_15_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_155_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_1_rs[3] , 
        \reg_apb_wrp_0/reg16x8_0/mem_1_[3]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_155_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_31_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_163_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_2_rs[3] , 
        \reg_apb_wrp_0/reg16x8_0/mem_2_[3]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_163_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_127_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_131_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_3_rs[3] , 
        \reg_apb_wrp_0/reg16x8_0/mem_3_[3]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_131_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_6_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_139_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_4_rs[3] , 
        \reg_apb_wrp_0/reg16x8_0/mem_4_[3]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_139_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_41_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_193_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_5_rs[3] , 
        \reg_apb_wrp_0/reg16x8_0/mem_5_[3]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_193_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_34_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_169_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_6_rs[3] , 
        \reg_apb_wrp_0/reg16x8_0/mem_6_[3]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_169_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_50_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_225_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_7_rs[3] , 
        \reg_apb_wrp_0/reg16x8_0/mem_7_[3]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_225_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_66_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_241_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_8_rs[3] , 
        \reg_apb_wrp_0/reg16x8_0/mem_8_[3]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_241_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_75_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_196_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_9_rs[3] , 
        \reg_apb_wrp_0/reg16x8_0/mem_9_[3]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_196_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_96_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_172_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_10_rs[3] , 
        \reg_apb_wrp_0/reg16x8_0/mem_10_[3]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_172_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_91_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_228_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_11_rs[3] , 
        \reg_apb_wrp_0/reg16x8_0/mem_11_[3]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_228_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_19_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_243_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_12_rs[3] , 
        \reg_apb_wrp_0/reg16x8_0/mem_12_[3]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_243_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_107_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_211_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_13_rs[3] , 
        \reg_apb_wrp_0/reg16x8_0/mem_13_[3]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_211_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_115_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_219_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_14_rs[3] , 
        \reg_apb_wrp_0/reg16x8_0/mem_14_[3]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_219_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_56_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_250_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_15_rs[3] , 
        \reg_apb_wrp_0/reg16x8_0/mem_15_[3]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_250_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_29_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_162_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_2_rs[2] , 
        \reg_apb_wrp_0/reg16x8_0/mem_2_[2]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_162_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_125_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_130_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_3_rs[2] , 
        \reg_apb_wrp_0/reg16x8_0/mem_3_[2]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_130_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_4_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_138_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_4_rs[2] , 
        \reg_apb_wrp_0/reg16x8_0/mem_4_[2]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_138_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_43_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_191_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_5_rs[2] , 
        \reg_apb_wrp_0/reg16x8_0/mem_5_[2]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_191_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_32_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_207_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_6_rs[2] , 
        \reg_apb_wrp_0/reg16x8_0/mem_6_[2]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_207_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_48_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_183_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_7_rs[2] , 
        \reg_apb_wrp_0/reg16x8_0/mem_7_[2]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_183_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_64_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_239_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_8_rs[2] , 
        \reg_apb_wrp_0/reg16x8_0/mem_8_[2]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_239_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_74_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_194_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_9_rs[2] , 
        \reg_apb_wrp_0/reg16x8_0/mem_9_[2]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_194_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_99_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_170_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_10_rs[2] , 
        \reg_apb_wrp_0/reg16x8_0/mem_10_[2]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_170_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_90_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_226_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_11_rs[2] , 
        \reg_apb_wrp_0/reg16x8_0/mem_11_[2]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_226_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_18_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_242_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_12_rs[2] , 
        \reg_apb_wrp_0/reg16x8_0/mem_12_[2]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_242_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_106_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_210_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_13_rs[2] , 
        \reg_apb_wrp_0/reg16x8_0/mem_13_[2]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_210_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_114_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_218_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_14_rs[2] , 
        \reg_apb_wrp_0/reg16x8_0/mem_14_[2]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_218_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_59_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_249_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_15_rs[2] , 
        \reg_apb_wrp_0/reg16x8_0/mem_15_[2]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_249_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_83_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_146_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_0_rs[3] , 
        \reg_apb_wrp_0/reg16x8_0/mem_0_[3]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_146_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_123_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_129_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_3_rs[1] , 
        \reg_apb_wrp_0/reg16x8_0/mem_3_[1]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_129_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_2_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_137_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_4_rs[1] , 
        \reg_apb_wrp_0/reg16x8_0/mem_4_[1]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_137_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_14_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_189_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_5_rs[1] , 
        \reg_apb_wrp_0/reg16x8_0/mem_5_[1]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_189_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_30_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_205_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_6_rs[1] , 
        \reg_apb_wrp_0/reg16x8_0/mem_6_[1]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_205_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_126_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_181_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_7_rs[1] , 
        \reg_apb_wrp_0/reg16x8_0/mem_7_[1]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_181_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_5_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_237_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_8_rs[1] , 
        \reg_apb_wrp_0/reg16x8_0/mem_8_[1]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_237_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_73_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_192_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_9_rs[1] , 
        \reg_apb_wrp_0/reg16x8_0/mem_9_[1]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_192_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_98_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_168_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_10_rs[1] , 
        \reg_apb_wrp_0/reg16x8_0/mem_10_[1]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_168_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_89_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_224_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_11_rs[1] , 
        \reg_apb_wrp_0/reg16x8_0/mem_11_[1]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_224_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_17_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_240_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_12_rs[1] , 
        \reg_apb_wrp_0/reg16x8_0/mem_12_[1]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_240_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_105_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_209_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_13_rs[1] , 
        \reg_apb_wrp_0/reg16x8_0/mem_13_[1]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_209_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_113_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_217_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_14_rs[1] , 
        \reg_apb_wrp_0/reg16x8_0/mem_14_[1]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_217_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_58_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_248_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_15_rs[1] , 
        \reg_apb_wrp_0/reg16x8_0/mem_15_[1]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_248_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_82_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_145_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_0_rs[2] , 
        \reg_apb_wrp_0/reg16x8_0/mem_0_[2]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_145_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_13_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_154_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_1_rs[2] , 
        \reg_apb_wrp_0/reg16x8_0/mem_1_[2]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_154_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_136_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_4_rs[0] , 
        \reg_apb_wrp_0/reg16x8_0/mem_4_[0]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_136_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_12_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_187_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_5_rs[0] , 
        \reg_apb_wrp_0/reg16x8_0/mem_5_[0]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_187_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_28_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_203_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_6_rs[0] , 
        \reg_apb_wrp_0/reg16x8_0/mem_6_[0]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_203_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_124_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_179_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_7_rs[0] , 
        \reg_apb_wrp_0/reg16x8_0/mem_7_[0]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_179_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_7_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_235_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_8_rs[0] , 
        \reg_apb_wrp_0/reg16x8_0/mem_8_[0]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_235_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_72_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_190_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_9_rs[0] , 
        \reg_apb_wrp_0/reg16x8_0/mem_9_[0]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_190_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_97_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_206_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_10_rs[0] , 
        \reg_apb_wrp_0/reg16x8_0/mem_10_[0]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_206_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_88_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_182_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_11_rs[0] , 
        \reg_apb_wrp_0/reg16x8_0/mem_11_[0]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_182_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_16_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_238_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_12_rs[0] , 
        \reg_apb_wrp_0/reg16x8_0/mem_12_[0]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_238_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_104_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_208_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_13_rs[0] , 
        \reg_apb_wrp_0/reg16x8_0/mem_13_[0]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_208_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_112_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_216_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_14_rs[0] , 
        \reg_apb_wrp_0/reg16x8_0/mem_14_[0]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_216_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_57_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_251_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_15_rs[0] , 
        \reg_apb_wrp_0/reg16x8_0/mem_15_[0]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_251_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_81_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_144_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_0_rs[1] , 
        \reg_apb_wrp_0/reg16x8_0/mem_0_[1]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_144_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_11_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_153_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_1_rs[1] , 
        \reg_apb_wrp_0/reg16x8_0/mem_1_[1]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_153_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_27_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_161_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_2_rs[1] , 
        \reg_apb_wrp_0/reg16x8_0/mem_2_[1]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_161_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_80_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_147_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_0_rs[0] , 
        \reg_apb_wrp_0/reg16x8_0/mem_0_[0]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_147_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_9_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_152_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_1_rs[0] , 
        \reg_apb_wrp_0/reg16x8_0/mem_1_[0]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_152_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_25_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_160_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_2_rs[0] , 
        \reg_apb_wrp_0/reg16x8_0/mem_2_[0]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_160_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_121_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_128_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_3_rs[0] , 
        \reg_apb_wrp_0/reg16x8_0/mem_3_[0]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_128_i , 
        \reg_apb_wrp_0/reg16x8_0/N_655 , 
        \reg_apb_wrp_0/reg16x8_0/N_654 , 
        \reg_apb_wrp_0/reg16x8_0/N_653 , 
        \reg_apb_wrp_0/reg16x8_0/N_652 , 
        \reg_apb_wrp_0/reg16x8_0/N_651 , 
        \reg_apb_wrp_0/reg16x8_0/N_650 , 
        \reg_apb_wrp_0/reg16x8_0/N_649 , 
        \reg_apb_wrp_0/reg16x8_0/N_648 , 
        \reg_apb_wrp_0/reg16x8_0/N_647 , 
        \reg_apb_wrp_0/reg16x8_0/N_646 , 
        \reg_apb_wrp_0/reg16x8_0/N_645 , 
        \reg_apb_wrp_0/reg16x8_0/N_644 , 
        \reg_apb_wrp_0/reg16x8_0/N_643 , 
        \reg_apb_wrp_0/reg16x8_0/N_642 , 
        \reg_apb_wrp_0/reg16x8_0/N_641 , 
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_7[3]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_6[3]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_5[3]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_4[3]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_3[3]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_2[3]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_1[3]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_0[3]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_7[2]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_6[2]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_5[2]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_4[2]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_3[2]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_2[2]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_1[2]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_0[2]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_7[1]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_6[1]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_5[1]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_4[1]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_3[1]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_2[1]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_1[1]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_0[1]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_7[4]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_6[4]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_5[4]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_4[4]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_3[4]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_2[4]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_1[4]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_0[4]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_7[0]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_6[0]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_5[0]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_4[0]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_3[0]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_2[0]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_1[0]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_0[0]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_0_7[6]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_0_6[6]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_0_5[6]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_0_4[6]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_0_3[6]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_0_2[6]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_0_1[6]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_0_0[6]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_7[7]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_6[7]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_5[7]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_4[7]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_3[7]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_2[7]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_1[7]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_0[7]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_7[5]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_6[5]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_5[5]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_4[5]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_3[5]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_2[5]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_1[5]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_0[5]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_13[3]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_12[3]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_13[2]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_12[2]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_13[1]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_12[1]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_13[4]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_12[4]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_13[0]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_12[0]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_0_13[6]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_0_12[6]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_13[7]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_12[7]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_13[5]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_12[5]_net_1 , 
        \CoreGPIO_0/GPOUT_reg35 , \COREAPBLSRAM_0/PREADY_reg6_i_0 , 
        \COREAPBLSRAM_0/PREADY_reg6_0_a2_0_net_1 , 
        \COREAPBLSRAM_0/wen , ff_to_start_net, 
        \hello_regs_MSS_0/MSS_ADLIB_INST/CAN_RXBUS_F2H_SCP_net , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/CAN_TX_EBL_F2H_SCP_net , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/CAN_TXBUS_F2H_SCP_net , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/COLF_net , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/CRSF_net , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F2_DMAREADY_net[1] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F2_DMAREADY_net[0] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[15] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[14] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[13] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[12] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[11] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[10] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[9] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[8] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[7] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[6] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[5] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[4] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[3] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[2] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[1] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[0] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F2HCALIB_net , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_DMAREADY_net[1] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_DMAREADY_net[0] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[31] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[30] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[29] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[28] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[27] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[26] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[25] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[24] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[23] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[22] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[21] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[20] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[19] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[18] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[17] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[16] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[15] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[14] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[13] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[12] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[11] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[10] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[9] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[8] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[7] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[6] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[5] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[4] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[3] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[2] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[1] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[0] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_ENABLE_net , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_MASTLOCK_net , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_READY_net , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_SEL_net , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_SIZE_net[1] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_SIZE_net[0] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_TRANS1_net , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[31] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[30] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[29] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[28] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[27] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[26] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[25] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[24] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[23] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[22] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[21] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[20] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[19] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[18] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[17] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[16] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[15] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[14] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[13] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[12] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[11] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[10] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[9] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[8] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[7] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[6] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[5] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[4] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[3] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[2] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[1] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[0] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_WRITE_net , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[31] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[30] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[29] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[28] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[27] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[26] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[25] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[24] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[23] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[22] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[21] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[20] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[19] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[18] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[17] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[16] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[15] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[14] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[13] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[12] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[11] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[10] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[9] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[8] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[7] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[6] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[5] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[4] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[3] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[2] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[1] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[0] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_HM0_READY_net , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_HM0_RESP_net , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/FAB_AVALID_net , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/FAB_HOSTDISCON_net , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/FAB_IDDIG_net , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/FAB_LINESTATE_net[1] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/FAB_LINESTATE_net[0] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/FAB_M3_RESET_N_net , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/FAB_PLL_LOCK_net , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/FAB_RXACTIVE_net , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/FAB_RXERROR_net , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/FAB_RXVALID_net , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/FAB_RXVALIDH_net , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/FAB_SESSEND_net , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/FAB_TXREADY_net , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/FAB_VBUSVALID_net , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/FAB_VSTATUS_net[7] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/FAB_VSTATUS_net[6] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/FAB_VSTATUS_net[5] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/FAB_VSTATUS_net[4] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/FAB_VSTATUS_net[3] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/FAB_VSTATUS_net[2] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/FAB_VSTATUS_net[1] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/FAB_VSTATUS_net[0] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/FAB_XDATAIN_net[7] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/FAB_XDATAIN_net[6] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/FAB_XDATAIN_net[5] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/FAB_XDATAIN_net[4] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/FAB_XDATAIN_net[3] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/FAB_XDATAIN_net[2] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/FAB_XDATAIN_net[1] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/FAB_XDATAIN_net[0] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/GTX_CLKPF_net , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/I2C0_BCLK_net , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/I2C0_SCL_F2H_SCP_net , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/I2C0_SDA_F2H_SCP_net , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/I2C1_BCLK_net , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/I2C1_SCL_F2H_SCP_net , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/I2C1_SDA_F2H_SCP_net , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/MDIF_net , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/MGPIO0A_F2H_GPIN_net , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/MGPIO10A_F2H_GPIN_net , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/MGPIO11A_F2H_GPIN_net , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/MGPIO11B_F2H_GPIN_net , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/MGPIO12A_F2H_GPIN_net , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/MGPIO13A_F2H_GPIN_net , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/MGPIO14A_F2H_GPIN_net , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/MGPIO15A_F2H_GPIN_net , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/MGPIO16A_F2H_GPIN_net , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/MGPIO17B_F2H_GPIN_net , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/MGPIO18B_F2H_GPIN_net , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/MGPIO19B_F2H_GPIN_net , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/MGPIO1A_F2H_GPIN_net , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/MGPIO20B_F2H_GPIN_net , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/MGPIO21B_F2H_GPIN_net , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/MGPIO22B_F2H_GPIN_net , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/MGPIO24B_F2H_GPIN_net , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/MGPIO25B_F2H_GPIN_net , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/MGPIO26B_F2H_GPIN_net , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/MGPIO27B_F2H_GPIN_net , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/MGPIO28B_F2H_GPIN_net , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/MGPIO29B_F2H_GPIN_net , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/MGPIO2A_F2H_GPIN_net , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/MGPIO30B_F2H_GPIN_net , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/MGPIO31B_F2H_GPIN_net , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/MGPIO3A_F2H_GPIN_net , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/MGPIO4A_F2H_GPIN_net , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/MGPIO5A_F2H_GPIN_net , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/MGPIO6A_F2H_GPIN_net , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/MGPIO7A_F2H_GPIN_net , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/MGPIO8A_F2H_GPIN_net , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/MGPIO9A_F2H_GPIN_net , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/MMUART0_CTS_F2H_SCP_net , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/MMUART0_DCD_F2H_SCP_net , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/MMUART0_DSR_F2H_SCP_net , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/MMUART0_DTR_F2H_SCP_net , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/MMUART0_RI_F2H_SCP_net , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/MMUART0_RTS_F2H_SCP_net , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/MMUART0_RXD_F2H_SCP_net , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/MMUART0_SCK_F2H_SCP_net , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/MMUART0_TXD_F2H_SCP_net , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/MMUART1_CTS_F2H_SCP_net , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/MMUART1_DCD_F2H_SCP_net , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/MMUART1_DSR_F2H_SCP_net , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/MMUART1_RI_F2H_SCP_net , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/MMUART1_RTS_F2H_SCP_net , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/MMUART1_RXD_F2H_SCP_net , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/MMUART1_SCK_F2H_SCP_net , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/MMUART1_TXD_F2H_SCP_net , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[31] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[30] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[29] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[28] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[27] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[26] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[25] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[24] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[23] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[22] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[21] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[20] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[19] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[18] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[17] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[16] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[15] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[14] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[13] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[12] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[11] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[10] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[9] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[8] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[7] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[6] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[5] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[4] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[3] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[2] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[1] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[0] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PREADY_net , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PSLVERR_net , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/RCGF_net[9] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/RCGF_net[8] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/RCGF_net[7] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/RCGF_net[6] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/RCGF_net[5] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/RCGF_net[4] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/RCGF_net[3] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/RCGF_net[2] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/RCGF_net[1] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/RCGF_net[0] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/RX_CLKPF_net , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/RX_DVF_net , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/RX_ERRF_net , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/RX_EV_net , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/RXDF_net[7] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/RXDF_net[6] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/RXDF_net[5] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/RXDF_net[4] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/RXDF_net[3] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/RXDF_net[2] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/RXDF_net[1] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/RXDF_net[0] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/SLEEPHOLDREQ_net , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/SMBALERT_NI0_net , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/SMBALERT_NI1_net , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/SMBSUS_NI0_net , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/SMBSUS_NI1_net , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/SPI0_CLK_IN_net , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/SPI0_SDI_F2H_SCP_net , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/SPI0_SDO_F2H_SCP_net , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/SPI0_SS0_F2H_SCP_net , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/SPI0_SS1_F2H_SCP_net , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/SPI0_SS2_F2H_SCP_net , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/SPI0_SS3_F2H_SCP_net , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/SPI1_CLK_IN_net , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/SPI1_SDI_F2H_SCP_net , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/SPI1_SDO_F2H_SCP_net , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/SPI1_SS0_F2H_SCP_net , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/SPI1_SS1_F2H_SCP_net , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/SPI1_SS2_F2H_SCP_net , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/SPI1_SS3_F2H_SCP_net , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/TX_CLKPF_net , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/USER_MSS_GPIO_RESET_N_net , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/USER_MSS_RESET_N_net , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/XCLK_FAB_net , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/CLK_BASE_net , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/CLK_MDDR_APB_net , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[31] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[30] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[29] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[28] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[27] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[26] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[25] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[24] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[23] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[22] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[21] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[20] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[19] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[18] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[17] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[16] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[15] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[14] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[13] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[12] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[11] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[10] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[9] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[8] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[7] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[6] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[5] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[4] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[3] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[2] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[1] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[0] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_ARBURST_HTRANS1_net[1] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_ARBURST_HTRANS1_net[0] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_ARID_HSEL1_net[3] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_ARID_HSEL1_net[2] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_ARID_HSEL1_net[1] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_ARID_HSEL1_net[0] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_ARLEN_HBURST1_net[3] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_ARLEN_HBURST1_net[2] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_ARLEN_HBURST1_net[1] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_ARLEN_HBURST1_net[0] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_ARLOCK_HMASTLOCK1_net[1] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_ARLOCK_HMASTLOCK1_net[0] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_ARSIZE_HSIZE1_net[1] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_ARSIZE_HSIZE1_net[0] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_ARVALID_HWRITE1_net , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[31] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[30] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[29] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[28] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[27] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[26] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[25] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[24] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[23] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[22] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[21] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[20] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[19] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[18] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[17] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[16] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[15] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[14] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[13] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[12] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[11] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[10] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[9] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[8] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[7] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[6] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[5] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[4] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[3] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[2] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[1] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[0] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_AWBURST_HTRANS0_net[1] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_AWBURST_HTRANS0_net[0] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_AWID_HSEL0_net[3] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_AWID_HSEL0_net[2] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_AWID_HSEL0_net[1] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_AWID_HSEL0_net[0] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_AWLEN_HBURST0_net[3] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_AWLEN_HBURST0_net[2] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_AWLEN_HBURST0_net[1] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_AWLEN_HBURST0_net[0] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_AWLOCK_HMASTLOCK0_net[1] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_AWLOCK_HMASTLOCK0_net[0] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_AWSIZE_HSIZE0_net[1] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_AWSIZE_HSIZE0_net[0] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_AWVALID_HWRITE0_net , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_BREADY_net , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_RMW_AXI_net , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_RREADY_net , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[63] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[62] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[61] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[60] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[59] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[58] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[57] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[56] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[55] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[54] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[53] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[52] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[51] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[50] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[49] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[48] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[47] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[46] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[45] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[44] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[43] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[42] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[41] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[40] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[39] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[38] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[37] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[36] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[35] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[34] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[33] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[32] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[31] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[30] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[29] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[28] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[27] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[26] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[25] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[24] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[23] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[22] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[21] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[20] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[19] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[18] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[17] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[16] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[15] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[14] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[13] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[12] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[11] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[10] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[9] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[8] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[7] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[6] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[5] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[4] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[3] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[2] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[1] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[0] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WID_HREADY01_net[3] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WID_HREADY01_net[2] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WID_HREADY01_net[1] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WID_HREADY01_net[0] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WLAST_net , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WSTRB_net[7] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WSTRB_net[6] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WSTRB_net[5] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WSTRB_net[4] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WSTRB_net[3] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WSTRB_net[2] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WSTRB_net[1] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WSTRB_net[0] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WVALID_net , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/FPGA_MDDR_ARESET_N_net , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PADDR_net[10] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PADDR_net[9] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PADDR_net[8] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PADDR_net[7] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PADDR_net[6] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PADDR_net[5] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PADDR_net[4] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PADDR_net[3] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PADDR_net[2] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PENABLE_net , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PSEL_net , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[15] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[14] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[13] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[12] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[11] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[10] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[9] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[8] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[7] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[6] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[5] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[4] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[3] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[2] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[1] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[0] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWRITE_net , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/PRESET_N_net , 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/A_CLK_net , 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/A_DOUT_CLK_net , 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/A_ARST_N_net , 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/A_DOUT_EN_net , 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/A_BLK_net[2] , 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/A_BLK_net[1] , 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/A_BLK_net[0] , 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/A_DOUT_ARST_N_net , 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/A_DOUT_SRST_N_net , 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/A_DIN_net[17] , 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/A_DIN_net[16] , 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/A_DIN_net[15] , 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/A_DIN_net[14] , 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/A_DIN_net[13] , 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/A_DIN_net[12] , 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/A_DIN_net[11] , 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/A_DIN_net[10] , 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/A_DIN_net[9] , 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/A_DIN_net[8] , 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/A_DIN_net[7] , 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/A_DIN_net[6] , 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/A_DIN_net[5] , 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/A_DIN_net[4] , 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/A_DIN_net[3] , 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/A_DIN_net[2] , 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/A_DIN_net[1] , 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/A_DIN_net[0] , 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/A_ADDR_net[13] , 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/A_ADDR_net[12] , 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/A_ADDR_net[11] , 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/A_ADDR_net[10] , 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/A_ADDR_net[9] , 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/A_ADDR_net[8] , 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/A_ADDR_net[7] , 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/A_ADDR_net[6] , 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/A_ADDR_net[5] , 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/A_ADDR_net[4] , 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/A_ADDR_net[3] , 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/A_ADDR_net[2] , 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/A_ADDR_net[1] , 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/A_ADDR_net[0] , 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/A_WEN_net[1] , 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/A_WEN_net[0] , 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/B_CLK_net , 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/B_DOUT_CLK_net , 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/B_ARST_N_net , 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/B_DOUT_EN_net , 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/B_BLK_net[2] , 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/B_BLK_net[1] , 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/B_BLK_net[0] , 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/B_DOUT_ARST_N_net , 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/B_DOUT_SRST_N_net , 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/B_DIN_net[17] , 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/B_DIN_net[16] , 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/B_DIN_net[15] , 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/B_DIN_net[14] , 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/B_DIN_net[13] , 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/B_DIN_net[12] , 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/B_DIN_net[11] , 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/B_DIN_net[10] , 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/B_DIN_net[9] , 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/B_DIN_net[8] , 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/B_DIN_net[7] , 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/B_DIN_net[6] , 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/B_DIN_net[5] , 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/B_DIN_net[4] , 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/B_DIN_net[3] , 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/B_DIN_net[2] , 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/B_DIN_net[1] , 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/B_DIN_net[0] , 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/B_ADDR_net[13] , 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/B_ADDR_net[12] , 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/B_ADDR_net[11] , 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/B_ADDR_net[10] , 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/B_ADDR_net[9] , 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/B_ADDR_net[8] , 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/B_ADDR_net[7] , 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/B_ADDR_net[6] , 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/B_ADDR_net[5] , 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/B_ADDR_net[4] , 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/B_ADDR_net[3] , 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/B_ADDR_net[2] , 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/B_ADDR_net[1] , 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/B_ADDR_net[0] , 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/B_WEN_net[1] , 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/B_WEN_net[0] , 
        \GPIO_OUT_1_obuf[4]/U0/DOUT1 , \GPIO_OUT_1_obuf[4]/U0/DOUT , 
        \GPIO_OUT_1_obuf[4]/U0/EOUT1 , \GPIO_OUT_1_obuf[4]/U0/EOUT , 
        \GPIO_OUT_1_obuf[0]/U0/DOUT1 , \GPIO_OUT_1_obuf[0]/U0/DOUT , 
        \GPIO_OUT_1_obuf[0]/U0/EOUT1 , \GPIO_OUT_1_obuf[0]/U0/EOUT , 
        \GPIO_OUT_1_obuf[3]/U0/DOUT1 , \GPIO_OUT_1_obuf[3]/U0/DOUT , 
        \GPIO_OUT_1_obuf[3]/U0/EOUT1 , \GPIO_OUT_1_obuf[3]/U0/EOUT , 
        \FCCC_0/CCC_INST/CLK0_net , \FCCC_0/CCC_INST/CLK1_net , 
        \FCCC_0/CCC_INST/CLK2_net , \FCCC_0/CCC_INST/CLK3_net , 
        \FCCC_0/CCC_INST/NGMUX0_SEL_net , 
        \FCCC_0/CCC_INST/NGMUX1_SEL_net , 
        \FCCC_0/CCC_INST/NGMUX2_SEL_net , 
        \FCCC_0/CCC_INST/NGMUX3_SEL_net , 
        \FCCC_0/CCC_INST/NGMUX0_HOLD_N_net , 
        \FCCC_0/CCC_INST/NGMUX1_HOLD_N_net , 
        \FCCC_0/CCC_INST/NGMUX2_HOLD_N_net , 
        \FCCC_0/CCC_INST/NGMUX3_HOLD_N_net , 
        \FCCC_0/CCC_INST/NGMUX0_ARST_N_net , 
        \FCCC_0/CCC_INST/NGMUX1_ARST_N_net , 
        \FCCC_0/CCC_INST/NGMUX2_ARST_N_net , 
        \FCCC_0/CCC_INST/NGMUX3_ARST_N_net , 
        \FCCC_0/CCC_INST/PLL_BYPASS_N_net , 
        \FCCC_0/CCC_INST/PLL_ARST_N_net , 
        \FCCC_0/CCC_INST/PLL_POWERDOWN_N_net , 
        \FCCC_0/CCC_INST/GPD0_ARST_N_net , 
        \FCCC_0/CCC_INST/GPD1_ARST_N_net , 
        \FCCC_0/CCC_INST/GPD2_ARST_N_net , 
        \FCCC_0/CCC_INST/GPD3_ARST_N_net , 
        \FCCC_0/CCC_INST/PRESET_N_net , \FCCC_0/CCC_INST/PCLK_net , 
        \FCCC_0/CCC_INST/PSEL_net , \FCCC_0/CCC_INST/PENABLE_net , 
        \FCCC_0/CCC_INST/PWRITE_net , \FCCC_0/CCC_INST/PADDR_net[7] , 
        \FCCC_0/CCC_INST/PADDR_net[6] , \FCCC_0/CCC_INST/PADDR_net[5] , 
        \FCCC_0/CCC_INST/PADDR_net[4] , \FCCC_0/CCC_INST/PADDR_net[3] , 
        \FCCC_0/CCC_INST/PADDR_net[2] , 
        \FCCC_0/CCC_INST/PWDATA_net[7] , 
        \FCCC_0/CCC_INST/PWDATA_net[6] , 
        \FCCC_0/CCC_INST/PWDATA_net[5] , 
        \FCCC_0/CCC_INST/PWDATA_net[4] , 
        \FCCC_0/CCC_INST/PWDATA_net[3] , 
        \FCCC_0/CCC_INST/PWDATA_net[2] , 
        \FCCC_0/CCC_INST/PWDATA_net[1] , 
        \FCCC_0/CCC_INST/PWDATA_net[0] , \GPIO_OUT_1_obuf[2]/U0/DOUT1 , 
        \GPIO_OUT_1_obuf[2]/U0/DOUT , \GPIO_OUT_1_obuf[2]/U0/EOUT1 , 
        \GPIO_OUT_1_obuf[2]/U0/EOUT , \GPIO_OUT_1_obuf[7]/U0/DOUT1 , 
        \GPIO_OUT_1_obuf[7]/U0/DOUT , \GPIO_OUT_1_obuf[7]/U0/EOUT1 , 
        \GPIO_OUT_1_obuf[7]/U0/EOUT , \GPIO_OUT_1_obuf[5]/U0/DOUT1 , 
        \GPIO_OUT_1_obuf[5]/U0/DOUT , \GPIO_OUT_1_obuf[5]/U0/EOUT1 , 
        \GPIO_OUT_1_obuf[5]/U0/EOUT , 
        \hello_regs_MSS_0/MMUART_0_RXD_PAD/YIN , 
        \GPIO_OUT_1_obuf[6]/U0/DOUT1 , \GPIO_OUT_1_obuf[6]/U0/DOUT , 
        \GPIO_OUT_1_obuf[6]/U0/EOUT1 , \GPIO_OUT_1_obuf[6]/U0/EOUT , 
        \GPIO_OUT_1_obuf[1]/U0/DOUT1 , \GPIO_OUT_1_obuf[1]/U0/DOUT , 
        \GPIO_OUT_1_obuf[1]/U0/EOUT1 , \GPIO_OUT_1_obuf[1]/U0/EOUT , 
        \MSS_RESET_N_M2F_obuf/U0/DOUT1 , 
        \MSS_RESET_N_M2F_obuf/U0/DOUT , 
        \MSS_RESET_N_M2F_obuf/U0/EOUT1 , 
        \MSS_RESET_N_M2F_obuf/U0/EOUT , CFG0_GND_INST_NET, 
        \FCCC_0/GL1_INST/U0_RGB1_YR , 
        \FCCC_0/GL1_INST/U0_RGB1_RGB0_rgbr_net_1 , 
        \FCCC_0/GL1_INST/U0_RGB1_RGB1_rgbr_net_1 , 
        \FCCC_0/GL1_INST/U0_RGB1_RGB2_rgbr_net_1 , 
        \FCCC_0/GL1_INST/U0_RGB1_RGB3_rgbr_net_1 , 
        \FCCC_0/GL1_INST/U0_RGB1_RGB4_rgbr_net_1 , 
        \FCCC_0/GL1_INST/U0_RGB1_RGB5_rgbr_net_1 , 
        \FCCC_0/GL1_INST/U0_RGB1_RGB5_rgbl_net_1 , 
        \FCCC_0/GL1_INST/U0_RGB1_RGB6_rgbr_net_1 , 
        \FCCC_0/GL1_INST/U0_RGB1_RGB6_rgbl_net_1 , 
        \FCCC_0/GL1_INST/U0_RGB1_RGB7_rgbr_net_1 , 
        \FCCC_0/GL1_INST/U0_RGB1_RGB7_rgbl_net_1 , 
        \FCCC_0/GL1_INST/U0_RGB1_RGB8_rgbr_net_1 , 
        \FCCC_0/GL1_INST/U0_RGB1_RGB8_rgbl_net_1 , 
        \FCCC_0/GL1_INST/U0_RGB1_RGB9_rgbr_net_1 , 
        \FCCC_0/GL1_INST/U0_RGB1_RGB9_rgbl_net_1 , 
        \FCCC_0/GL1_INST/U0_RGB1_RGB10_rgbr_net_1 , 
        \FCCC_0/GL1_INST/U0_RGB1_RGB10_rgbl_net_1 , 
        \FCCC_0/GL1_INST/U0_RGB1_RGB11_rgbr_net_1 , 
        \FCCC_0/GL1_INST/U0_RGB1_RGB11_rgbl_net_1 , 
        \FCCC_0/GL1_INST/U0_RGB1_RGB12_rgbr_net_1 , 
        \FCCC_0/GL1_INST/U0_RGB1_RGB12_rgbl_net_1 , 
        \FCCC_0/GL1_INST/U0_RGB1_RGB13_rgbr_net_1 , 
        \FCCC_0/GL1_INST/U0_RGB1_RGB13_rgbl_net_1 , 
        \FCCC_0/GL1_INST/U0_RGB1_RGB14_rgbr_net_1 , 
        \FCCC_0/GL1_INST/U0_RGB1_RGB14_rgbl_net_1 , 
        \FCCC_0/GL1_INST/U0_RGB1_RGB15_rgbr_net_1 , 
        \FCCC_0/GL1_INST/U0_RGB1_RGB15_rgbl_net_1 , 
        \FCCC_0/GL1_INST/U0_RGB1_RGB16_rgbr_net_1 , 
        \FCCC_0/GL1_INST/U0_RGB1_RGB16_rgbl_net_1 , 
        \FCCC_0/GL1_INST/U0_RGB1_RGB17_rgbr_net_1 , 
        \FCCC_0/GL1_INST/U0_RGB1_RGB17_rgbl_net_1 , 
        \FCCC_0/GL1_INST/U0_RGB1_RGB18_rgbr_net_1 , 
        \FCCC_0/GL1_INST/U0_RGB1_RGB18_rgbl_net_1 , 
        \FCCC_0/GL1_INST/U0_RGB1_RGB19_rgbr_net_1 , 
        \hello_regs_MSS_0/MSS_ADLIB_INST_RNIUO3B/U0_RGB1_YR , 
        \hello_regs_MSS_0/MSS_ADLIB_INST_RNIUO3B/U0_RGB1_RGB0_rgbr_net_1 , 
        \hello_regs_MSS_0/MSS_ADLIB_INST_RNIUO3B/U0_RGB1_RGB1_rgbr_net_1 , 
        \hello_regs_MSS_0/MSS_ADLIB_INST_RNIUO3B/U0_RGB1_RGB2_rgbr_net_1 , 
        \hello_regs_MSS_0/MSS_ADLIB_INST_RNIUO3B/U0_RGB1_RGB3_rgbr_net_1 , 
        \hello_regs_MSS_0/MSS_ADLIB_INST_RNIUO3B/U0_RGB1_RGB4_rgbr_net_1 , 
        \hello_regs_MSS_0/MSS_ADLIB_INST_RNIUO3B/U0_RGB1_RGB5_rgbr_net_1 , 
        \hello_regs_MSS_0/MSS_ADLIB_INST_RNIUO3B/U0_RGB1_RGB6_rgbr_net_1 , 
        \hello_regs_MSS_0/MSS_ADLIB_INST_RNIUO3B/U0_YNn_GSouth , 
        \FCCC_0/GL1_INST/U0_YNn_GSouth , AFLSDF_VCC, AFLSDF_GND, 
        AFLSDF_INV_0_net_1, AFLSDF_INV_1_net_1, AFLSDF_INV_2_net_1, 
        AFLSDF_INV_3_net_1, AFLSDF_INV_4_net_1, AFLSDF_INV_5_net_1, 
        AFLSDF_INV_6_net_1, AFLSDF_INV_7_net_1, AFLSDF_INV_8_net_1, 
        AFLSDF_INV_9_net_1, AFLSDF_INV_10_net_1, AFLSDF_INV_11_net_1, 
        AFLSDF_INV_12_net_1, AFLSDF_INV_13_net_1, AFLSDF_INV_14_net_1, 
        AFLSDF_INV_15_net_1, AFLSDF_INV_16_net_1, AFLSDF_INV_17_net_1, 
        AFLSDF_INV_18_net_1, AFLSDF_INV_19_net_1, AFLSDF_INV_20_net_1, 
        AFLSDF_INV_21_net_1, AFLSDF_INV_22_net_1, AFLSDF_INV_23_net_1, 
        AFLSDF_INV_24_net_1, AFLSDF_INV_25_net_1, AFLSDF_INV_26_net_1, 
        AFLSDF_INV_27_net_1, AFLSDF_INV_28_net_1, AFLSDF_INV_29_net_1, 
        AFLSDF_INV_30_net_1, AFLSDF_INV_31_net_1, AFLSDF_INV_32_net_1, 
        AFLSDF_INV_33_net_1, AFLSDF_INV_34_net_1, AFLSDF_INV_35_net_1, 
        AFLSDF_INV_36_net_1, AFLSDF_INV_37_net_1, AFLSDF_INV_38_net_1, 
        AFLSDF_INV_39_net_1, AFLSDF_INV_40_net_1, AFLSDF_INV_41_net_1, 
        AFLSDF_INV_42_net_1, AFLSDF_INV_43_net_1, AFLSDF_INV_44_net_1, 
        AFLSDF_INV_45_net_1, AFLSDF_INV_46_net_1, AFLSDF_INV_47_net_1, 
        AFLSDF_INV_48_net_1, AFLSDF_INV_49_net_1, AFLSDF_INV_50_net_1, 
        AFLSDF_INV_51_net_1, AFLSDF_INV_52_net_1, AFLSDF_INV_53_net_1, 
        AFLSDF_INV_54_net_1, AFLSDF_INV_55_net_1, AFLSDF_INV_56_net_1, 
        AFLSDF_INV_57_net_1, AFLSDF_INV_58_net_1, AFLSDF_INV_59_net_1, 
        AFLSDF_INV_60_net_1, AFLSDF_INV_61_net_1, AFLSDF_INV_62_net_1, 
        AFLSDF_INV_63_net_1, AFLSDF_INV_64_net_1, AFLSDF_INV_65_net_1, 
        AFLSDF_INV_66_net_1, AFLSDF_INV_67_net_1, AFLSDF_INV_68_net_1, 
        AFLSDF_INV_69_net_1, AFLSDF_INV_70_net_1, AFLSDF_INV_71_net_1, 
        AFLSDF_INV_72_net_1, AFLSDF_INV_73_net_1, AFLSDF_INV_74_net_1, 
        AFLSDF_INV_75_net_1, AFLSDF_INV_76_net_1, AFLSDF_INV_77_net_1, 
        AFLSDF_INV_78_net_1, AFLSDF_INV_79_net_1, AFLSDF_INV_80_net_1, 
        AFLSDF_INV_81_net_1, AFLSDF_INV_82_net_1, AFLSDF_INV_83_net_1, 
        AFLSDF_INV_84_net_1, AFLSDF_INV_85_net_1, AFLSDF_INV_86_net_1, 
        AFLSDF_INV_87_net_1, AFLSDF_INV_88_net_1, AFLSDF_INV_89_net_1, 
        AFLSDF_INV_90_net_1, AFLSDF_INV_91_net_1, AFLSDF_INV_92_net_1, 
        AFLSDF_INV_93_net_1, AFLSDF_INV_94_net_1, AFLSDF_INV_95_net_1, 
        AFLSDF_INV_96_net_1, AFLSDF_INV_97_net_1, AFLSDF_INV_98_net_1, 
        AFLSDF_INV_99_net_1, AFLSDF_INV_100_net_1, 
        AFLSDF_INV_101_net_1, AFLSDF_INV_102_net_1, 
        AFLSDF_INV_103_net_1, AFLSDF_INV_104_net_1, 
        AFLSDF_INV_105_net_1, AFLSDF_INV_106_net_1, 
        AFLSDF_INV_107_net_1, AFLSDF_INV_108_net_1, 
        AFLSDF_INV_109_net_1, AFLSDF_INV_110_net_1, 
        AFLSDF_INV_111_net_1, AFLSDF_INV_112_net_1, 
        AFLSDF_INV_113_net_1, AFLSDF_INV_114_net_1, 
        AFLSDF_INV_115_net_1, AFLSDF_INV_116_net_1, 
        AFLSDF_INV_117_net_1, AFLSDF_INV_118_net_1, 
        AFLSDF_INV_119_net_1, AFLSDF_INV_120_net_1, 
        AFLSDF_INV_121_net_1, AFLSDF_INV_122_net_1, 
        AFLSDF_INV_123_net_1, AFLSDF_INV_124_net_1, 
        AFLSDF_INV_125_net_1, AFLSDF_INV_126_net_1, 
        AFLSDF_INV_127_net_1, AFLSDF_INV_128_net_1, 
        AFLSDF_INV_129_net_1, AFLSDF_INV_130_net_1, 
        AFLSDF_INV_131_net_1, AFLSDF_INV_132_net_1, 
        AFLSDF_INV_133_net_1, AFLSDF_INV_134_net_1, 
        AFLSDF_INV_135_net_1, AFLSDF_INV_136_net_1, 
        AFLSDF_INV_137_net_1, AFLSDF_INV_138_net_1, 
        AFLSDF_INV_139_net_1, AFLSDF_INV_140_net_1, 
        AFLSDF_INV_141_net_1, AFLSDF_INV_142_net_1, 
        AFLSDF_INV_143_net_1, AFLSDF_INV_144_net_1, 
        AFLSDF_INV_145_net_1, AFLSDF_INV_146_net_1, 
        AFLSDF_INV_147_net_1;
    wire GND_power_net1;
    wire VCC_power_net1;
    assign GND = GND_power_net1;
    assign AFLSDF_GND = GND_power_net1;
    assign VCC = VCC_power_net1;
    assign AFLSDF_VCC = VCC_power_net1;
    
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_80_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB13_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_0__1_sqmuxa ), .ALn(
        AFLSDF_INV_0_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(GND), 
        .Q(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_80_set_net_1 ));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_285  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PADDR_net[8] ), 
        .IPB(
        \hello_regs_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[12] ), 
        .IPC());
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_142  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(), .IPB(
        \hello_regs_MSS_0/MSS_ADLIB_INST/SPI1_CLK_IN_net ), .IPC());
    CFG3 #( .INIT(8'h80) )  
        \reg_apb_wrp_0/reg16x8_0/mem_4__1_sqmuxa_0_a2  (.A(
        \reg_apb_wrp_0/reg16x8_0/N_648 ), .B(N_637), .C(N_638), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_4__1_sqmuxa ));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_66  (.A(
        GND), .B(VCC), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[27] ), .IPB(
        \hello_regs_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[0] ), 
        .IPC());
    SLE \COREAPBLSRAM_0/PRDATA_reg[20]  (.D(
        \COREAPBLSRAM_0.lsram_width32_PRDATA[20] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB10_rgbr_net_1 ), .EN(
        \COREAPBLSRAM_0.PRDATA4 ), .ALn(
        \hello_regs_MSS_0/MSS_ADLIB_INST_RNIUO3B/U0_RGB1_RGB2_rgbr_net_1 )
        , .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \COREAPBLSRAM_0.PRDATA_reg[20] ));
    SLE \COREAPBLSRAM_0/PRDATA_reg[19]  (.D(
        \COREAPBLSRAM_0.lsram_width32_PRDATA[19] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB9_rgbr_net_1 ), .EN(
        \COREAPBLSRAM_0.PRDATA4 ), .ALn(
        \hello_regs_MSS_0/MSS_ADLIB_INST_RNIUO3B/U0_RGB1_RGB1_rgbr_net_1 )
        , .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \COREAPBLSRAM_0.PRDATA_reg[19] ));
    CFG2_IP_BC 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/CFG_23  
        (.B(\CoreAPB3_0_APBmslave5_PWDATA[29] ), .C(
        \COREAPBLSRAM_0/wen ), .IPB(
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/B_DIN_net[14] )
        , .IPC(
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/B_WEN_net[1] )
        );
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/mem_10__RNISPDJ[2]  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_99_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_170_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_10_rs[2] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_10_[2]_net_1 ));
    INV_BA AFLSDF_INV_64 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_74_net_1 ), .Y(
        AFLSDF_INV_64_net_1));
    CFG3 #( .INIT(8'hF2) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_179  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_7_[0]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_641 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_179_i ));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_93  (.A(
        VCC), .B(VCC), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/RX_DVF_net ), .IPB(), .IPC());
    sdf_IOPAD_TRI \GPIO_OUT_1_obuf[6]/U0/U_IOPAD  (.PAD(GPIO_OUT_1[6]), 
        .D(\GPIO_OUT_1_obuf[6]/U0/DOUT ), .E(
        \GPIO_OUT_1_obuf[6]/U0/EOUT ));
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_data_out8_46  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_1_[7]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_651 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_46_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_10_[0]  (.D(
        \CoreAPB3_0_APBmslave5_PWDATA[0] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB8_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_10__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_206_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_10_rs[0] ));
    CFG4 #( .INIT(16'hFFFE) )  
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_12[4]  (.A(
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_1[4]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_3[4]_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_2[4]_net_1 ), .D(
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_0[4]_net_1 ), .Y(
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_12[4]_net_1 ));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_50  (.A(
        GND), .B(VCC), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[4] ), .IPB(), 
        .IPC());
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_185  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/MMUART0_RXD_F2H_SCP_net ), 
        .IPB(\hello_regs_MSS_0/MSS_ADLIB_INST/I2C0_SCL_F2H_SCP_net ), 
        .IPC());
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_50_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB15_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_7__1_sqmuxa ), .ALn(
        AFLSDF_INV_1_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(GND), 
        .Q(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_50_set_net_1 ));
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_data_out8_31  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_2_[3]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_642 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_31_net_1 ));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_52_set_RNIC2OE  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_52_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_227_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_7_rs[4] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_7_[4]_net_1 ));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_187  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/MMUART0_SCK_F2H_SCP_net ), 
        .IPB(), .IPC());
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_78  (.A(
        VCC), .B(VCC), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[12] ), 
        .IPB(
        \hello_regs_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[19] ), 
        .IPC());
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_246  (
        .A(VCC), .B(GND), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[58] ), 
        .IPB(\hello_regs_MSS_0/MSS_ADLIB_INST/F_WSTRB_net[6] ), .IPC());
    CFG4 #( .INIT(16'hFFFE) )  
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_12[1]  (.A(
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_1[1]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_3[1]_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_2[1]_net_1 ), .D(
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_0[1]_net_1 ), .Y(
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_12[1]_net_1 ));
    SLE_IP_EN 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/FF_12  
        (.EN(VCC), .IPENn());
    CFG2_IP_BC 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/CFG_1  
        (.B(\CoreAPB3_0_APBmslave5_PWDATA[16] ), .C(GND), .IPB(
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/B_DIN_net[0] )
        , .IPC(
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/B_ADDR_net[0] )
        );
    SLE \reg_apb_wrp_0/reg16x8_0/mem_9_[5]  (.D(
        \CoreAPB3_0_APBmslave5_PWDATA[5] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB14_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_9__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_200_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_9_rs[5] ));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_221  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[5] ), 
        .IPB(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[17] ), 
        .IPC());
    SLE_IP_EN 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/FF_2  
        (.EN(VCC), .IPENn());
    CFG3 #( .INIT(8'hF2) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_196  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_9_[3]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_643 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_196_i ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_112_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB16_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_14__1_sqmuxa ), .ALn(
        AFLSDF_INV_2_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(GND), 
        .Q(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_112_set_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_29_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB6_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_2__1_sqmuxa ), .ALn(
        AFLSDF_INV_3_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(GND), 
        .Q(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_29_set_net_1 ));
    INV_BA AFLSDF_INV_53 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_59_net_1 ), .Y(
        AFLSDF_INV_53_net_1));
    CFG3 #( .INIT(8'hF2) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_130  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_3_[2]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_655 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_130_i ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_226_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_90_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_226_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_226_rs_net_1 ));
    CFG4 #( .INIT(16'h7530) )  
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_6[1]  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_4_[1]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/mem_1_[1]_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/N_651 ), .D(
        \reg_apb_wrp_0/reg16x8_0/N_648 ), .Y(
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_6[1]_net_1 ));
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_data_out8_92  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_11_[4]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_649 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_92_net_1 ));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_48  (.A(
        GND), .B(VCC), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[2] ), .IPB(), 
        .IPC());
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_125_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB12_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_3__1_sqmuxa ), .ALn(
        AFLSDF_INV_4_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(GND), 
        .Q(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_125_set_net_1 ));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_92  (.A(
        VCC), .B(VCC), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/RX_CLKPF_net ), .IPB(
        \hello_regs_MSS_0/MSS_ADLIB_INST/RX_ERRF_net ), .IPC());
    SLE_IP_EN 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/FF_34  
        (.EN(VCC), .IPENn(AFLSDF_INV_5_net_1));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_5_[3]  (.D(
        \CoreAPB3_0_APBmslave5_PWDATA[3] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB8_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_5__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_193_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_5_rs[3] ));
    IOENFF_BYPASS \GPIO_OUT_1_obuf[0]/U0/U_IOENFF  (.A(
        \GPIO_OUT_1_obuf[0]/U0/EOUT1 ), .Y(
        \GPIO_OUT_1_obuf[0]/U0/EOUT ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_42_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB11_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_1__1_sqmuxa ), .ALn(
        AFLSDF_INV_6_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(GND), 
        .Q(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_42_set_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_127_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB15_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_3__1_sqmuxa ), .ALn(
        AFLSDF_INV_7_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(GND), 
        .Q(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_127_set_net_1 ));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_0  (.A(
        N_537_i_0), .B(VCC), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_HM0_READY_net ), .IPB(), 
        .IPC());
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_23  (.A(
        VCC), .B(GND), .C(VCC), .IPA(), .IPB(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_TRANS1_net ), .IPC());
    CFG3 #( .INIT(8'h02) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_119  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_14_[7]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_650 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_119_net_1 ));
    CFG2_IP_BC 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/CFG_2  
        (.B(\CoreAPB3_0_APBmslave5_PWDATA[8] ), .C(GND), .IPB(
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/A_DIN_net[9] )
        , .IPC(
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/A_ADDR_net[1] )
        );
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_data_out8_89  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_11_[1]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_649 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_89_net_1 ));
    CFG3 #( .INIT(8'hF2) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_182  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_11_[0]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_649 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_182_i ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_162_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_29_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_162_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_162_rs_net_1 ));
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_data_out8_8  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_4_[6]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_648 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_8_net_1 ));
    CFG3 #( .INIT(8'hF2) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_230  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_11_[4]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_649 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_230_i ));
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_data_out8_23  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_12_[7]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_644 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_23_net_1 ));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_182  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/MGPIO27B_F2H_GPIN_net ), .IPB(
        ), .IPC());
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_148  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/MGPIO1A_F2H_GPIN_net ), .IPB(
        \hello_regs_MSS_0/MSS_ADLIB_INST/CAN_TX_EBL_F2H_SCP_net ), 
        .IPC());
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_134  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/I2C0_BCLK_net ), .IPB(), .IPC(
        ));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_151_rs_RNIC10H  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_87_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_151_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_0_rs[7] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_0_[7]_net_1 ));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_111  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/FAB_XDATAIN_net[3] ), .IPB(
        \hello_regs_MSS_0/MSS_ADLIB_INST/FAB_VSTATUS_net[0] ), .IPC());
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_225_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_50_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_225_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_225_rs_net_1 ));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_34  (.A(
        VCC), .B(GND), .C(VCC), .IPA(), .IPB(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[17] ), .IPC());
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_231_rs_RNILT5G  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_3_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_231_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_7_rs[6] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_7_[6]_net_1 ));
    CFG4 #( .INIT(16'h7350) )  
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_1[2]  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_15_[2]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/mem_14_[2]_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/N_654 ), .D(
        \reg_apb_wrp_0/reg16x8_0/N_650 ), .Y(
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_1[2]_net_1 ));
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_data_out8_90  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_11_[2]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_649 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_90_net_1 ));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_215_rs_RNI5OUS  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_111_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_215_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_13_rs[7] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_13_[7]_net_1 ));
    RGB \FCCC_0/GL1_INST/U0_RGB1_RGB9  (.An(\FCCC_0/GL1_INST/U0_YNn ), 
        .ENn(GND), .YL(\FCCC_0/GL1_INST/U0_RGB1_RGB9_rgbl_net_1 ), .YR(
        \FCCC_0/GL1_INST/U0_RGB1_RGB9_rgbr_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_5_[4]  (.D(
        \CoreAPB3_0_APBmslave5_PWDATA[4] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB8_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_5__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_195_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_5_rs[4] ));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_9_[7]  (.D(
        \CoreAPB3_0_APBmslave5_PWDATA[7] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB18_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_9__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_204_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_9_rs[7] ));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_279  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PADDR_net[2] ), 
        .IPB(
        \hello_regs_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[6] ), 
        .IPC());
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_56_set_RNIQBFK  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_56_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_250_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_15_rs[3] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_15_[3]_net_1 ));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_65  (.A(
        GND), .B(VCC), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[26] ), .IPB(
        \hello_regs_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PSLVERR_net ), 
        .IPC());
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_286  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PADDR_net[9] ), 
        .IPB(
        \hello_regs_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[13] ), 
        .IPC());
    INV_BA AFLSDF_INV_55 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_113_net_1 ), .Y(
        AFLSDF_INV_55_net_1));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_22  (.A(
        VCC), .B(GND), .C(VCC), .IPA(), .IPB(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_SIZE_net[1] ), .IPC());
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_36_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB10_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_6__1_sqmuxa ), .ALn(
        AFLSDF_INV_8_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(GND), 
        .Q(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_36_set_net_1 ));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/mem_14__RNI44NB[1]  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_113_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_217_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_14_rs[1] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_14_[1]_net_1 ));
    IP_INTERFACE \FCCC_0/CCC_INST/IP_INTERFACE_3  (.A(GND), .B(GND), 
        .C(VCC), .IPA(\FCCC_0/CCC_INST/PRESET_N_net ), .IPB(
        \FCCC_0/CCC_INST/NGMUX1_SEL_net ), .IPC(
        \FCCC_0/CCC_INST/PWDATA_net[1] ));
    INV_BA AFLSDF_INV_20 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_110_net_1 ), .Y(
        AFLSDF_INV_20_net_1));
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_data_out8_12  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_5_[0]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_653 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_12_net_1 ));
    SLE_IP_EN 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/FF_23  
        (.EN(VCC), .IPENn());
    INV_BA AFLSDF_INV_140 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_12_net_1 ), .Y(
        AFLSDF_INV_140_net_1));
    IP_INTERFACE \FCCC_0/CCC_INST/IP_INTERFACE_2  (.A(VCC), .B(GND), 
        .C(VCC), .IPA(\FCCC_0/CCC_INST/PCLK_net ), .IPB(
        \FCCC_0/CCC_INST/NGMUX0_SEL_net ), .IPC(
        \FCCC_0/CCC_INST/PWDATA_net[0] ));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_106  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(), .IPB(
        \hello_regs_MSS_0/MSS_ADLIB_INST/FAB_TXREADY_net ), .IPC());
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_103_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB8_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_10__1_sqmuxa ), .ALn(
        AFLSDF_INV_9_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(GND), 
        .Q(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_103_set_net_1 ));
    RGB \hello_regs_MSS_0/MSS_ADLIB_INST_RNIUO3B/U0_RGB1_RGB1  (.An(
        \hello_regs_MSS_0/MSS_ADLIB_INST_RNIUO3B/U0_YNn ), .ENn(GND), 
        .YL(), .YR(
        \hello_regs_MSS_0/MSS_ADLIB_INST_RNIUO3B/U0_RGB1_RGB1_rgbr_net_1 )
        );
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_124  (
        .A(VCC), .B(GND), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/FAB_IDDIG_net ), .IPB(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[6] ), .IPC()
        );
    SLE \reg_apb_wrp_0/reg16x8_0/mem_11_[5]  (.D(
        \CoreAPB3_0_APBmslave5_PWDATA[5] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB4_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_11__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_232_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_11_rs[5] ));
    INV_BA AFLSDF_INV_47 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_85_net_1 ), .Y(
        AFLSDF_INV_47_net_1));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_136_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_net_1 ), .EN(VCC), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_136_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_136_rs_net_1 ));
    SLE_IP_EN 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/FF_14  
        (.EN(VCC), .IPENn());
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_278  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[2] ), 
        .IPB(
        \hello_regs_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[5] ), 
        .IPC());
    CFG4 #( .INIT(16'hECA0) )  \CoreAPB3_0/u_mux_p_to_b3/PRDATA_0[8]  
        (.A(\CoreAPB3_0/u_mux_p_to_b3/N_636 ), .B(
        \COREAPBLSRAM_0.PRDATA4 ), .C(\COREAPBLSRAM_0.PRDATA_reg[8] ), 
        .D(\COREAPBLSRAM_0.lsram_width32_PRDATA[8] ), .Y(
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[8] ));
    CFG1_IP_B 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/CFG_34  
        (.B(GND), .IPB(
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/A_DIN_net[17] )
        );
    CFG3 #( .INIT(8'hF2) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_181  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_7_[1]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_641 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_181_i ));
    CFG3 #( .INIT(8'hF2) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_156  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_1_[4]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_651 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_156_i ));
    CFG3 #( .INIT(8'hF2) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_134  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_3_[6]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_655 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_134_i ));
    INV_BA AFLSDF_INV_9 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_103_net_1 ), .Y(
        AFLSDF_INV_9_net_1));
    CFG3 #( .INIT(8'hF2) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_235  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_8_[0]_net_1 ), .B(N_639), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_235_i ));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_set_RNIU3D21  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_136_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_4_rs[0] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_4_[0]_net_1 ));
    CFG4 #( .INIT(16'h7350) )  
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_0[1]  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_11_[1]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/mem_10_[1]_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/N_649 ), .D(
        \reg_apb_wrp_0/reg16x8_0/N_647 ), .Y(
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_0[1]_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_218_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_114_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_218_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_218_rs_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_5_[0]  (.D(
        \CoreAPB3_0_APBmslave5_PWDATA[0] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB9_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_5__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_187_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_5_rs[0] ));
    IP_INTERFACE \FCCC_0/CCC_INST/IP_INTERFACE_5  (.A(VCC), .B(VCC), 
        .C(VCC), .IPA(), .IPB(\FCCC_0/CCC_INST/NGMUX1_HOLD_N_net ), 
        .IPC(\FCCC_0/CCC_INST/PWDATA_net[3] ));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_83  (.A(
        VCC), .B(VCC), .C(VCC), .IPA(), .IPB(
        \hello_regs_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[24] ), 
        .IPC());
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_140_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_65_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_140_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_140_rs_net_1 ));
    CFG2 #( .INIT(4'h8) )  
        \CoreAPB3_0/u_mux_p_to_b3/PRDATA_0_iv_0_a2_2_0[6]  (.A(N_639), 
        .B(\GPIO_OUT_1_c[6] ), .Y(
        \CoreAPB3_0/u_mux_p_to_b3/PRDATA_0_iv_0_a2_2_0[6]_net_1 ));
    CFG4 #( .INIT(16'hECA0) )  \CoreAPB3_0/u_mux_p_to_b3/PRDATA_0[15]  
        (.A(\CoreAPB3_0/u_mux_p_to_b3/N_636 ), .B(
        \COREAPBLSRAM_0.PRDATA4 ), .C(\COREAPBLSRAM_0.PRDATA_reg[15] ), 
        .D(\COREAPBLSRAM_0.lsram_width32_PRDATA[15] ), .Y(
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[15] ));
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_data_out8_10  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_4_[7]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_648 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_10_net_1 ));
    CFG4 #( .INIT(16'h7350) )  
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_5[4]  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_0_[4]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/mem_7_[4]_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/N_645 ), .D(
        \reg_apb_wrp_0/reg16x8_0/N_641 ), .Y(
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_5[4]_net_1 ));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_188  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/MGPIO30B_F2H_GPIN_net ), .IPB(
        ), .IPC());
    CFG2_IP_BC 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/CFG_12  
        (.B(\CoreAPB3_0_APBmslave5_PWDATA[3] ), .C(
        \CoreAPB3_0_APBmslave5_PADDR[0] ), .IPB(
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/A_DIN_net[3] )
        , .IPC(
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/A_ADDR_net[5] )
        );
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_255_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_61_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_255_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_255_rs_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_115_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB15_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_14__1_sqmuxa ), .ALn(
        AFLSDF_INV_10_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(GND)
        , .Q(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_115_set_net_1 ));
    CFG4 #( .INIT(16'h0080) )  
        \reg_apb_wrp_0/reg16x8_0/WRITE_GEN.mem_13__2_i_a2[5]  (.A(
        \CoreAPB3_0_APBmslave5_PADDR[2] ), .B(
        \CoreAPB3_0_APBmslave5_PADDR[5] ), .C(
        \CoreAPB3_0_APBmslave5_PADDR[4] ), .D(
        \CoreAPB3_0_APBmslave5_PADDR[3] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/N_646 ));
    CFG4 #( .INIT(16'h7350) )  
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_0[2]  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_11_[2]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/mem_10_[2]_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/N_649 ), .D(
        \reg_apb_wrp_0/reg16x8_0/N_647 ), .Y(
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_0[2]_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_117_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB11_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_14__1_sqmuxa ), .ALn(
        AFLSDF_INV_11_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(GND)
        , .Q(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_117_set_net_1 ));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_38  (.A(
        GND), .B(VCC), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[21] ), .IPB(), 
        .IPC());
    INV_BA AFLSDF_INV_76 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_13_net_1 ), .Y(
        AFLSDF_INV_76_net_1));
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_data_out8_85  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_0_[5]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_645 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_85_net_1 ));
    IOOUTFF_BYPASS \GPIO_OUT_1_obuf[6]/U0/U_IOOUTFF  (.A(
        \GPIO_OUT_1_obuf[6]/U0/DOUT1 ), .Y(
        \GPIO_OUT_1_obuf[6]/U0/DOUT ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_233_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_1_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_233_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_233_rs_net_1 ));
    CFG4 #( .INIT(16'h7530) )  
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_3[0]  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_2_[0]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/mem_13_[0]_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/N_646 ), .D(
        \reg_apb_wrp_0/reg16x8_0/N_642 ), .Y(
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_3[0]_net_1 ));
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_data_out8_64  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_8_[2]_net_1 ), .B(N_639), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_64_net_1 ));
    SLE_IP_CLK 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/FF_25  
        (.CLK(VCC), .IPCLKn(AFLSDF_INV_12_net_1));
    INV_BA AFLSDF_INV_49 (.A(AFLSDF_INV_49_net_1), .Y(
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/A_BLK_net[2] )
        );
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_120_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB12_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_6__1_sqmuxa ), .ALn(
        AFLSDF_INV_13_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(GND)
        , .Q(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_120_set_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_197_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_45_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_197_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_197_rs_net_1 ));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_76_set_RNIRUK01  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_76_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_198_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_9_rs[4] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_9_[4]_net_1 ));
    CFG3 #( .INIT(8'h80) )  
        \CoreGPIO_0/xhdl1.GEN_BITS[0].APB_8.GPOUT_reg35_0_a2  (.A(
        N_639), .B(\CoreAPB3_0.u_mux_p_to_b3.PRDATA_0_iv_0_a2_3_5[1] ), 
        .C(N_638), .Y(\CoreGPIO_0/GPOUT_reg35 ));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_11_[0]  (.D(
        \CoreAPB3_0_APBmslave5_PWDATA[0] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB6_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_11__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_182_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_11_rs[0] ));
    CFG2_IP_BC 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/CFG_8  
        (.B(\CoreAPB3_0_APBmslave5_PWDATA[2] ), .C(GND), .IPB(
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/A_DIN_net[2] )
        , .IPC(
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/A_ADDR_net[4] )
        );
    CFG2_IP_BC 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/CFG_22  
        (.B(\CoreAPB3_0_APBmslave5_PWDATA[13] ), .C(
        \COREAPBLSRAM_0/wen ), .IPB(
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/A_DIN_net[14] )
        , .IPC(
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/B_WEN_net[0] )
        );
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_131_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_127_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_131_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_131_rs_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_194_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_74_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_194_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_194_rs_net_1 ));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_82  (.A(
        VCC), .B(VCC), .C(VCC), .IPA(), .IPB(
        \hello_regs_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[23] ), 
        .IPC());
    SLE_IP_EN 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/FF_20  
        (.EN(VCC), .IPENn());
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_data_out8_33  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_2_[4]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_642 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_33_net_1 ));
    SLE \COREAPBLSRAM_0/PREADY_reg  (.D(
        \COREAPBLSRAM_0/PREADY_reg6_i_0 ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB8_rgbr_net_1 ), .EN(VCC), .ALn(
        \hello_regs_MSS_0/MSS_ADLIB_INST_RNIUO3B/U0_RGB1_RGB0_rgbr_net_1 )
        , .ADn(GND), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        CoreAPB3_0_APBmslave7_PREADY));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_14_set_RNIC4GM  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_14_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_189_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_5_rs[1] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_5_[1]_net_1 ));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_272  (
        .A(GND), .B(GND), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_ARLEN_HBURST1_net[0] ), 
        .IPB(\hello_regs_MSS_0/MSS_ADLIB_INST/F_RMW_AXI_net ), .IPC());
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_data_out8_67  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_4_[5]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_648 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_67_net_1 ));
    CFG3 #( .INIT(8'hF2) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_192  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_9_[1]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_643 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_192_i ));
    MSS_010_IP #( .INIT(1438'h00000000003612000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000F00000000F000000000000000000000000000000007FFFFFFFB000001007C33C000000006092C0104003FFFFE400000000000010000000000F81C000001FEDFDC010842108421000001FE34001FF8000000400000000020091007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF)
        , .ACT_UBITS(56'hFFFFFFFFFFFFFF), .MEMORYFILE("ENVM_init.mem")
        , .RTC_MAIN_XTL_FREQ(0.0), .RTC_MAIN_XTL_MODE("") )  
        \hello_regs_MSS_0/MSS_ADLIB_INST/INST_MSS_010_IP  (
        .CAN_RXBUS_MGPIO3A_H2F_A(), .CAN_RXBUS_MGPIO3A_H2F_B(), 
        .CAN_TX_EBL_MGPIO4A_H2F_A(), .CAN_TX_EBL_MGPIO4A_H2F_B(), 
        .CAN_TXBUS_MGPIO2A_H2F_A(), .CAN_TXBUS_MGPIO2A_H2F_B(), 
        .CLK_CONFIG_APB(), .COMMS_INT(), .CONFIG_PRESET_N(), 
        .EDAC_ERROR({nc0, nc1, nc2, nc3, nc4, nc5, nc6, nc7}), 
        .F_FM0_RDATA({nc8, nc9, nc10, nc11, nc12, nc13, nc14, nc15, 
        nc16, nc17, nc18, nc19, nc20, nc21, nc22, nc23, nc24, nc25, 
        nc26, nc27, nc28, nc29, nc30, nc31, nc32, nc33, nc34, nc35, 
        nc36, nc37, nc38, nc39}), .F_FM0_READYOUT(), .F_FM0_RESP(), 
        .F_HM0_ADDR({nc40, nc41, nc42, nc43, nc44, nc45, nc46, nc47, 
        nc48, nc49, nc50, nc51, 
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PADDR[19] , 
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PADDR[18] , 
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PADDR[17] , 
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PADDR[16] , nc52, nc53, 
        nc54, nc55, nc56, nc57, nc58, \CoreAPB3_0_APBmslave5_PADDR[8] , 
        \CoreAPB3_0_APBmslave5_PADDR[7] , 
        \CoreAPB3_0_APBmslave5_PADDR[6] , 
        \CoreAPB3_0_APBmslave5_PADDR[5] , 
        \CoreAPB3_0_APBmslave5_PADDR[4] , 
        \CoreAPB3_0_APBmslave5_PADDR[3] , 
        \CoreAPB3_0_APBmslave5_PADDR[2] , 
        \CoreAPB3_0_APBmslave5_PADDR[1] , 
        \CoreAPB3_0_APBmslave5_PADDR[0] }), .F_HM0_ENABLE(
        CoreAPB3_0_APBmslave5_PENABLE), .F_HM0_SEL(
        hello_regs_MSS_0_FIC_0_APB_MASTER_PSELx), .F_HM0_SIZE({nc59, 
        nc60}), .F_HM0_TRANS1(), .F_HM0_WDATA({
        \CoreAPB3_0_APBmslave5_PWDATA[31] , 
        \CoreAPB3_0_APBmslave5_PWDATA[30] , 
        \CoreAPB3_0_APBmslave5_PWDATA[29] , 
        \CoreAPB3_0_APBmslave5_PWDATA[28] , 
        \CoreAPB3_0_APBmslave5_PWDATA[27] , 
        \CoreAPB3_0_APBmslave5_PWDATA[26] , 
        \CoreAPB3_0_APBmslave5_PWDATA[25] , 
        \CoreAPB3_0_APBmslave5_PWDATA[24] , 
        \CoreAPB3_0_APBmslave5_PWDATA[23] , 
        \CoreAPB3_0_APBmslave5_PWDATA[22] , 
        \CoreAPB3_0_APBmslave5_PWDATA[21] , 
        \CoreAPB3_0_APBmslave5_PWDATA[20] , 
        \CoreAPB3_0_APBmslave5_PWDATA[19] , 
        \CoreAPB3_0_APBmslave5_PWDATA[18] , 
        \CoreAPB3_0_APBmslave5_PWDATA[17] , 
        \CoreAPB3_0_APBmslave5_PWDATA[16] , 
        \CoreAPB3_0_APBmslave5_PWDATA[15] , 
        \CoreAPB3_0_APBmslave5_PWDATA[14] , 
        \CoreAPB3_0_APBmslave5_PWDATA[13] , 
        \CoreAPB3_0_APBmslave5_PWDATA[12] , 
        \CoreAPB3_0_APBmslave5_PWDATA[11] , 
        \CoreAPB3_0_APBmslave5_PWDATA[10] , 
        \CoreAPB3_0_APBmslave5_PWDATA[9] , 
        \CoreAPB3_0_APBmslave5_PWDATA[8] , 
        \CoreAPB3_0_APBmslave5_PWDATA[7] , 
        \CoreAPB3_0_APBmslave5_PWDATA[6] , 
        \CoreAPB3_0_APBmslave5_PWDATA[5] , 
        \CoreAPB3_0_APBmslave5_PWDATA[4] , 
        \CoreAPB3_0_APBmslave5_PWDATA[3] , 
        \CoreAPB3_0_APBmslave5_PWDATA[2] , 
        \CoreAPB3_0_APBmslave5_PWDATA[1] , 
        \CoreAPB3_0_APBmslave5_PWDATA[0] }), .F_HM0_WRITE(
        CoreAPB3_0_APBmslave5_PWRITE), .FAB_CHRGVBUS(), 
        .FAB_DISCHRGVBUS(), .FAB_DMPULLDOWN(), .FAB_DPPULLDOWN(), 
        .FAB_DRVVBUS(), .FAB_IDPULLUP(), .FAB_OPMODE({nc61, nc62}), 
        .FAB_SUSPENDM(), .FAB_TERMSEL(), .FAB_TXVALID(), .FAB_VCONTROL({
        nc63, nc64, nc65, nc66}), .FAB_VCONTROLLOADM(), .FAB_XCVRSEL({
        nc67, nc68}), .FAB_XDATAOUT({nc69, nc70, nc71, nc72, nc73, 
        nc74, nc75, nc76}), .FACC_GLMUX_SEL(), .FIC32_0_MASTER({nc77, 
        nc78}), .FIC32_1_MASTER({nc79, nc80}), .FPGA_RESET_N(
        \hello_regs_MSS_0/FPGA_RESET_N ), .GTX_CLK(), .H2F_INTERRUPT({
        nc81, nc82, nc83, nc84, nc85, nc86, nc87, nc88, nc89, nc90, 
        nc91, nc92, nc93, nc94, nc95, nc96}), .H2F_NMI(), .H2FCALIB(), 
        .I2C0_SCL_MGPIO31B_H2F_A(), .I2C0_SCL_MGPIO31B_H2F_B(), 
        .I2C0_SDA_MGPIO30B_H2F_A(), .I2C0_SDA_MGPIO30B_H2F_B(), 
        .I2C1_SCL_MGPIO1A_H2F_A(), .I2C1_SCL_MGPIO1A_H2F_B(), 
        .I2C1_SDA_MGPIO0A_H2F_A(), .I2C1_SDA_MGPIO0A_H2F_B(), .MDCF(), 
        .MDOENF(), .MDOF(), .MMUART0_CTS_MGPIO19B_H2F_A(), 
        .MMUART0_CTS_MGPIO19B_H2F_B(), .MMUART0_DCD_MGPIO22B_H2F_A(), 
        .MMUART0_DCD_MGPIO22B_H2F_B(), .MMUART0_DSR_MGPIO20B_H2F_A(), 
        .MMUART0_DSR_MGPIO20B_H2F_B(), .MMUART0_DTR_MGPIO18B_H2F_A(), 
        .MMUART0_DTR_MGPIO18B_H2F_B(), .MMUART0_RI_MGPIO21B_H2F_A(), 
        .MMUART0_RI_MGPIO21B_H2F_B(), .MMUART0_RTS_MGPIO17B_H2F_A(), 
        .MMUART0_RTS_MGPIO17B_H2F_B(), .MMUART0_RXD_MGPIO28B_H2F_A(), 
        .MMUART0_RXD_MGPIO28B_H2F_B(), .MMUART0_SCK_MGPIO29B_H2F_A(), 
        .MMUART0_SCK_MGPIO29B_H2F_B(), .MMUART0_TXD_MGPIO27B_H2F_A(), 
        .MMUART0_TXD_MGPIO27B_H2F_B(), .MMUART1_DTR_MGPIO12B_H2F_A(), 
        .MMUART1_RTS_MGPIO11B_H2F_A(), .MMUART1_RTS_MGPIO11B_H2F_B(), 
        .MMUART1_RXD_MGPIO26B_H2F_A(), .MMUART1_RXD_MGPIO26B_H2F_B(), 
        .MMUART1_SCK_MGPIO25B_H2F_A(), .MMUART1_SCK_MGPIO25B_H2F_B(), 
        .MMUART1_TXD_MGPIO24B_H2F_A(), .MMUART1_TXD_MGPIO24B_H2F_B(), 
        .MPLL_LOCK(), .PER2_FABRIC_PADDR({nc97, nc98, nc99, nc100, 
        nc101, nc102, nc103, nc104, nc105, nc106, nc107, nc108, nc109, 
        nc110}), .PER2_FABRIC_PENABLE(), .PER2_FABRIC_PSEL(), 
        .PER2_FABRIC_PWDATA({nc111, nc112, nc113, nc114, nc115, nc116, 
        nc117, nc118, nc119, nc120, nc121, nc122, nc123, nc124, nc125, 
        nc126, nc127, nc128, nc129, nc130, nc131, nc132, nc133, nc134, 
        nc135, nc136, nc137, nc138, nc139, nc140, nc141, nc142}), 
        .PER2_FABRIC_PWRITE(), .RTC_MATCH(), .SLEEPDEEP(), 
        .SLEEPHOLDACK(), .SLEEPING(), .SMBALERT_NO0(), .SMBALERT_NO1(), 
        .SMBSUS_NO0(), .SMBSUS_NO1(), .SPI0_CLK_OUT(), 
        .SPI0_SDI_MGPIO5A_H2F_A(), .SPI0_SDI_MGPIO5A_H2F_B(), 
        .SPI0_SDO_MGPIO6A_H2F_A(), .SPI0_SDO_MGPIO6A_H2F_B(), 
        .SPI0_SS0_MGPIO7A_H2F_A(), .SPI0_SS0_MGPIO7A_H2F_B(), 
        .SPI0_SS1_MGPIO8A_H2F_A(), .SPI0_SS1_MGPIO8A_H2F_B(), 
        .SPI0_SS2_MGPIO9A_H2F_A(), .SPI0_SS2_MGPIO9A_H2F_B(), 
        .SPI0_SS3_MGPIO10A_H2F_A(), .SPI0_SS3_MGPIO10A_H2F_B(), 
        .SPI0_SS4_MGPIO19A_H2F_A(), .SPI0_SS5_MGPIO20A_H2F_A(), 
        .SPI0_SS6_MGPIO21A_H2F_A(), .SPI0_SS7_MGPIO22A_H2F_A(), 
        .SPI1_CLK_OUT(), .SPI1_SDI_MGPIO11A_H2F_A(), 
        .SPI1_SDI_MGPIO11A_H2F_B(), .SPI1_SDO_MGPIO12A_H2F_A(), 
        .SPI1_SDO_MGPIO12A_H2F_B(), .SPI1_SS0_MGPIO13A_H2F_A(), 
        .SPI1_SS0_MGPIO13A_H2F_B(), .SPI1_SS1_MGPIO14A_H2F_A(), 
        .SPI1_SS1_MGPIO14A_H2F_B(), .SPI1_SS2_MGPIO15A_H2F_A(), 
        .SPI1_SS2_MGPIO15A_H2F_B(), .SPI1_SS3_MGPIO16A_H2F_A(), 
        .SPI1_SS3_MGPIO16A_H2F_B(), .SPI1_SS4_MGPIO17A_H2F_A(), 
        .SPI1_SS5_MGPIO18A_H2F_A(), .SPI1_SS6_MGPIO23A_H2F_A(), 
        .SPI1_SS7_MGPIO24A_H2F_A(), .TCGF({nc143, nc144, nc145, nc146, 
        nc147, nc148, nc149, nc150, nc151, nc152}), .TRACECLK(), 
        .TRACEDATA({nc153, nc154, nc155, nc156}), .TX_CLK(), .TX_ENF(), 
        .TX_ERRF(), .TXCTL_EN_RIF(), .TXD_RIF({nc157, nc158, nc159, 
        nc160}), .TXDF({nc161, nc162, nc163, nc164, nc165, nc166, 
        nc167, nc168}), .TXEV(), .WDOGTIMEOUT(), .F_ARREADY_HREADYOUT1(
        ), .F_AWREADY_HREADYOUT0(), .F_BID({nc169, nc170, nc171, nc172})
        , .F_BRESP_HRESP0({nc173, nc174}), .F_BVALID(), 
        .F_RDATA_HRDATA01({nc175, nc176, nc177, nc178, nc179, nc180, 
        nc181, nc182, nc183, nc184, nc185, nc186, nc187, nc188, nc189, 
        nc190, nc191, nc192, nc193, nc194, nc195, nc196, nc197, nc198, 
        nc199, nc200, nc201, nc202, nc203, nc204, nc205, nc206, nc207, 
        nc208, nc209, nc210, nc211, nc212, nc213, nc214, nc215, nc216, 
        nc217, nc218, nc219, nc220, nc221, nc222, nc223, nc224, nc225, 
        nc226, nc227, nc228, nc229, nc230, nc231, nc232, nc233, nc234, 
        nc235, nc236, nc237, nc238}), .F_RID({nc239, nc240, nc241, 
        nc242}), .F_RLAST(), .F_RRESP_HRESP1({nc243, nc244}), 
        .F_RVALID(), .F_WREADY(), .MDDR_FABRIC_PRDATA({nc245, nc246, 
        nc247, nc248, nc249, nc250, nc251, nc252, nc253, nc254, nc255, 
        nc256, nc257, nc258, nc259, nc260}), .MDDR_FABRIC_PREADY(), 
        .MDDR_FABRIC_PSLVERR(), .CAN_RXBUS_F2H_SCP(
        \hello_regs_MSS_0/MSS_ADLIB_INST/CAN_RXBUS_F2H_SCP_net ), 
        .CAN_TX_EBL_F2H_SCP(
        \hello_regs_MSS_0/MSS_ADLIB_INST/CAN_TX_EBL_F2H_SCP_net ), 
        .CAN_TXBUS_F2H_SCP(
        \hello_regs_MSS_0/MSS_ADLIB_INST/CAN_TXBUS_F2H_SCP_net ), 
        .COLF(\hello_regs_MSS_0/MSS_ADLIB_INST/COLF_net ), .CRSF(
        \hello_regs_MSS_0/MSS_ADLIB_INST/CRSF_net ), .F2_DMAREADY({
        \hello_regs_MSS_0/MSS_ADLIB_INST/F2_DMAREADY_net[1] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F2_DMAREADY_net[0] }), 
        .F2H_INTERRUPT({
        \hello_regs_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[15] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[14] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[13] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[12] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[11] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[10] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[9] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[8] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[7] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[6] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[5] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[4] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[3] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[2] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[1] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[0] }), 
        .F2HCALIB(\hello_regs_MSS_0/MSS_ADLIB_INST/F2HCALIB_net ), 
        .F_DMAREADY({
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_DMAREADY_net[1] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_DMAREADY_net[0] }), 
        .F_FM0_ADDR({
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[31] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[30] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[29] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[28] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[27] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[26] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[25] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[24] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[23] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[22] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[21] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[20] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[19] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[18] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[17] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[16] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[15] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[14] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[13] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[12] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[11] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[10] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[9] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[8] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[7] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[6] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[5] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[4] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[3] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[2] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[1] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[0] }), 
        .F_FM0_ENABLE(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_ENABLE_net ), 
        .F_FM0_MASTLOCK(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_MASTLOCK_net ), 
        .F_FM0_READY(\hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_READY_net )
        , .F_FM0_SEL(\hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_SEL_net ), 
        .F_FM0_SIZE({
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_SIZE_net[1] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_SIZE_net[0] }), 
        .F_FM0_TRANS1(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_TRANS1_net ), 
        .F_FM0_WDATA({
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[31] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[30] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[29] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[28] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[27] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[26] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[25] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[24] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[23] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[22] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[21] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[20] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[19] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[18] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[17] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[16] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[15] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[14] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[13] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[12] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[11] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[10] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[9] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[8] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[7] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[6] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[5] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[4] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[3] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[2] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[1] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[0] }), 
        .F_FM0_WRITE(\hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_WRITE_net )
        , .F_HM0_RDATA({
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[31] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[30] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[29] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[28] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[27] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[26] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[25] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[24] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[23] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[22] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[21] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[20] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[19] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[18] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[17] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[16] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[15] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[14] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[13] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[12] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[11] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[10] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[9] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[8] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[7] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[6] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[5] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[4] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[3] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[2] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[1] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[0] }), 
        .F_HM0_READY(\hello_regs_MSS_0/MSS_ADLIB_INST/F_HM0_READY_net )
        , .F_HM0_RESP(\hello_regs_MSS_0/MSS_ADLIB_INST/F_HM0_RESP_net )
        , .FAB_AVALID(\hello_regs_MSS_0/MSS_ADLIB_INST/FAB_AVALID_net )
        , .FAB_HOSTDISCON(
        \hello_regs_MSS_0/MSS_ADLIB_INST/FAB_HOSTDISCON_net ), 
        .FAB_IDDIG(\hello_regs_MSS_0/MSS_ADLIB_INST/FAB_IDDIG_net ), 
        .FAB_LINESTATE({
        \hello_regs_MSS_0/MSS_ADLIB_INST/FAB_LINESTATE_net[1] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/FAB_LINESTATE_net[0] }), 
        .FAB_M3_RESET_N(
        \hello_regs_MSS_0/MSS_ADLIB_INST/FAB_M3_RESET_N_net ), 
        .FAB_PLL_LOCK(
        \hello_regs_MSS_0/MSS_ADLIB_INST/FAB_PLL_LOCK_net ), 
        .FAB_RXACTIVE(
        \hello_regs_MSS_0/MSS_ADLIB_INST/FAB_RXACTIVE_net ), 
        .FAB_RXERROR(\hello_regs_MSS_0/MSS_ADLIB_INST/FAB_RXERROR_net )
        , .FAB_RXVALID(
        \hello_regs_MSS_0/MSS_ADLIB_INST/FAB_RXVALID_net ), 
        .FAB_RXVALIDH(
        \hello_regs_MSS_0/MSS_ADLIB_INST/FAB_RXVALIDH_net ), 
        .FAB_SESSEND(\hello_regs_MSS_0/MSS_ADLIB_INST/FAB_SESSEND_net )
        , .FAB_TXREADY(
        \hello_regs_MSS_0/MSS_ADLIB_INST/FAB_TXREADY_net ), 
        .FAB_VBUSVALID(
        \hello_regs_MSS_0/MSS_ADLIB_INST/FAB_VBUSVALID_net ), 
        .FAB_VSTATUS({
        \hello_regs_MSS_0/MSS_ADLIB_INST/FAB_VSTATUS_net[7] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/FAB_VSTATUS_net[6] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/FAB_VSTATUS_net[5] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/FAB_VSTATUS_net[4] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/FAB_VSTATUS_net[3] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/FAB_VSTATUS_net[2] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/FAB_VSTATUS_net[1] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/FAB_VSTATUS_net[0] }), 
        .FAB_XDATAIN({
        \hello_regs_MSS_0/MSS_ADLIB_INST/FAB_XDATAIN_net[7] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/FAB_XDATAIN_net[6] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/FAB_XDATAIN_net[5] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/FAB_XDATAIN_net[4] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/FAB_XDATAIN_net[3] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/FAB_XDATAIN_net[2] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/FAB_XDATAIN_net[1] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/FAB_XDATAIN_net[0] }), 
        .GTX_CLKPF(\hello_regs_MSS_0/MSS_ADLIB_INST/GTX_CLKPF_net ), 
        .I2C0_BCLK(\hello_regs_MSS_0/MSS_ADLIB_INST/I2C0_BCLK_net ), 
        .I2C0_SCL_F2H_SCP(
        \hello_regs_MSS_0/MSS_ADLIB_INST/I2C0_SCL_F2H_SCP_net ), 
        .I2C0_SDA_F2H_SCP(
        \hello_regs_MSS_0/MSS_ADLIB_INST/I2C0_SDA_F2H_SCP_net ), 
        .I2C1_BCLK(\hello_regs_MSS_0/MSS_ADLIB_INST/I2C1_BCLK_net ), 
        .I2C1_SCL_F2H_SCP(
        \hello_regs_MSS_0/MSS_ADLIB_INST/I2C1_SCL_F2H_SCP_net ), 
        .I2C1_SDA_F2H_SCP(
        \hello_regs_MSS_0/MSS_ADLIB_INST/I2C1_SDA_F2H_SCP_net ), .MDIF(
        \hello_regs_MSS_0/MSS_ADLIB_INST/MDIF_net ), .MGPIO0A_F2H_GPIN(
        \hello_regs_MSS_0/MSS_ADLIB_INST/MGPIO0A_F2H_GPIN_net ), 
        .MGPIO10A_F2H_GPIN(
        \hello_regs_MSS_0/MSS_ADLIB_INST/MGPIO10A_F2H_GPIN_net ), 
        .MGPIO11A_F2H_GPIN(
        \hello_regs_MSS_0/MSS_ADLIB_INST/MGPIO11A_F2H_GPIN_net ), 
        .MGPIO11B_F2H_GPIN(
        \hello_regs_MSS_0/MSS_ADLIB_INST/MGPIO11B_F2H_GPIN_net ), 
        .MGPIO12A_F2H_GPIN(
        \hello_regs_MSS_0/MSS_ADLIB_INST/MGPIO12A_F2H_GPIN_net ), 
        .MGPIO13A_F2H_GPIN(
        \hello_regs_MSS_0/MSS_ADLIB_INST/MGPIO13A_F2H_GPIN_net ), 
        .MGPIO14A_F2H_GPIN(
        \hello_regs_MSS_0/MSS_ADLIB_INST/MGPIO14A_F2H_GPIN_net ), 
        .MGPIO15A_F2H_GPIN(
        \hello_regs_MSS_0/MSS_ADLIB_INST/MGPIO15A_F2H_GPIN_net ), 
        .MGPIO16A_F2H_GPIN(
        \hello_regs_MSS_0/MSS_ADLIB_INST/MGPIO16A_F2H_GPIN_net ), 
        .MGPIO17B_F2H_GPIN(
        \hello_regs_MSS_0/MSS_ADLIB_INST/MGPIO17B_F2H_GPIN_net ), 
        .MGPIO18B_F2H_GPIN(
        \hello_regs_MSS_0/MSS_ADLIB_INST/MGPIO18B_F2H_GPIN_net ), 
        .MGPIO19B_F2H_GPIN(
        \hello_regs_MSS_0/MSS_ADLIB_INST/MGPIO19B_F2H_GPIN_net ), 
        .MGPIO1A_F2H_GPIN(
        \hello_regs_MSS_0/MSS_ADLIB_INST/MGPIO1A_F2H_GPIN_net ), 
        .MGPIO20B_F2H_GPIN(
        \hello_regs_MSS_0/MSS_ADLIB_INST/MGPIO20B_F2H_GPIN_net ), 
        .MGPIO21B_F2H_GPIN(
        \hello_regs_MSS_0/MSS_ADLIB_INST/MGPIO21B_F2H_GPIN_net ), 
        .MGPIO22B_F2H_GPIN(
        \hello_regs_MSS_0/MSS_ADLIB_INST/MGPIO22B_F2H_GPIN_net ), 
        .MGPIO24B_F2H_GPIN(
        \hello_regs_MSS_0/MSS_ADLIB_INST/MGPIO24B_F2H_GPIN_net ), 
        .MGPIO25B_F2H_GPIN(
        \hello_regs_MSS_0/MSS_ADLIB_INST/MGPIO25B_F2H_GPIN_net ), 
        .MGPIO26B_F2H_GPIN(
        \hello_regs_MSS_0/MSS_ADLIB_INST/MGPIO26B_F2H_GPIN_net ), 
        .MGPIO27B_F2H_GPIN(
        \hello_regs_MSS_0/MSS_ADLIB_INST/MGPIO27B_F2H_GPIN_net ), 
        .MGPIO28B_F2H_GPIN(
        \hello_regs_MSS_0/MSS_ADLIB_INST/MGPIO28B_F2H_GPIN_net ), 
        .MGPIO29B_F2H_GPIN(
        \hello_regs_MSS_0/MSS_ADLIB_INST/MGPIO29B_F2H_GPIN_net ), 
        .MGPIO2A_F2H_GPIN(
        \hello_regs_MSS_0/MSS_ADLIB_INST/MGPIO2A_F2H_GPIN_net ), 
        .MGPIO30B_F2H_GPIN(
        \hello_regs_MSS_0/MSS_ADLIB_INST/MGPIO30B_F2H_GPIN_net ), 
        .MGPIO31B_F2H_GPIN(
        \hello_regs_MSS_0/MSS_ADLIB_INST/MGPIO31B_F2H_GPIN_net ), 
        .MGPIO3A_F2H_GPIN(
        \hello_regs_MSS_0/MSS_ADLIB_INST/MGPIO3A_F2H_GPIN_net ), 
        .MGPIO4A_F2H_GPIN(
        \hello_regs_MSS_0/MSS_ADLIB_INST/MGPIO4A_F2H_GPIN_net ), 
        .MGPIO5A_F2H_GPIN(
        \hello_regs_MSS_0/MSS_ADLIB_INST/MGPIO5A_F2H_GPIN_net ), 
        .MGPIO6A_F2H_GPIN(
        \hello_regs_MSS_0/MSS_ADLIB_INST/MGPIO6A_F2H_GPIN_net ), 
        .MGPIO7A_F2H_GPIN(
        \hello_regs_MSS_0/MSS_ADLIB_INST/MGPIO7A_F2H_GPIN_net ), 
        .MGPIO8A_F2H_GPIN(
        \hello_regs_MSS_0/MSS_ADLIB_INST/MGPIO8A_F2H_GPIN_net ), 
        .MGPIO9A_F2H_GPIN(
        \hello_regs_MSS_0/MSS_ADLIB_INST/MGPIO9A_F2H_GPIN_net ), 
        .MMUART0_CTS_F2H_SCP(
        \hello_regs_MSS_0/MSS_ADLIB_INST/MMUART0_CTS_F2H_SCP_net ), 
        .MMUART0_DCD_F2H_SCP(
        \hello_regs_MSS_0/MSS_ADLIB_INST/MMUART0_DCD_F2H_SCP_net ), 
        .MMUART0_DSR_F2H_SCP(
        \hello_regs_MSS_0/MSS_ADLIB_INST/MMUART0_DSR_F2H_SCP_net ), 
        .MMUART0_DTR_F2H_SCP(
        \hello_regs_MSS_0/MSS_ADLIB_INST/MMUART0_DTR_F2H_SCP_net ), 
        .MMUART0_RI_F2H_SCP(
        \hello_regs_MSS_0/MSS_ADLIB_INST/MMUART0_RI_F2H_SCP_net ), 
        .MMUART0_RTS_F2H_SCP(
        \hello_regs_MSS_0/MSS_ADLIB_INST/MMUART0_RTS_F2H_SCP_net ), 
        .MMUART0_RXD_F2H_SCP(
        \hello_regs_MSS_0/MSS_ADLIB_INST/MMUART0_RXD_F2H_SCP_net ), 
        .MMUART0_SCK_F2H_SCP(
        \hello_regs_MSS_0/MSS_ADLIB_INST/MMUART0_SCK_F2H_SCP_net ), 
        .MMUART0_TXD_F2H_SCP(
        \hello_regs_MSS_0/MSS_ADLIB_INST/MMUART0_TXD_F2H_SCP_net ), 
        .MMUART1_CTS_F2H_SCP(
        \hello_regs_MSS_0/MSS_ADLIB_INST/MMUART1_CTS_F2H_SCP_net ), 
        .MMUART1_DCD_F2H_SCP(
        \hello_regs_MSS_0/MSS_ADLIB_INST/MMUART1_DCD_F2H_SCP_net ), 
        .MMUART1_DSR_F2H_SCP(
        \hello_regs_MSS_0/MSS_ADLIB_INST/MMUART1_DSR_F2H_SCP_net ), 
        .MMUART1_RI_F2H_SCP(
        \hello_regs_MSS_0/MSS_ADLIB_INST/MMUART1_RI_F2H_SCP_net ), 
        .MMUART1_RTS_F2H_SCP(
        \hello_regs_MSS_0/MSS_ADLIB_INST/MMUART1_RTS_F2H_SCP_net ), 
        .MMUART1_RXD_F2H_SCP(
        \hello_regs_MSS_0/MSS_ADLIB_INST/MMUART1_RXD_F2H_SCP_net ), 
        .MMUART1_SCK_F2H_SCP(
        \hello_regs_MSS_0/MSS_ADLIB_INST/MMUART1_SCK_F2H_SCP_net ), 
        .MMUART1_TXD_F2H_SCP(
        \hello_regs_MSS_0/MSS_ADLIB_INST/MMUART1_TXD_F2H_SCP_net ), 
        .PER2_FABRIC_PRDATA({
        \hello_regs_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[31] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[30] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[29] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[28] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[27] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[26] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[25] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[24] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[23] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[22] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[21] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[20] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[19] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[18] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[17] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[16] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[15] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[14] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[13] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[12] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[11] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[10] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[9] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[8] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[7] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[6] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[5] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[4] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[3] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[2] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[1] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[0] }), 
        .PER2_FABRIC_PREADY(
        \hello_regs_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PREADY_net ), 
        .PER2_FABRIC_PSLVERR(
        \hello_regs_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PSLVERR_net ), 
        .RCGF({\hello_regs_MSS_0/MSS_ADLIB_INST/RCGF_net[9] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/RCGF_net[8] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/RCGF_net[7] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/RCGF_net[6] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/RCGF_net[5] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/RCGF_net[4] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/RCGF_net[3] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/RCGF_net[2] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/RCGF_net[1] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/RCGF_net[0] }), .RX_CLKPF(
        \hello_regs_MSS_0/MSS_ADLIB_INST/RX_CLKPF_net ), .RX_DVF(
        \hello_regs_MSS_0/MSS_ADLIB_INST/RX_DVF_net ), .RX_ERRF(
        \hello_regs_MSS_0/MSS_ADLIB_INST/RX_ERRF_net ), .RX_EV(
        \hello_regs_MSS_0/MSS_ADLIB_INST/RX_EV_net ), .RXDF({
        \hello_regs_MSS_0/MSS_ADLIB_INST/RXDF_net[7] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/RXDF_net[6] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/RXDF_net[5] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/RXDF_net[4] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/RXDF_net[3] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/RXDF_net[2] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/RXDF_net[1] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/RXDF_net[0] }), .SLEEPHOLDREQ(
        \hello_regs_MSS_0/MSS_ADLIB_INST/SLEEPHOLDREQ_net ), 
        .SMBALERT_NI0(
        \hello_regs_MSS_0/MSS_ADLIB_INST/SMBALERT_NI0_net ), 
        .SMBALERT_NI1(
        \hello_regs_MSS_0/MSS_ADLIB_INST/SMBALERT_NI1_net ), 
        .SMBSUS_NI0(\hello_regs_MSS_0/MSS_ADLIB_INST/SMBSUS_NI0_net ), 
        .SMBSUS_NI1(\hello_regs_MSS_0/MSS_ADLIB_INST/SMBSUS_NI1_net ), 
        .SPI0_CLK_IN(\hello_regs_MSS_0/MSS_ADLIB_INST/SPI0_CLK_IN_net )
        , .SPI0_SDI_F2H_SCP(
        \hello_regs_MSS_0/MSS_ADLIB_INST/SPI0_SDI_F2H_SCP_net ), 
        .SPI0_SDO_F2H_SCP(
        \hello_regs_MSS_0/MSS_ADLIB_INST/SPI0_SDO_F2H_SCP_net ), 
        .SPI0_SS0_F2H_SCP(
        \hello_regs_MSS_0/MSS_ADLIB_INST/SPI0_SS0_F2H_SCP_net ), 
        .SPI0_SS1_F2H_SCP(
        \hello_regs_MSS_0/MSS_ADLIB_INST/SPI0_SS1_F2H_SCP_net ), 
        .SPI0_SS2_F2H_SCP(
        \hello_regs_MSS_0/MSS_ADLIB_INST/SPI0_SS2_F2H_SCP_net ), 
        .SPI0_SS3_F2H_SCP(
        \hello_regs_MSS_0/MSS_ADLIB_INST/SPI0_SS3_F2H_SCP_net ), 
        .SPI1_CLK_IN(\hello_regs_MSS_0/MSS_ADLIB_INST/SPI1_CLK_IN_net )
        , .SPI1_SDI_F2H_SCP(
        \hello_regs_MSS_0/MSS_ADLIB_INST/SPI1_SDI_F2H_SCP_net ), 
        .SPI1_SDO_F2H_SCP(
        \hello_regs_MSS_0/MSS_ADLIB_INST/SPI1_SDO_F2H_SCP_net ), 
        .SPI1_SS0_F2H_SCP(
        \hello_regs_MSS_0/MSS_ADLIB_INST/SPI1_SS0_F2H_SCP_net ), 
        .SPI1_SS1_F2H_SCP(
        \hello_regs_MSS_0/MSS_ADLIB_INST/SPI1_SS1_F2H_SCP_net ), 
        .SPI1_SS2_F2H_SCP(
        \hello_regs_MSS_0/MSS_ADLIB_INST/SPI1_SS2_F2H_SCP_net ), 
        .SPI1_SS3_F2H_SCP(
        \hello_regs_MSS_0/MSS_ADLIB_INST/SPI1_SS3_F2H_SCP_net ), 
        .TX_CLKPF(\hello_regs_MSS_0/MSS_ADLIB_INST/TX_CLKPF_net ), 
        .USER_MSS_GPIO_RESET_N(
        \hello_regs_MSS_0/MSS_ADLIB_INST/USER_MSS_GPIO_RESET_N_net ), 
        .USER_MSS_RESET_N(
        \hello_regs_MSS_0/MSS_ADLIB_INST/USER_MSS_RESET_N_net ), 
        .XCLK_FAB(\hello_regs_MSS_0/MSS_ADLIB_INST/XCLK_FAB_net ), 
        .CLK_BASE(\hello_regs_MSS_0/MSS_ADLIB_INST/CLK_BASE_net ), 
        .CLK_MDDR_APB(
        \hello_regs_MSS_0/MSS_ADLIB_INST/CLK_MDDR_APB_net ), 
        .F_ARADDR_HADDR1({
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[31] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[30] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[29] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[28] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[27] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[26] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[25] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[24] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[23] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[22] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[21] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[20] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[19] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[18] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[17] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[16] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[15] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[14] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[13] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[12] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[11] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[10] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[9] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[8] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[7] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[6] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[5] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[4] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[3] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[2] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[1] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[0] }), 
        .F_ARBURST_HTRANS1({
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_ARBURST_HTRANS1_net[1] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_ARBURST_HTRANS1_net[0] }), 
        .F_ARID_HSEL1({
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_ARID_HSEL1_net[3] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_ARID_HSEL1_net[2] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_ARID_HSEL1_net[1] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_ARID_HSEL1_net[0] }), 
        .F_ARLEN_HBURST1({
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_ARLEN_HBURST1_net[3] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_ARLEN_HBURST1_net[2] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_ARLEN_HBURST1_net[1] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_ARLEN_HBURST1_net[0] }), 
        .F_ARLOCK_HMASTLOCK1({
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_ARLOCK_HMASTLOCK1_net[1] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_ARLOCK_HMASTLOCK1_net[0] }), 
        .F_ARSIZE_HSIZE1({
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_ARSIZE_HSIZE1_net[1] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_ARSIZE_HSIZE1_net[0] }), 
        .F_ARVALID_HWRITE1(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_ARVALID_HWRITE1_net ), 
        .F_AWADDR_HADDR0({
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[31] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[30] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[29] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[28] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[27] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[26] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[25] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[24] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[23] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[22] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[21] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[20] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[19] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[18] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[17] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[16] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[15] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[14] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[13] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[12] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[11] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[10] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[9] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[8] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[7] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[6] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[5] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[4] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[3] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[2] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[1] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[0] }), 
        .F_AWBURST_HTRANS0({
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_AWBURST_HTRANS0_net[1] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_AWBURST_HTRANS0_net[0] }), 
        .F_AWID_HSEL0({
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_AWID_HSEL0_net[3] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_AWID_HSEL0_net[2] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_AWID_HSEL0_net[1] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_AWID_HSEL0_net[0] }), 
        .F_AWLEN_HBURST0({
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_AWLEN_HBURST0_net[3] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_AWLEN_HBURST0_net[2] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_AWLEN_HBURST0_net[1] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_AWLEN_HBURST0_net[0] }), 
        .F_AWLOCK_HMASTLOCK0({
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_AWLOCK_HMASTLOCK0_net[1] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_AWLOCK_HMASTLOCK0_net[0] }), 
        .F_AWSIZE_HSIZE0({
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_AWSIZE_HSIZE0_net[1] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_AWSIZE_HSIZE0_net[0] }), 
        .F_AWVALID_HWRITE0(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_AWVALID_HWRITE0_net ), 
        .F_BREADY(\hello_regs_MSS_0/MSS_ADLIB_INST/F_BREADY_net ), 
        .F_RMW_AXI(\hello_regs_MSS_0/MSS_ADLIB_INST/F_RMW_AXI_net ), 
        .F_RREADY(\hello_regs_MSS_0/MSS_ADLIB_INST/F_RREADY_net ), 
        .F_WDATA_HWDATA01({
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[63] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[62] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[61] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[60] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[59] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[58] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[57] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[56] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[55] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[54] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[53] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[52] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[51] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[50] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[49] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[48] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[47] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[46] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[45] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[44] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[43] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[42] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[41] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[40] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[39] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[38] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[37] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[36] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[35] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[34] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[33] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[32] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[31] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[30] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[29] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[28] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[27] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[26] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[25] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[24] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[23] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[22] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[21] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[20] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[19] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[18] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[17] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[16] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[15] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[14] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[13] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[12] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[11] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[10] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[9] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[8] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[7] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[6] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[5] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[4] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[3] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[2] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[1] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[0] }), 
        .F_WID_HREADY01({
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WID_HREADY01_net[3] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WID_HREADY01_net[2] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WID_HREADY01_net[1] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WID_HREADY01_net[0] }), 
        .F_WLAST(\hello_regs_MSS_0/MSS_ADLIB_INST/F_WLAST_net ), 
        .F_WSTRB({\hello_regs_MSS_0/MSS_ADLIB_INST/F_WSTRB_net[7] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WSTRB_net[6] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WSTRB_net[5] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WSTRB_net[4] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WSTRB_net[3] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WSTRB_net[2] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WSTRB_net[1] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WSTRB_net[0] }), .F_WVALID(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WVALID_net ), 
        .FPGA_MDDR_ARESET_N(
        \hello_regs_MSS_0/MSS_ADLIB_INST/FPGA_MDDR_ARESET_N_net ), 
        .MDDR_FABRIC_PADDR({
        \hello_regs_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PADDR_net[10] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PADDR_net[9] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PADDR_net[8] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PADDR_net[7] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PADDR_net[6] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PADDR_net[5] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PADDR_net[4] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PADDR_net[3] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PADDR_net[2] }), 
        .MDDR_FABRIC_PENABLE(
        \hello_regs_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PENABLE_net ), 
        .MDDR_FABRIC_PSEL(
        \hello_regs_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PSEL_net ), 
        .MDDR_FABRIC_PWDATA({
        \hello_regs_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[15] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[14] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[13] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[12] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[11] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[10] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[9] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[8] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[7] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[6] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[5] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[4] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[3] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[2] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[1] , 
        \hello_regs_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[0] }), 
        .MDDR_FABRIC_PWRITE(
        \hello_regs_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWRITE_net ), 
        .PRESET_N(\hello_regs_MSS_0/MSS_ADLIB_INST/PRESET_N_net ), 
        .CAN_RXBUS_USBA_DATA1_MGPIO3A_IN(GND), 
        .CAN_TX_EBL_USBA_DATA2_MGPIO4A_IN(GND), 
        .CAN_TXBUS_USBA_DATA0_MGPIO2A_IN(GND), .DM_IN({GND, GND, GND}), 
        .DRAM_DQ_IN({GND, GND, GND, GND, GND, GND, GND, GND, GND, GND, 
        GND, GND, GND, GND, GND, GND, GND, GND}), .DRAM_DQS_IN({GND, 
        GND, GND}), .DRAM_FIFO_WE_IN({GND, GND}), 
        .I2C0_SCL_USBC_DATA1_MGPIO31B_IN(GND), 
        .I2C0_SDA_USBC_DATA0_MGPIO30B_IN(GND), 
        .I2C1_SCL_USBA_DATA4_MGPIO1A_IN(GND), 
        .I2C1_SDA_USBA_DATA3_MGPIO0A_IN(GND), 
        .MMUART0_CTS_USBC_DATA7_MGPIO19B_IN(GND), 
        .MMUART0_DCD_MGPIO22B_IN(GND), .MMUART0_DSR_MGPIO20B_IN(GND), 
        .MMUART0_DTR_USBC_DATA6_MGPIO18B_IN(GND), 
        .MMUART0_RI_MGPIO21B_IN(GND), 
        .MMUART0_RTS_USBC_DATA5_MGPIO17B_IN(GND), 
        .MMUART0_RXD_USBC_STP_MGPIO28B_IN(
        \hello_regs_MSS_0/MMUART_0_RXD_PAD_Y ), 
        .MMUART0_SCK_USBC_NXT_MGPIO29B_IN(GND), 
        .MMUART0_TXD_USBC_DIR_MGPIO27B_IN(GND), 
        .MMUART1_RXD_USBC_DATA3_MGPIO26B_IN(GND), 
        .MMUART1_SCK_USBC_DATA4_MGPIO25B_IN(GND), 
        .MMUART1_TXD_USBC_DATA2_MGPIO24B_IN(GND), 
        .RGMII_GTX_CLK_RMII_CLK_USBB_XCLK_IN(GND), 
        .RGMII_MDC_RMII_MDC_IN(GND), 
        .RGMII_MDIO_RMII_MDIO_USBB_DATA7_IN(GND), .RGMII_RX_CLK_IN(GND)
        , .RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_IN(GND), 
        .RGMII_RXD0_RMII_RXD0_USBB_DATA0_IN(GND), 
        .RGMII_RXD1_RMII_RXD1_USBB_DATA1_IN(GND), 
        .RGMII_RXD2_RMII_RX_ER_USBB_DATA3_IN(GND), 
        .RGMII_RXD3_USBB_DATA4_IN(GND), .RGMII_TX_CLK_IN(GND), 
        .RGMII_TX_CTL_RMII_TX_EN_USBB_NXT_IN(GND), 
        .RGMII_TXD0_RMII_TXD0_USBB_DIR_IN(GND), 
        .RGMII_TXD1_RMII_TXD1_USBB_STP_IN(GND), 
        .RGMII_TXD2_USBB_DATA5_IN(GND), .RGMII_TXD3_USBB_DATA6_IN(GND), 
        .SPI0_SCK_USBA_XCLK_IN(GND), .SPI0_SDI_USBA_DIR_MGPIO5A_IN(GND)
        , .SPI0_SDO_USBA_STP_MGPIO6A_IN(GND), 
        .SPI0_SS0_USBA_NXT_MGPIO7A_IN(GND), 
        .SPI0_SS1_USBA_DATA5_MGPIO8A_IN(GND), 
        .SPI0_SS2_USBA_DATA6_MGPIO9A_IN(GND), 
        .SPI0_SS3_USBA_DATA7_MGPIO10A_IN(GND), .SPI1_SCK_IN(GND), 
        .SPI1_SDI_MGPIO11A_IN(GND), .SPI1_SDO_MGPIO12A_IN(GND), 
        .SPI1_SS0_MGPIO13A_IN(GND), .SPI1_SS1_MGPIO14A_IN(GND), 
        .SPI1_SS2_MGPIO15A_IN(GND), .SPI1_SS3_MGPIO16A_IN(GND), 
        .SPI1_SS4_MGPIO17A_IN(GND), .SPI1_SS5_MGPIO18A_IN(GND), 
        .SPI1_SS6_MGPIO23A_IN(GND), .SPI1_SS7_MGPIO24A_IN(GND), 
        .USBC_XCLK_IN(GND), .CAN_RXBUS_USBA_DATA1_MGPIO3A_OUT(), 
        .CAN_TX_EBL_USBA_DATA2_MGPIO4A_OUT(), 
        .CAN_TXBUS_USBA_DATA0_MGPIO2A_OUT(), .DRAM_ADDR({nc261, nc262, 
        nc263, nc264, nc265, nc266, nc267, nc268, nc269, nc270, nc271, 
        nc272, nc273, nc274, nc275, nc276}), .DRAM_BA({nc277, nc278, 
        nc279}), .DRAM_CASN(), .DRAM_CKE(), .DRAM_CLK(), .DRAM_CSN(), 
        .DRAM_DM_RDQS_OUT({nc280, nc281, nc282}), .DRAM_DQ_OUT({nc283, 
        nc284, nc285, nc286, nc287, nc288, nc289, nc290, nc291, nc292, 
        nc293, nc294, nc295, nc296, nc297, nc298, nc299, nc300}), 
        .DRAM_DQS_OUT({nc301, nc302, nc303}), .DRAM_FIFO_WE_OUT({nc304, 
        nc305}), .DRAM_ODT(), .DRAM_RASN(), .DRAM_RSTN(), .DRAM_WEN(), 
        .I2C0_SCL_USBC_DATA1_MGPIO31B_OUT(), 
        .I2C0_SDA_USBC_DATA0_MGPIO30B_OUT(), 
        .I2C1_SCL_USBA_DATA4_MGPIO1A_OUT(), 
        .I2C1_SDA_USBA_DATA3_MGPIO0A_OUT(), 
        .MMUART0_CTS_USBC_DATA7_MGPIO19B_OUT(), 
        .MMUART0_DCD_MGPIO22B_OUT(), .MMUART0_DSR_MGPIO20B_OUT(), 
        .MMUART0_DTR_USBC_DATA6_MGPIO18B_OUT(), 
        .MMUART0_RI_MGPIO21B_OUT(), 
        .MMUART0_RTS_USBC_DATA5_MGPIO17B_OUT(), 
        .MMUART0_RXD_USBC_STP_MGPIO28B_OUT(), 
        .MMUART0_SCK_USBC_NXT_MGPIO29B_OUT(), 
        .MMUART0_TXD_USBC_DIR_MGPIO27B_OUT(
        \hello_regs_MSS_0/MSS_ADLIB_INST_MMUART0_TXD_USBC_DIR_MGPIO27B_OUT )
        , .MMUART1_RXD_USBC_DATA3_MGPIO26B_OUT(), 
        .MMUART1_SCK_USBC_DATA4_MGPIO25B_OUT(), 
        .MMUART1_TXD_USBC_DATA2_MGPIO24B_OUT(), 
        .RGMII_GTX_CLK_RMII_CLK_USBB_XCLK_OUT(), 
        .RGMII_MDC_RMII_MDC_OUT(), 
        .RGMII_MDIO_RMII_MDIO_USBB_DATA7_OUT(), .RGMII_RX_CLK_OUT(), 
        .RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_OUT(), 
        .RGMII_RXD0_RMII_RXD0_USBB_DATA0_OUT(), 
        .RGMII_RXD1_RMII_RXD1_USBB_DATA1_OUT(), 
        .RGMII_RXD2_RMII_RX_ER_USBB_DATA3_OUT(), 
        .RGMII_RXD3_USBB_DATA4_OUT(), .RGMII_TX_CLK_OUT(), 
        .RGMII_TX_CTL_RMII_TX_EN_USBB_NXT_OUT(), 
        .RGMII_TXD0_RMII_TXD0_USBB_DIR_OUT(), 
        .RGMII_TXD1_RMII_TXD1_USBB_STP_OUT(), 
        .RGMII_TXD2_USBB_DATA5_OUT(), .RGMII_TXD3_USBB_DATA6_OUT(), 
        .SPI0_SCK_USBA_XCLK_OUT(), .SPI0_SDI_USBA_DIR_MGPIO5A_OUT(), 
        .SPI0_SDO_USBA_STP_MGPIO6A_OUT(), 
        .SPI0_SS0_USBA_NXT_MGPIO7A_OUT(), 
        .SPI0_SS1_USBA_DATA5_MGPIO8A_OUT(), 
        .SPI0_SS2_USBA_DATA6_MGPIO9A_OUT(), 
        .SPI0_SS3_USBA_DATA7_MGPIO10A_OUT(), .SPI1_SCK_OUT(), 
        .SPI1_SDI_MGPIO11A_OUT(), .SPI1_SDO_MGPIO12A_OUT(), 
        .SPI1_SS0_MGPIO13A_OUT(), .SPI1_SS1_MGPIO14A_OUT(), 
        .SPI1_SS2_MGPIO15A_OUT(), .SPI1_SS3_MGPIO16A_OUT(), 
        .SPI1_SS4_MGPIO17A_OUT(), .SPI1_SS5_MGPIO18A_OUT(), 
        .SPI1_SS6_MGPIO23A_OUT(), .SPI1_SS7_MGPIO24A_OUT(), 
        .USBC_XCLK_OUT(), .CAN_RXBUS_USBA_DATA1_MGPIO3A_OE(), 
        .CAN_TX_EBL_USBA_DATA2_MGPIO4A_OE(), 
        .CAN_TXBUS_USBA_DATA0_MGPIO2A_OE(), .DM_OE({nc306, nc307, 
        nc308}), .DRAM_DQ_OE({nc309, nc310, nc311, nc312, nc313, nc314, 
        nc315, nc316, nc317, nc318, nc319, nc320, nc321, nc322, nc323, 
        nc324, nc325, nc326}), .DRAM_DQS_OE({nc327, nc328, nc329}), 
        .I2C0_SCL_USBC_DATA1_MGPIO31B_OE(), 
        .I2C0_SDA_USBC_DATA0_MGPIO30B_OE(), 
        .I2C1_SCL_USBA_DATA4_MGPIO1A_OE(), 
        .I2C1_SDA_USBA_DATA3_MGPIO0A_OE(), 
        .MMUART0_CTS_USBC_DATA7_MGPIO19B_OE(), 
        .MMUART0_DCD_MGPIO22B_OE(), .MMUART0_DSR_MGPIO20B_OE(), 
        .MMUART0_DTR_USBC_DATA6_MGPIO18B_OE(), .MMUART0_RI_MGPIO21B_OE(
        ), .MMUART0_RTS_USBC_DATA5_MGPIO17B_OE(), 
        .MMUART0_RXD_USBC_STP_MGPIO28B_OE(), 
        .MMUART0_SCK_USBC_NXT_MGPIO29B_OE(), 
        .MMUART0_TXD_USBC_DIR_MGPIO27B_OE(
        \hello_regs_MSS_0/MSS_ADLIB_INST_MMUART0_TXD_USBC_DIR_MGPIO27B_OE )
        , .MMUART1_RXD_USBC_DATA3_MGPIO26B_OE(), 
        .MMUART1_SCK_USBC_DATA4_MGPIO25B_OE(), 
        .MMUART1_TXD_USBC_DATA2_MGPIO24B_OE(), 
        .RGMII_GTX_CLK_RMII_CLK_USBB_XCLK_OE(), .RGMII_MDC_RMII_MDC_OE(
        ), .RGMII_MDIO_RMII_MDIO_USBB_DATA7_OE(), .RGMII_RX_CLK_OE(), 
        .RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_OE(), 
        .RGMII_RXD0_RMII_RXD0_USBB_DATA0_OE(), 
        .RGMII_RXD1_RMII_RXD1_USBB_DATA1_OE(), 
        .RGMII_RXD2_RMII_RX_ER_USBB_DATA3_OE(), 
        .RGMII_RXD3_USBB_DATA4_OE(), .RGMII_TX_CLK_OE(), 
        .RGMII_TX_CTL_RMII_TX_EN_USBB_NXT_OE(), 
        .RGMII_TXD0_RMII_TXD0_USBB_DIR_OE(), 
        .RGMII_TXD1_RMII_TXD1_USBB_STP_OE(), .RGMII_TXD2_USBB_DATA5_OE(
        ), .RGMII_TXD3_USBB_DATA6_OE(), .SPI0_SCK_USBA_XCLK_OE(), 
        .SPI0_SDI_USBA_DIR_MGPIO5A_OE(), .SPI0_SDO_USBA_STP_MGPIO6A_OE(
        ), .SPI0_SS0_USBA_NXT_MGPIO7A_OE(), 
        .SPI0_SS1_USBA_DATA5_MGPIO8A_OE(), 
        .SPI0_SS2_USBA_DATA6_MGPIO9A_OE(), 
        .SPI0_SS3_USBA_DATA7_MGPIO10A_OE(), .SPI1_SCK_OE(), 
        .SPI1_SDI_MGPIO11A_OE(), .SPI1_SDO_MGPIO12A_OE(), 
        .SPI1_SS0_MGPIO13A_OE(), .SPI1_SS1_MGPIO14A_OE(), 
        .SPI1_SS2_MGPIO15A_OE(), .SPI1_SS3_MGPIO16A_OE(), 
        .SPI1_SS4_MGPIO17A_OE(), .SPI1_SS5_MGPIO18A_OE(), 
        .SPI1_SS6_MGPIO23A_OE(), .SPI1_SS7_MGPIO24A_OE(), 
        .USBC_XCLK_OE());
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_273  (
        .A(GND), .B(VCC), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_ARLEN_HBURST1_net[1] ), 
        .IPB(\hello_regs_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PSEL_net ), 
        .IPC());
    CFG4 #( .INIT(16'h7350) )  
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_0_2[6]  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_12_[6]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/mem_9_[6]_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/N_644 ), .D(
        \reg_apb_wrp_0/reg16x8_0/N_643 ), .Y(
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_0_2[6]_net_1 ));
    SLE \COREAPBLSRAM_0/PRDATA_reg[7]  (.D(
        \COREAPBLSRAM_0.lsram_width32_PRDATA[7] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB10_rgbr_net_1 ), .EN(
        \COREAPBLSRAM_0.PRDATA4 ), .ALn(
        \hello_regs_MSS_0/MSS_ADLIB_INST_RNIUO3B/U0_RGB1_RGB2_rgbr_net_1 )
        , .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \COREAPBLSRAM_0.PRDATA_reg[7] ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_200_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_77_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_200_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_200_rs_net_1 ));
    CFG2 #( .INIT(4'hD) )  \COREAPBLSRAM_0/g0_1  (.A(
        CoreAPB3_0_APBmslave5_PENABLE), .B(
        CoreAPB3_0_APBmslave5_PWRITE), .Y(N_354));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_2_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB16_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_4__1_sqmuxa ), .ALn(
        AFLSDF_INV_14_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(GND)
        , .Q(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_2_set_net_1 ));
    CFG4 #( .INIT(16'h7350) )  
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_2[5]  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_12_[5]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/mem_9_[5]_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/N_644 ), .D(
        \reg_apb_wrp_0/reg16x8_0/N_643 ), .Y(
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_2[5]_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_1_[3]  (.D(
        \CoreAPB3_0_APBmslave5_PWDATA[3] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB17_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_1__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_155_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_1_rs[3] ));
    INV_BA AFLSDF_INV_106 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_105_net_1 ), .Y(
        AFLSDF_INV_106_net_1));
    INV_BA AFLSDF_INV_52 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_89_net_1 ), .Y(
        AFLSDF_INV_52_net_1));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_249_rs_RNI4ENM  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_59_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_249_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_15_rs[2] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_15_[2]_net_1 ));
    RGB \FCCC_0/GL1_INST/U0_RGB1_RGB2  (.An(\FCCC_0/GL1_INST/U0_YNn ), 
        .ENn(GND), .YL(), .YR(
        \FCCC_0/GL1_INST/U0_RGB1_RGB2_rgbr_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_157_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_42_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_157_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_157_rs_net_1 ));
    SLE \COREAPBLSRAM_0/PRDATA_reg[10]  (.D(
        \COREAPBLSRAM_0.lsram_width32_PRDATA[10] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB8_rgbr_net_1 ), .EN(
        \COREAPBLSRAM_0.PRDATA4 ), .ALn(
        \hello_regs_MSS_0/MSS_ADLIB_INST_RNIUO3B/U0_RGB1_RGB0_rgbr_net_1 )
        , .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \COREAPBLSRAM_0.PRDATA_reg[10] ));
    CFG4 #( .INIT(16'hECA0) )  \CoreAPB3_0/u_mux_p_to_b3/PRDATA_0[28]  
        (.A(\CoreAPB3_0/u_mux_p_to_b3/N_636 ), .B(
        \COREAPBLSRAM_0.PRDATA4 ), .C(\COREAPBLSRAM_0.PRDATA_reg[28] ), 
        .D(\COREAPBLSRAM_0.lsram_width32_PRDATA[28] ), .Y(
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[28] ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_26_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB6_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_5__1_sqmuxa ), .ALn(
        AFLSDF_INV_15_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(GND)
        , .Q(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_26_set_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_10_[6]  (.D(
        \CoreAPB3_0_APBmslave5_PWDATA[6] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB8_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_10__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_178_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_10_rs[6] ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_165_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_35_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_165_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_165_rs_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_154_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_13_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_154_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_154_rs_net_1 ));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_148_rs_RNIC3TN  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_84_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_148_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_0_rs[4] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_0_[4]_net_1 ));
    CFG3 #( .INIT(8'hF2) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_139  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_4_[3]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_648 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_139_i ));
    INV_BA AFLSDF_INV_16 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_83_net_1 ), .Y(
        AFLSDF_INV_16_net_1));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_90_set_RNIMSQD  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_90_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_226_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_11_rs[2] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_11_[2]_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_83_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB17_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_0__1_sqmuxa ), .ALn(
        AFLSDF_INV_16_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(GND)
        , .Q(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_83_set_net_1 ));
    CFG3 #( .INIT(8'hF2) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_251  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_15_[0]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_654 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_251_i ));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_216_rs_RNI1SD6  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_112_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_216_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_14_rs[0] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_14_[0]_net_1 ));
    INV_BA AFLSDF_INV_104 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_76_net_1 ), .Y(
        AFLSDF_INV_104_net_1));
    IOOUTFF_BYPASS \GPIO_OUT_1_obuf[2]/U0/U_IOOUTFF  (.A(
        \GPIO_OUT_1_obuf[2]/U0/DOUT1 ), .Y(
        \GPIO_OUT_1_obuf[2]/U0/DOUT ));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_1_[4]  (.D(
        \CoreAPB3_0_APBmslave5_PWDATA[4] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB15_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_1__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_156_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_1_rs[4] ));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/mem_6__RNIGGAL[5]  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_38_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_173_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_6_rs[5] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_6_[5]_net_1 ));
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_data_out8_61  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_15_[4]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_654 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_61_net_1 ));
    CFG3 #( .INIT(8'hF2) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_223  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_14_[7]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_650 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_223_i ));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_103  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/RCGF_net[3] ), .IPB(
        \hello_regs_MSS_0/MSS_ADLIB_INST/XCLK_FAB_net ), .IPC());
    INV_BA AFLSDF_INV_66 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_63_net_1 ), .Y(
        AFLSDF_INV_66_net_1));
    CFG3 #( .INIT(8'hF2) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_191  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_5_[2]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_653 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_191_i ));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_130  (
        .A(VCC), .B(GND), .C(VCC), .IPA(), .IPB(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[12] ), .IPC(
        ));
    INV_BA AFLSDF_INV_101 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_68_net_1 ), .Y(
        AFLSDF_INV_101_net_1));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_53_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB11_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_3__1_sqmuxa ), .ALn(
        AFLSDF_INV_17_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(GND)
        , .Q(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_53_set_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_101_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB8_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_10__1_sqmuxa ), .ALn(
        AFLSDF_INV_18_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(GND)
        , .Q(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_101_set_net_1 ));
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_data_out8_56  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_15_[3]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_654 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_56_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_32_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB11_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_6__1_sqmuxa ), .ALn(
        AFLSDF_INV_19_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(GND)
        , .Q(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_32_set_net_1 ));
    SLE \COREAPBLSRAM_0/PRDATA_reg[8]  (.D(
        \COREAPBLSRAM_0.lsram_width32_PRDATA[8] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB13_rgbr_net_1 ), .EN(
        \COREAPBLSRAM_0.PRDATA4 ), .ALn(
        \hello_regs_MSS_0/MSS_ADLIB_INST_RNIUO3B/U0_RGB1_RGB5_rgbr_net_1 )
        , .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \COREAPBLSRAM_0.PRDATA_reg[8] ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_149_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_85_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_149_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_149_rs_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_5_[2]  (.D(
        \CoreAPB3_0_APBmslave5_PWDATA[2] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB5_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_5__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_191_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_5_rs[2] ));
    CFG2_IP_BC 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/CFG_17  
        (.B(\CoreAPB3_0_APBmslave5_PWDATA[20] ), .C(
        \CoreAPB3_0_APBmslave5_PADDR[2] ), .IPB(
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/B_DIN_net[4] )
        , .IPC(
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/B_ADDR_net[7] )
        );
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_110_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB9_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_13__1_sqmuxa ), .ALn(
        AFLSDF_INV_20_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(GND)
        , .Q(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_110_set_net_1 ));
    CFG4 #( .INIT(16'h7530) )  
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_3[5]  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_2_[5]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/mem_13_[5]_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/N_646 ), .D(
        \reg_apb_wrp_0/reg16x8_0/N_642 ), .Y(
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_3[5]_net_1 ));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_235  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[33] ), 
        .IPB(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[45] ), 
        .IPC());
    CFG4 #( .INIT(16'hECA0) )  \CoreAPB3_0/u_mux_p_to_b3/PRDATA_0[17]  
        (.A(\CoreAPB3_0/u_mux_p_to_b3/N_636 ), .B(
        \COREAPBLSRAM_0.PRDATA4 ), .C(\COREAPBLSRAM_0.PRDATA_reg[17] ), 
        .D(\COREAPBLSRAM_0.lsram_width32_PRDATA[17] ), .Y(
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[17] ));
    CFG4 #( .INIT(16'h0400) )  
        \reg_apb_wrp_0/reg16x8_0/WRITE_GEN.mem_10__2_i_a2[5]  (.A(
        \CoreAPB3_0_APBmslave5_PADDR[2] ), .B(
        \CoreAPB3_0_APBmslave5_PADDR[5] ), .C(
        \CoreAPB3_0_APBmslave5_PADDR[4] ), .D(
        \CoreAPB3_0_APBmslave5_PADDR[3] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/N_647 ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_193_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_41_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_193_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_193_rs_net_1 ));
    CFG3 #( .INIT(8'hF2) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_203  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_6_[0]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_652 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_203_i ));
    CFG3 #( .INIT(8'hF2) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_152  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_1_[0]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_651 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_152_i ));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_1_[0]  (.D(
        \CoreAPB3_0_APBmslave5_PWDATA[0] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB10_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_1__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_152_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_1_rs[0] ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_180_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_100_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_180_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_180_rs_net_1 ));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_135  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/SMBALERT_NI0_net ), .IPB(
        \hello_regs_MSS_0/MSS_ADLIB_INST/USER_MSS_RESET_N_net ), .IPC()
        );
    INV_BA AFLSDF_INV_44 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_58_net_1 ), .Y(
        AFLSDF_INV_44_net_1));
    CFG4 #( .INIT(16'h4000) )  
        \reg_apb_wrp_0/reg16x8_0/WRITE_GEN.mem_14__2_i_0_0_a2[6]  (.A(
        \CoreAPB3_0_APBmslave5_PADDR[2] ), .B(
        \CoreAPB3_0_APBmslave5_PADDR[5] ), .C(
        \CoreAPB3_0_APBmslave5_PADDR[4] ), .D(
        \CoreAPB3_0_APBmslave5_PADDR[3] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/N_650 ));
    CFG2_IP_BC 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/CFG_27  
        (.B(\CoreAPB3_0_APBmslave5_PWDATA[30] ), .C(
        \CoreAPB3_0_APBmslave5_PADDR[5] ), .IPB(
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/B_DIN_net[15] )
        , .IPC(
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/B_ADDR_net[10] )
        );
    INV_BA AFLSDF_INV_97 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_102_net_1 ), .Y(
        AFLSDF_INV_97_net_1));
    RGB \hello_regs_MSS_0/MSS_ADLIB_INST_RNIUO3B/U0_RGB1_RGB2  (.An(
        \hello_regs_MSS_0/MSS_ADLIB_INST_RNIUO3B/U0_YNn ), .ENn(GND), 
        .YL(), .YR(
        \hello_regs_MSS_0/MSS_ADLIB_INST_RNIUO3B/U0_RGB1_RGB2_rgbr_net_1 )
        );
    INV_BA AFLSDF_INV_51 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_60_net_1 ), .Y(
        AFLSDF_INV_51_net_1));
    INV_BA AFLSDF_INV_38 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_51_net_1 ), .Y(
        AFLSDF_INV_38_net_1));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_217  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[1] ), 
        .IPB(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[13] ), 
        .IPC(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[25] ));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_120  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/FAB_VBUSVALID_net ), .IPB(), 
        .IPC());
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_137  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/I2C1_BCLK_net ), .IPB(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_DMAREADY_net[1] ), .IPC());
    IOOUTFF_BYPASS \GPIO_OUT_1_obuf[5]/U0/U_IOOUTFF  (.A(
        \GPIO_OUT_1_obuf[5]/U0/DOUT1 ), .Y(
        \GPIO_OUT_1_obuf[5]/U0/DOUT ));
    SLE_IP_EN 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/FF_17  
        (.EN(VCC), .IPENn());
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_73  (.A(
        VCC), .B(VCC), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[7] ), 
        .IPB(), .IPC());
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_161  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/SPI1_SDI_F2H_SCP_net ), .IPB(
        \hello_regs_MSS_0/MSS_ADLIB_INST/SPI1_SS1_F2H_SCP_net ), .IPC()
        );
    CFG2 #( .INIT(4'h7) )  
        \CoreAPB3_0/u_mux_p_to_b3/PRDATA_0_iv_0_1_0[6]  (.A(N_637), .B(
        \CoreAPB3_0_APBmslave5_PRDATA[6] ), .Y(
        \CoreAPB3_0/u_mux_p_to_b3/PRDATA_0_iv_0_1_0[6]_net_1 ));
    CFG4 #( .INIT(16'h8C00) )  
        \CoreAPB3_0/u_mux_p_to_b3/PRDATA_0_a2_1[29]  (.A(
        CoreAPB3_0_APBmslave5_PWRITE), .B(
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PADDR[17] ), .C(
        CoreAPB3_0_APBmslave5_PENABLE), .D(N_625), .Y(
        \CoreAPB3_0/u_mux_p_to_b3/N_636 ));
    CFG3 #( .INIT(8'hF2) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_145  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_0_[2]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_645 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_145_i ));
    CFG3 #( .INIT(8'h80) )  
        \reg_apb_wrp_0/reg16x8_0/mem_15__1_sqmuxa_0_a2  (.A(
        \reg_apb_wrp_0/reg16x8_0/N_654 ), .B(N_637), .C(N_638), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_15__1_sqmuxa ));
    CFG3 #( .INIT(8'hF2) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_160  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_2_[0]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_642 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_160_i ));
    sdf_IOPAD_TRI \GPIO_OUT_1_obuf[1]/U0/U_IOPAD  (.PAD(GPIO_OUT_1[1]), 
        .D(\GPIO_OUT_1_obuf[1]/U0/DOUT ), .E(
        \GPIO_OUT_1_obuf[1]/U0/EOUT ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_244_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_20_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_244_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_244_rs_net_1 ));
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_data_out8_78  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_9_[6]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_643 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_78_net_1 ));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/mem_6__RNI4FVN[0]  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_28_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_203_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_6_rs[0] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_6_[0]_net_1 ));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_225  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[9] ), 
        .IPB(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[21] ), 
        .IPC());
    CFG4 #( .INIT(16'h7350) )  
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_5[1]  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_0_[1]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/mem_7_[1]_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/N_645 ), .D(
        \reg_apb_wrp_0/reg16x8_0/N_641 ), .Y(
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_5[1]_net_1 ));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_270  (
        .A(VCC), .B(GND), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[30] ), 
        .IPB(\hello_regs_MSS_0/MSS_ADLIB_INST/F_RREADY_net ), .IPC());
    SLE_IP_EN 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/FF_3  
        (.EN(VCC), .IPENn());
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_94_set_RNITEJG  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_94_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_234_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_11_rs[6] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_11_[6]_net_1 ));
    CFG3 #( .INIT(8'h80) )  
        \CoreAPB3_0/u_mux_p_to_b3/PRDATA_0_iv_0_a2_1[1]  (.A(
        \COREAPBLSRAM_0.PRDATA4_0_a2_0 ), .B(N_625), .C(
        \COREAPBLSRAM_0.lsram_width32_PRDATA[1] ), .Y(
        \CoreAPB3_0/u_mux_p_to_b3/N_585 ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_153_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_11_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_153_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_153_rs_net_1 ));
    INV_BA AFLSDF_INV_135 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_38_net_1 ), .Y(
        AFLSDF_INV_135_net_1));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_44_set_RNICP0N  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_44_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_158_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_1_rs[6] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_1_[6]_net_1 ));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_43  (.A(
        GND), .B(GND), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[26] ), .IPB(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_SEL_net ), .IPC());
    CFG3 #( .INIT(8'hF2) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_175  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_6_[6]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_652 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_175_i ));
    CFG3 #( .INIT(8'hF2) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_143  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_4_[6]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_648 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_143_i ));
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_data_out8_26  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_5_[7]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_653 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_26_net_1 ));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_51  (.A(
        GND), .B(GND), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[5] ), .IPB(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[12] ), .IPC());
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_125  (
        .A(GND), .B(GND), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[0] ), .IPB(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[7] ), .IPC()
        );
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_217_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_113_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_217_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_217_rs_net_1 ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[2].APB_8.GPOUT_reg[2]  (.D(
        \CoreAPB3_0_APBmslave5_PWDATA[2] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB12_rgbr_net_1 ), .EN(
        \CoreGPIO_0/GPOUT_reg35 ), .ALn(
        \hello_regs_MSS_0/MSS_ADLIB_INST_RNIUO3B/U0_RGB1_RGB4_rgbr_net_1 )
        , .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \GPIO_OUT_1_c[2] ));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_19_set_RNIOS9Q  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_19_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_243_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_12_rs[3] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_12_[3]_net_1 ));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/mem_14__RNI42QK[4]  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_116_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_220_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_14_rs[4] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_14_[4]_net_1 ));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_64  (.A(
        GND), .B(VCC), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[25] ), .IPB(
        \hello_regs_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PREADY_net ), 
        .IPC());
    CFG4 #( .INIT(16'h7350) )  
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_0_0[6]  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_11_[6]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/mem_10_[6]_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/N_649 ), .D(
        \reg_apb_wrp_0/reg16x8_0/N_647 ), .Y(
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_0_0[6]_net_1 ));
    CFG3 #( .INIT(8'hF2) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_151  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_0_[7]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_645 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_151_i ));
    INV_BA AFLSDF_INV_99 (.A(AFLSDF_INV_99_net_1), .Y(
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/A_DOUT_EN_net )
        );
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_127  (
        .A(GND), .B(GND), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[2] ), .IPB(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[9] ), .IPC()
        );
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_72  (.A(
        VCC), .B(VCC), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[6] ), 
        .IPB(), .IPC());
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_132  (
        .A(GND), .B(VCC), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[14] ), .IPB(
        ), .IPC());
    CFG4 #( .INIT(16'h7530) )  
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_3[7]  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_2_[7]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/mem_13_[7]_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/N_646 ), .D(
        \reg_apb_wrp_0/reg16x8_0/N_642 ), .Y(
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_3[7]_net_1 ));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/mem_15__RNIR8701[5]  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_62_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_252_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_15_rs[5] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_15_[5]_net_1 ));
    IP_INTERFACE \FCCC_0/CCC_INST/IP_INTERFACE_9  (.A(VCC), .B(GND), 
        .C(VCC), .IPA(\FCCC_0/CCC_INST/PLL_BYPASS_N_net ), .IPB(
        \FCCC_0/CCC_INST/NGMUX3_SEL_net ), .IPC(
        \FCCC_0/CCC_INST/PWDATA_net[7] ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_192_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_73_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_192_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_192_rs_net_1 ));
    CFG2 #( .INIT(4'h8) )  
        \CoreAPB3_0/u_mux_p_to_b3/PRDATA_0_iv_0_a2_2_0[7]  (.A(N_639), 
        .B(\GPIO_OUT_1_c[7] ), .Y(
        \CoreAPB3_0/u_mux_p_to_b3/PRDATA_0_iv_0_a2_2_0[7]_net_1 ));
    INV_BA AFLSDF_INV_102 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_17_net_1 ), .Y(
        AFLSDF_INV_102_net_1));
    CFG2_IP_BC 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/CFG_16  
        (.B(\CoreAPB3_0_APBmslave5_PWDATA[4] ), .C(
        \CoreAPB3_0_APBmslave5_PADDR[2] ), .IPB(
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/A_DIN_net[4] )
        , .IPC(
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/A_ADDR_net[7] )
        );
    CFG3 #( .INIT(8'hF2) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_173  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_6_[5]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_652 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_173_i ));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_68_set_RNIGNVU  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_68_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_142_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_8_rs[4] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_8_[4]_net_1 ));
    CFG3 #( .INIT(8'hF2) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_148  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_0_[4]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_645 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_148_i ));
    CFG4 #( .INIT(16'h7530) )  
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_3[3]  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_2_[3]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/mem_13_[3]_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/N_646 ), .D(
        \reg_apb_wrp_0/reg16x8_0/N_642 ), .Y(
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_3[3]_net_1 ));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_109  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/FAB_XDATAIN_net[1] ), .IPB(), 
        .IPC());
    CFG2_IP_BC 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/CFG_33  
        (.B(GND), .C(\CoreAPB3_0_APBmslave5_PADDR[8] ), .IPB(
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/B_DIN_net[8] )
        , .IPC(
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/B_ADDR_net[13] )
        );
    INV_BA AFLSDF_INV_33 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_70_net_1 ), .Y(
        AFLSDF_INV_33_net_1));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_42  (.A(
        GND), .B(GND), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[25] ), .IPB(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_WRITE_net ), .IPC());
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_10  (.A(
        VCC), .B(\hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[15] ), .C(
        VCC), .IPA(), .IPB(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[15] ), .IPC());
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_22_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB16_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_12__1_sqmuxa ), .ALn(
        AFLSDF_INV_21_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(GND)
        , .Q(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_22_set_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_209_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_105_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_209_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_209_rs_net_1 ));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_236  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[34] ), 
        .IPB(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[46] ), 
        .IPC());
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_108_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB1_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_13__1_sqmuxa ), .ALn(
        AFLSDF_INV_22_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(GND)
        , .Q(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_108_set_net_1 ));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/mem_7__RNIQQ531[1]  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_126_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_181_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_7_rs[1] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_7_[1]_net_1 ));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_274  (
        .A(GND), .B(VCC), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_ARLEN_HBURST1_net[2] ), 
        .IPB(\hello_regs_MSS_0/MSS_ADLIB_INST/CLK_MDDR_APB_net ), .IPC(
        ));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/mem_3__RNIHIVR[0]  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_121_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_128_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_3_rs[0] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_3_[0]_net_1 ));
    SLE_IP_CLK 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/FF_1  
        (.CLK(VCC), .IPCLKn(AFLSDF_INV_23_net_1));
    CFG3 #( .INIT(8'h02) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_115  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_14_[3]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_650 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_115_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_238_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_16_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_238_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_238_rs_net_1 ));
    CFG2_IP_BC 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/CFG_26  
        (.B(\CoreAPB3_0_APBmslave5_PWDATA[14] ), .C(
        \CoreAPB3_0_APBmslave5_PADDR[5] ), .IPB(
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/A_DIN_net[15] )
        , .IPC(
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/A_ADDR_net[10] )
        );
    CFG3 #( .INIT(8'hF2) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_178  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_10_[6]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_647 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_178_i ));
    CFG3 #( .INIT(8'hF2) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_164  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_2_[4]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_642 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_164_i ));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_122  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/FAB_SESSEND_net ), .IPB(), 
        .IPC());
    SLE \reg_apb_wrp_0/reg16x8_0/mem_11_[6]  (.D(
        \CoreAPB3_0_APBmslave5_PWDATA[6] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB6_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_11__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_234_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_11_rs[6] ));
    CFG3 #( .INIT(8'h80) )  \COREAPBLSRAM_0/wen_0_a2  (.A(
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PADDR[17] ), .B(N_638), .C(
        N_625), .Y(\COREAPBLSRAM_0/wen ));
    SLE \COREAPBLSRAM_0/PRDATA_reg[5]  (.D(
        \COREAPBLSRAM_0.lsram_width32_PRDATA[5] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB8_rgbr_net_1 ), .EN(
        \COREAPBLSRAM_0.PRDATA4 ), .ALn(
        \hello_regs_MSS_0/MSS_ADLIB_INST_RNIUO3B/U0_RGB1_RGB0_rgbr_net_1 )
        , .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \COREAPBLSRAM_0.PRDATA_reg[5] ));
    SLE_IP_EN 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/FF_33  
        (.EN(VCC), .IPENn(AFLSDF_INV_24_net_1));
    FLASH_FREEZE \flash_freeze_inst/INST_FLASH_FREEZE_IP  (
        .FF_TO_START(ff_to_start_net), .FF_DONE());
    CFG3 #( .INIT(8'hF2) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_244  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_12_[4]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_644 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_244_i ));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_13_[4]  (.D(
        \CoreAPB3_0_APBmslave5_PWDATA[4] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB1_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_13__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_212_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_13_rs[4] ));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_151  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/CAN_TXBUS_F2H_SCP_net ), .IPB(
        \hello_regs_MSS_0/MSS_ADLIB_INST/MGPIO6A_F2H_GPIN_net ), .IPC()
        );
    INV_BA AFLSDF_INV_70 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_91_net_1 ), .Y(
        AFLSDF_INV_70_net_1));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_152_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_9_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_152_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_152_rs_net_1 ));
    CFG2 #( .INIT(4'h1) )  \reg_apb_wrp_0/reg16x8_0/data_out_RNO[6]  (
        .A(\reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_0_13[6]_net_1 ), 
        .B(\reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_0_12[6]_net_1 ), 
        .Y(\reg_apb_wrp_0/reg16x8_0/N_22_i_0 ));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_5_[5]  (.D(
        \CoreAPB3_0_APBmslave5_PWDATA[5] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB9_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_5__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_197_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_5_rs[5] ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_189_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_14_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_189_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_189_rs_net_1 ));
    INV_BA AFLSDF_INV_108 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_11_net_1 ), .Y(
        AFLSDF_INV_108_net_1));
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_data_out8_63  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_15_[6]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_654 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_63_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_1_[2]  (.D(
        \CoreAPB3_0_APBmslave5_PWDATA[2] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB15_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_1__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_154_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_1_rs[2] ));
    CFG3 #( .INIT(8'h02) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_113  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_14_[1]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_650 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_113_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_15_[3]  (.D(
        \CoreAPB3_0_APBmslave5_PWDATA[3] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB16_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_15__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_250_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_15_rs[3] ));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_12_[4]  (.D(
        \CoreAPB3_0_APBmslave5_PWDATA[4] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB13_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_12__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_244_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_12_rs[4] ));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_68  (.A(
        GND), .B(VCC), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[29] ), .IPB(
        \hello_regs_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[2] ), 
        .IPC());
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_166_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_37_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_166_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_166_rs_net_1 ));
    CFG4 #( .INIT(16'h1000) )  
        \reg_apb_wrp_0/reg16x8_0/WRITE_GEN.mem_6__2_i_0_0_a2[6]  (.A(
        \CoreAPB3_0_APBmslave5_PADDR[2] ), .B(
        \CoreAPB3_0_APBmslave5_PADDR[5] ), .C(
        \CoreAPB3_0_APBmslave5_PADDR[4] ), .D(
        \CoreAPB3_0_APBmslave5_PADDR[3] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/N_652 ));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_104_set_RNI2T9U  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_104_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_208_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_13_rs[0] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_13_[0]_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_119_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB15_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_14__1_sqmuxa ), .ALn(
        AFLSDF_INV_25_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(GND)
        , .Q(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_119_set_net_1 ));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_226  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[10] ), 
        .IPB(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[22] ), 
        .IPC());
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_138  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/SMBALERT_NI1_net ), .IPB(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F2_DMAREADY_net[0] ), .IPC());
    CFG4 #( .INIT(16'h4000) )  \COREAPBLSRAM_0/g0  (.A(
        CoreAPB3_0_APBmslave5_PWRITE), .B(
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PADDR[17] ), .C(
        CoreAPB3_0_APBmslave5_PENABLE), .D(N_625), .Y(
        \COREAPBLSRAM_0.PRDATA4 ));
    CFG4 #( .INIT(16'hFFFE) )  
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_0_13[6]  (.A(
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_0_4[6]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_0_5[6]_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_0_7[6]_net_1 ), .D(
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_0_6[6]_net_1 ), .Y(
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_0_13[6]_net_1 ));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_33  (.A(
        GND), .B(GND), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[9] ), .IPB(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[16] ), .IPC());
    CFG2_IP_BC 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/CFG_3  
        (.B(\CoreAPB3_0_APBmslave5_PWDATA[24] ), .C(GND), .IPB(
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/B_DIN_net[9] )
        , .IPC(
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/B_ADDR_net[1] )
        );
    INV_BA AFLSDF_INV_35 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_87_net_1 ), .Y(
        AFLSDF_INV_35_net_1));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_116  (
        .A(GND), .B(VCC), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/FAB_RXVALIDH_net ), .IPB(
        \hello_regs_MSS_0/MSS_ADLIB_INST/FAB_VSTATUS_net[5] ), .IPC());
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_data_out8_79  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_9_[7]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_643 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_79_net_1 ));
    IOINFF_BYPASS \hello_regs_MSS_0/MMUART_0_RXD_PAD/U_IOINFF  (.A(
        \hello_regs_MSS_0/MMUART_0_RXD_PAD_Y ), .Y(
        \hello_regs_MSS_0/MMUART_0_RXD_PAD/YIN ));
    CFG4 #( .INIT(16'h7350) )  
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_0[7]  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_11_[7]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/mem_10_[7]_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/N_649 ), .D(
        \reg_apb_wrp_0/reg16x8_0/N_647 ), .Y(
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_0[7]_net_1 ));
    IP_INTERFACE \FCCC_0/CCC_INST/IP_INTERFACE_10  (.A(VCC), .B(VCC), 
        .C(VCC), .IPA(\FCCC_0/CCC_INST/PLL_ARST_N_net ), .IPB(
        \FCCC_0/CCC_INST/NGMUX2_HOLD_N_net ), .IPC());
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_data_out8_7  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_8_[0]_net_1 ), .B(N_639), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_7_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_148_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_84_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_148_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_148_rs_net_1 ));
    CFG3 #( .INIT(8'h02) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_118  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_14_[6]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_650 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_118_net_1 ));
    RGB \FCCC_0/GL1_INST/U0_RGB1_RGB7  (.An(\FCCC_0/GL1_INST/U0_YNn ), 
        .ENn(GND), .YL(\FCCC_0/GL1_INST/U0_RGB1_RGB7_rgbl_net_1 ), .YR(
        \FCCC_0/GL1_INST/U0_RGB1_RGB7_rgbr_net_1 ));
    SLE_IP_EN 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/FF_35  
        (.EN(VCC), .IPENn(AFLSDF_INV_26_net_1));
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_data_out8_36  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_6_[4]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_652 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_36_net_1 ));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_194_rs_RNIJ8S31  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_74_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_194_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_9_rs[2] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_9_[2]_net_1 ));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_15_set_RNI42VO  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_15_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_155_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_1_rs[3] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_1_[3]_net_1 ));
    CFG4 #( .INIT(16'hE400) )  
        \CoreAPB3_0/u_mux_p_to_b3/PRDATA_0_iv_0_0[0]  (.A(
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PADDR[17] ), .B(
        \CoreAPB3_0_APBmslave5_PRDATA[0] ), .C(
        \CoreAPB3_0/u_mux_p_to_b3/PRDATA_N_8_0 ), .D(N_625), .Y(
        \CoreAPB3_0/u_mux_p_to_b3/PRDATA_0_iv_0_0[0]_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_14_[4]  (.D(
        \CoreAPB3_0_APBmslave5_PWDATA[4] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB11_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_14__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_220_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_14_rs[4] ));
    IOENFF_BYPASS \GPIO_OUT_1_obuf[2]/U0/U_IOENFF  (.A(
        \GPIO_OUT_1_obuf[2]/U0/EOUT1 ), .Y(
        \GPIO_OUT_1_obuf[2]/U0/EOUT ));
    SLE \reg_apb_wrp_0/reg16x8_0/data_out[7]  (.D(
        \reg_apb_wrp_0/reg16x8_0/N_84_i_0 ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB10_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/rd_enable ), .ALn(
        \hello_regs_MSS_0/MSS_ADLIB_INST_RNIUO3B/U0_RGB1_RGB2_rgbr_net_1 )
        , .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreAPB3_0_APBmslave5_PRDATA[7] ));
    CFG4 #( .INIT(16'hFFFE) )  
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_12[0]  (.A(
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_1[0]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_3[0]_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_2[0]_net_1 ), .D(
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_0[0]_net_1 ), .Y(
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_12[0]_net_1 ));
    SLE_IP_EN 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/FF_13  
        (.EN(VCC), .IPENn());
    SLE \reg_apb_wrp_0/reg16x8_0/mem_5_[7]  (.D(
        \CoreAPB3_0_APBmslave5_PWDATA[7] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB6_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_5__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_201_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_5_rs[7] ));
    SLE \COREAPBLSRAM_0/PRDATA_reg[31]  (.D(
        \COREAPBLSRAM_0.lsram_width32_PRDATA[31] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB10_rgbr_net_1 ), .EN(
        \COREAPBLSRAM_0.PRDATA4 ), .ALn(
        \hello_regs_MSS_0/MSS_ADLIB_INST_RNIUO3B/U0_RGB1_RGB2_rgbr_net_1 )
        , .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \COREAPBLSRAM_0.PRDATA_reg[31] ));
    INV_BA AFLSDF_INV_94 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_14_net_1 ), .Y(
        AFLSDF_INV_94_net_1));
    CFG3 #( .INIT(8'h80) )  
        \reg_apb_wrp_0/reg16x8_0/mem_2__1_sqmuxa_0_a2  (.A(
        \reg_apb_wrp_0/reg16x8_0/N_642 ), .B(N_637), .C(N_638), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_2__1_sqmuxa ));
    CFG4 #( .INIT(16'hECA0) )  \CoreAPB3_0/u_mux_p_to_b3/PRDATA_0[21]  
        (.A(\CoreAPB3_0/u_mux_p_to_b3/N_636 ), .B(
        \COREAPBLSRAM_0.PRDATA4 ), .C(\COREAPBLSRAM_0.PRDATA_reg[21] ), 
        .D(\COREAPBLSRAM_0.lsram_width32_PRDATA[21] ), .Y(
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[21] ));
    SLE_IP_EN 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/FF_30  
        (.EN(VCC), .IPENn(AFLSDF_INV_27_net_1));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_128  (
        .A(GND), .B(GND), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[3] ), .IPB(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[10] ), .IPC(
        ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_84_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB14_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_0__1_sqmuxa ), .ALn(
        AFLSDF_INV_28_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(GND)
        , .Q(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_84_set_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_177_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_122_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_177_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_177_rs_net_1 ));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_32  (.A(
        GND), .B(GND), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[8] ), .IPB(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[15] ), .IPC());
    INV_BA AFLSDF_INV_10 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_115_net_1 ), .Y(
        AFLSDF_INV_10_net_1));
    CFG4 #( .INIT(16'h0040) )  
        \reg_apb_wrp_0/reg16x8_0/WRITE_GEN.mem_12__2_i_a2[0]  (.A(
        \CoreAPB3_0_APBmslave5_PADDR[2] ), .B(
        \CoreAPB3_0_APBmslave5_PADDR[5] ), .C(
        \CoreAPB3_0_APBmslave5_PADDR[4] ), .D(
        \CoreAPB3_0_APBmslave5_PADDR[3] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/N_644 ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_161_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_27_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_161_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_161_rs_net_1 ));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_5  (.A(
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[3] ), .B(
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[10] ), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[3] ), .IPB(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[10] ), .IPC());
    CFG3 #( .INIT(8'hF2) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_214  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_13_[6]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_646 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_214_i ));
    SLE_IP_EN 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/FF_21  
        (.EN(VCC), .IPENn());
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_174_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_101_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_174_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_174_rs_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_221_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_117_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_221_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_221_rs_net_1 ));
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_data_out8_48  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_7_[2]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_641 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_48_net_1 ));
    CFG3 #( .INIT(8'hF2) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_169  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_6_[3]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_652 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_169_i ));
    INV_BA AFLSDF_INV_60 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_1_net_1 ), .Y(
        AFLSDF_INV_60_net_1));
    INV_BA AFLSDF_INV_125 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_45_net_1 ), .Y(
        AFLSDF_INV_125_net_1));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_54_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB15_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_7__1_sqmuxa ), .ALn(
        AFLSDF_INV_29_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(GND)
        , .Q(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_54_set_net_1 ));
    CFG4 #( .INIT(16'h4F00) )  
        \CoreAPB3_0/u_mux_p_to_b3/PRDATA_0_iv_0_1[4]  (.A(
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PADDR[17] ), .B(
        \CoreAPB3_0_APBmslave5_PRDATA[4] ), .C(
        \CoreAPB3_0/u_mux_p_to_b3/PRDATA_m3_i_0_net_1 ), .D(N_625), .Y(
        \CoreAPB3_0/u_mux_p_to_b3/PRDATA_0_iv_0_1[4]_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_202_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_78_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_202_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_202_rs_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_0_[1]  (.D(
        \CoreAPB3_0_APBmslave5_PWDATA[1] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB18_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_0__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_144_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_0_rs[1] ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_90_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB5_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_11__1_sqmuxa ), .ALn(
        AFLSDF_INV_30_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(GND)
        , .Q(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_90_set_net_1 ));
    CFG3 #( .INIT(8'h02) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_126  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_7_[1]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_641 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_126_net_1 ));
    CFG4 #( .INIT(16'h7530) )  
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_7[4]  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_8_[4]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/mem_5_[4]_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/N_653 ), .D(N_639), .Y(
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_7[4]_net_1 ));
    CFG4 #( .INIT(16'hECA0) )  \CoreAPB3_0/u_mux_p_to_b3/PRDATA_0[9]  
        (.A(\CoreAPB3_0/u_mux_p_to_b3/N_636 ), .B(
        \COREAPBLSRAM_0.PRDATA4 ), .C(\COREAPBLSRAM_0.PRDATA_reg[9] ), 
        .D(\COREAPBLSRAM_0.lsram_width32_PRDATA[9] ), .Y(
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[9] ));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_2_[3]  (.D(
        \CoreAPB3_0_APBmslave5_PWDATA[3] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB5_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_2__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_163_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_2_rs[3] ));
    RGB \FCCC_0/GL1_INST/U0_RGB1_RGB15  (.An(
        \FCCC_0/GL1_INST/U0_YNn_GSouth ), .ENn(GND), .YL(
        \FCCC_0/GL1_INST/U0_RGB1_RGB15_rgbl_net_1 ), .YR(
        \FCCC_0/GL1_INST/U0_RGB1_RGB15_rgbr_net_1 ));
    SLE_IP_EN 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/FF_15  
        (.EN(VCC), .IPENn());
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_209  (
        .A(VCC), .B(GND), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[27] ), 
        .IPB(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_AWBURST_HTRANS0_net[1] ), 
        .IPC());
    CFG4 #( .INIT(16'h7350) )  
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_5[5]  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_0_[5]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/mem_7_[5]_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/N_645 ), .D(
        \reg_apb_wrp_0/reg16x8_0/N_641 ), .Y(
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_5[5]_net_1 ));
    CFG4 #( .INIT(16'h7350) )  
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_2[3]  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_12_[3]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/mem_9_[3]_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/N_644 ), .D(
        \reg_apb_wrp_0/reg16x8_0/N_643 ), .Y(
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_2[3]_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_195_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_47_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_195_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_195_rs_net_1 ));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_267  (
        .A(VCC), .B(GND), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[27] ), 
        .IPB(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_ARLOCK_HMASTLOCK1_net[1] ), 
        .IPC());
    RGB \FCCC_0/GL1_INST/U0_RGB1_RGB0  (.An(\FCCC_0/GL1_INST/U0_YNn ), 
        .ENn(GND), .YL(), .YR(
        \FCCC_0/GL1_INST/U0_RGB1_RGB0_rgbr_net_1 ));
    IOTRI_OB_EB \GPIO_OUT_1_obuf[6]/U0/U_IOTRI  (.D(\GPIO_OUT_1_c[6] ), 
        .E(VCC), .DOUT(\GPIO_OUT_1_obuf[6]/U0/DOUT1 ), .EOUT(
        \GPIO_OUT_1_obuf[6]/U0/EOUT1 ));
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_data_out8_75  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_9_[3]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_643 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_75_net_1 ));
    INV_BA AFLSDF_INV_46 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_123_net_1 ), .Y(
        AFLSDF_INV_46_net_1));
    SLE_IP_EN 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/FF_10  
        (.EN(VCC), .IPENn(AFLSDF_INV_31_net_1));
    CFG4 #( .INIT(16'h8F0F) )  
        \CoreAPB3_0/u_mux_p_to_b3/PRDATA_0_iv_0[3]  (.A(N_639), .B(
        \GPIO_OUT_1_c[3] ), .C(
        \CoreAPB3_0/u_mux_p_to_b3/PRDATA_0_iv_0_1[3]_net_1 ), .D(
        \CoreAPB3_0.u_mux_p_to_b3.PRDATA_0_iv_0_a2_3_5[1] ), .Y(
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[3] ));
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_data_out8_82  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_0_[2]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_645 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_82_net_1 ));
    CFG3 #( .INIT(8'h02) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_106  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_13_[2]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_646 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_106_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_106_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB2_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_13__1_sqmuxa ), .ALn(
        AFLSDF_INV_32_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(GND)
        , .Q(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_106_set_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_2_[4]  (.D(
        \CoreAPB3_0_APBmslave5_PWDATA[4] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB0_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_2__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_164_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_2_rs[4] ));
    INV_BA AFLSDF_INV_32 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_106_net_1 ), .Y(
        AFLSDF_INV_32_net_1));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_208  (
        .A(VCC), .B(GND), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[26] ), 
        .IPB(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_AWBURST_HTRANS0_net[0] ), 
        .IPC());
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/mem_7__RNIMSVP[7]  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_1_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_233_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_7_rs[7] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_7_[7]_net_1 ));
    INV_BA AFLSDF_INV_5 (.A(AFLSDF_INV_5_net_1), .Y(
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/B_BLK_net[1] )
        );
    CFG2_IP_BC 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/CFG_32  
        (.B(GND), .C(\CoreAPB3_0_APBmslave5_PADDR[8] ), .IPB(
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/A_DIN_net[8] )
        , .IPC(
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/A_ADDR_net[13] )
        );
    SLE \reg_apb_wrp_0/reg16x8_0/mem_3_[1]  (.D(
        \CoreAPB3_0_APBmslave5_PWDATA[1] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB15_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_3__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_129_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_3_rs[1] ));
    CFG3 #( .INIT(8'hF2) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_135  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_3_[7]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_655 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_135_i ));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_1_[5]  (.D(
        \CoreAPB3_0_APBmslave5_PWDATA[5] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB10_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_1__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_157_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_1_rs[5] ));
    CFG2_IP_BC 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/CFG_18  
        (.B(\CoreAPB3_0_APBmslave5_PWDATA[12] ), .C(
        \CoreAPB3_0_APBmslave5_PADDR[3] ), .IPB(
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/A_DIN_net[13] )
        , .IPC(
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/A_ADDR_net[8] )
        );
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_110_set_RNI2GL71  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_110_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_214_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_13_rs[6] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_13_[6]_net_1 ));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_56  (.A(
        GND), .B(GND), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[10] ), .IPB(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[17] ), .IPC());
    CFG4 #( .INIT(16'hECA0) )  \CoreAPB3_0/u_mux_p_to_b3/PRDATA_0[13]  
        (.A(\CoreAPB3_0/u_mux_p_to_b3/N_636 ), .B(
        \COREAPBLSRAM_0.PRDATA4 ), .C(\COREAPBLSRAM_0.PRDATA_reg[13] ), 
        .D(\COREAPBLSRAM_0.lsram_width32_PRDATA[13] ), .Y(
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[13] ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_251_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_57_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_251_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_251_rs_net_1 ));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_113  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/FAB_XDATAIN_net[5] ), .IPB(
        \hello_regs_MSS_0/MSS_ADLIB_INST/FAB_VSTATUS_net[2] ), .IPC());
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_155_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_15_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_155_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_155_rs_net_1 ));
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_data_out8_80  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_0_[0]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_645 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_80_net_1 ));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_63_set_RNIUGGL  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_63_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_253_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_15_rs[6] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_15_[6]_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_7_[1]  (.D(
        \CoreAPB3_0_APBmslave5_PWDATA[1] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB16_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_7__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_181_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_7_rs[1] ));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_79_set_RNIL2ET  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_79_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_204_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_9_rs[7] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_9_[7]_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_173_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_38_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_173_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_173_rs_net_1 ));
    INV_BA AFLSDF_INV_115 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_72_net_1 ), .Y(
        AFLSDF_INV_115_net_1));
    CFG3 #( .INIT(8'hF2) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_133  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_3_[5]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_655 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_133_i ));
    sdf_IOPAD_TRI \hello_regs_MSS_0/MMUART_0_TXD_PAD/U_IOPAD  (.PAD(
        MMUART_0_TXD), .D(
        \hello_regs_MSS_0/MSS_ADLIB_INST_MMUART0_TXD_USBC_DIR_MGPIO27B_OUT )
        , .E(
        \hello_regs_MSS_0/MSS_ADLIB_INST_MMUART0_TXD_USBC_DIR_MGPIO27B_OE )
        );
    CFG4 #( .INIT(16'h7530) )  
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_0_4[6]  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_6_[6]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/mem_3_[6]_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/N_655 ), .D(
        \reg_apb_wrp_0/reg16x8_0/N_652 ), .Y(
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_0_4[6]_net_1 ));
    CFG2_IP_BC 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/CFG_28  
        (.B(\CoreAPB3_0_APBmslave5_PWDATA[7] ), .C(
        \CoreAPB3_0_APBmslave5_PADDR[6] ), .IPB(
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/A_DIN_net[7] )
        , .IPC(
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/A_ADDR_net[11] )
        );
    SLE \reg_apb_wrp_0/reg16x8_0/mem_2_[0]  (.D(
        \CoreAPB3_0_APBmslave5_PWDATA[0] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB5_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_2__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_160_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_2_rs[0] ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_237_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_5_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_237_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_237_rs_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_188_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_71_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_188_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_188_rs_net_1 ));
    CFG3 #( .INIT(8'h80) )  
        \reg_apb_wrp_0/reg16x8_0/mem_10__1_sqmuxa_0_a2  (.A(
        \reg_apb_wrp_0/reg16x8_0/N_647 ), .B(N_637), .C(N_638), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_10__1_sqmuxa ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_70_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB7_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_8__1_sqmuxa ), .ALn(
        AFLSDF_INV_33_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(GND)
        , .Q(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_70_set_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_8_[1]  (.D(
        \CoreAPB3_0_APBmslave5_PWDATA[1] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB5_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_8__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_237_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_8_rs[1] ));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/mem_3__RNI8EOO[6]  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_53_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_134_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_3_rs[6] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_3_[6]_net_1 ));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/mem_12__RNII1001[4]  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_20_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_244_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_12_rs[4] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_12_[4]_net_1 ));
    INV_BA AFLSDF_INV_100 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_33_net_1 ), .Y(
        AFLSDF_INV_100_net_1));
    CFG3 #( .INIT(8'hF2) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_252  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_15_[5]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_654 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_252_i ));
    CFG4 #( .INIT(16'h0008) )  
        \reg_apb_wrp_0/reg16x8_0/WRITE_GEN.mem_9__2_i_0_0_a2[6]  (.A(
        \CoreAPB3_0_APBmslave5_PADDR[2] ), .B(
        \CoreAPB3_0_APBmslave5_PADDR[5] ), .C(
        \CoreAPB3_0_APBmslave5_PADDR[4] ), .D(
        \CoreAPB3_0_APBmslave5_PADDR[3] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/N_643 ));
    CFG4 #( .INIT(16'h2000) )  
        \reg_apb_wrp_0/reg16x8_0/WRITE_GEN.mem_7__2_i_a2[1]  (.A(
        \CoreAPB3_0_APBmslave5_PADDR[2] ), .B(
        \CoreAPB3_0_APBmslave5_PADDR[5] ), .C(
        \CoreAPB3_0_APBmslave5_PADDR[4] ), .D(
        \CoreAPB3_0_APBmslave5_PADDR[3] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/N_641 ));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_97_set_RNIOAJE  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_97_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_206_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_10_rs[0] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_10_[0]_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_1_[7]  (.D(
        \CoreAPB3_0_APBmslave5_PWDATA[7] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB16_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_1__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_159_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_1_rs[7] ));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_202  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[6] ), 
        .IPB(\hello_regs_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[18] )
        , .IPC());
    CFG3 #( .INIT(8'hF2) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_221  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_14_[5]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_650 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_221_i ));
    CFG3 #( .INIT(8'hF2) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_138  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_4_[2]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_648 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_138_i ));
    IOOUTFF_BYPASS \GPIO_OUT_1_obuf[3]/U0/U_IOOUTFF  (.A(
        \GPIO_OUT_1_obuf[3]/U0/DOUT1 ), .Y(
        \GPIO_OUT_1_obuf[3]/U0/DOUT ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_104_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB4_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_13__1_sqmuxa ), .ALn(
        AFLSDF_INV_34_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(GND)
        , .Q(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_104_set_net_1 ));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_203  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[7] ), 
        .IPB(\hello_regs_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[19] )
        , .IPC());
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_230_rs_RNILOQJ  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_92_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_230_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_11_rs[4] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_11_[4]_net_1 ));
    RGB \FCCC_0/GL1_INST/U0_RGB1_RGB17  (.An(
        \FCCC_0/GL1_INST/U0_YNn_GSouth ), .ENn(GND), .YL(
        \FCCC_0/GL1_INST/U0_RGB1_RGB17_rgbl_net_1 ), .YR(
        \FCCC_0/GL1_INST/U0_RGB1_RGB17_rgbr_net_1 ));
    CCC #( .INIT(210'h0000007FB8000044D64000318C6318C1F18C61EC0404040400301)
        , .VCOFREQUENCY(800.0) )  \FCCC_0/CCC_INST/INST_CCC_IP  (.Y0(), 
        .Y1(), .Y2(), .Y3(), .PRDATA({nc330, nc331, nc332, nc333, 
        nc334, nc335, nc336, nc337}), .LOCK(FCCC_0_LOCK), .BUSY(), 
        .CLK0(\FCCC_0/CCC_INST/CLK0_net ), .CLK1(
        \FCCC_0/CCC_INST/CLK1_net ), .CLK2(\FCCC_0/CCC_INST/CLK2_net ), 
        .CLK3(\FCCC_0/CCC_INST/CLK3_net ), .NGMUX0_SEL(
        \FCCC_0/CCC_INST/NGMUX0_SEL_net ), .NGMUX1_SEL(
        \FCCC_0/CCC_INST/NGMUX1_SEL_net ), .NGMUX2_SEL(
        \FCCC_0/CCC_INST/NGMUX2_SEL_net ), .NGMUX3_SEL(
        \FCCC_0/CCC_INST/NGMUX3_SEL_net ), .NGMUX0_HOLD_N(
        \FCCC_0/CCC_INST/NGMUX0_HOLD_N_net ), .NGMUX1_HOLD_N(
        \FCCC_0/CCC_INST/NGMUX1_HOLD_N_net ), .NGMUX2_HOLD_N(
        \FCCC_0/CCC_INST/NGMUX2_HOLD_N_net ), .NGMUX3_HOLD_N(
        \FCCC_0/CCC_INST/NGMUX3_HOLD_N_net ), .NGMUX0_ARST_N(
        \FCCC_0/CCC_INST/NGMUX0_ARST_N_net ), .NGMUX1_ARST_N(
        \FCCC_0/CCC_INST/NGMUX1_ARST_N_net ), .NGMUX2_ARST_N(
        \FCCC_0/CCC_INST/NGMUX2_ARST_N_net ), .NGMUX3_ARST_N(
        \FCCC_0/CCC_INST/NGMUX3_ARST_N_net ), .PLL_BYPASS_N(
        \FCCC_0/CCC_INST/PLL_BYPASS_N_net ), .PLL_ARST_N(
        \FCCC_0/CCC_INST/PLL_ARST_N_net ), .PLL_POWERDOWN_N(
        \FCCC_0/CCC_INST/PLL_POWERDOWN_N_net ), .GPD0_ARST_N(
        \FCCC_0/CCC_INST/GPD0_ARST_N_net ), .GPD1_ARST_N(
        \FCCC_0/CCC_INST/GPD1_ARST_N_net ), .GPD2_ARST_N(
        \FCCC_0/CCC_INST/GPD2_ARST_N_net ), .GPD3_ARST_N(
        \FCCC_0/CCC_INST/GPD3_ARST_N_net ), .PRESET_N(
        \FCCC_0/CCC_INST/PRESET_N_net ), .PCLK(
        \FCCC_0/CCC_INST/PCLK_net ), .PSEL(\FCCC_0/CCC_INST/PSEL_net ), 
        .PENABLE(\FCCC_0/CCC_INST/PENABLE_net ), .PWRITE(
        \FCCC_0/CCC_INST/PWRITE_net ), .PADDR({
        \FCCC_0/CCC_INST/PADDR_net[7] , \FCCC_0/CCC_INST/PADDR_net[6] , 
        \FCCC_0/CCC_INST/PADDR_net[5] , \FCCC_0/CCC_INST/PADDR_net[4] , 
        \FCCC_0/CCC_INST/PADDR_net[3] , \FCCC_0/CCC_INST/PADDR_net[2] })
        , .PWDATA({\FCCC_0/CCC_INST/PWDATA_net[7] , 
        \FCCC_0/CCC_INST/PWDATA_net[6] , 
        \FCCC_0/CCC_INST/PWDATA_net[5] , 
        \FCCC_0/CCC_INST/PWDATA_net[4] , 
        \FCCC_0/CCC_INST/PWDATA_net[3] , 
        \FCCC_0/CCC_INST/PWDATA_net[2] , 
        \FCCC_0/CCC_INST/PWDATA_net[1] , 
        \FCCC_0/CCC_INST/PWDATA_net[0] }), .CLK0_PAD(GND), .CLK1_PAD(
        GND), .CLK2_PAD(GND), .CLK3_PAD(GND), .GL0(\FCCC_0/GL1_net ), 
        .GL1(), .GL2(), .GL3(), .RCOSC_25_50MHZ(
        OSC_0_RCOSC_25_50MHZ_CCC_OUT_RCOSC_25_50MHZ_CCC), .RCOSC_1MHZ(
        GND), .XTLOSC(GND));
    CFG2_IP_BC 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/CFG_4  
        (.B(\CoreAPB3_0_APBmslave5_PWDATA[1] ), .C(GND), .IPB(
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/A_DIN_net[1] )
        , .IPC(
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/A_ADDR_net[2] )
        );
    INV_BA AFLSDF_INV_133 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_8_net_1 ), .Y(
        AFLSDF_INV_133_net_1));
    CFG4 #( .INIT(16'hECA0) )  \CoreAPB3_0/u_mux_p_to_b3/PRDATA_0[25]  
        (.A(\CoreAPB3_0/u_mux_p_to_b3/N_636 ), .B(
        \COREAPBLSRAM_0.PRDATA4 ), .C(\COREAPBLSRAM_0.PRDATA_reg[25] ), 
        .D(\COREAPBLSRAM_0.lsram_width32_PRDATA[25] ), .Y(
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[25] ));
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_data_out8_49  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_3_[4]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_655 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_49_net_1 ));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_257  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[5] ), 
        .IPB(\hello_regs_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[17] )
        , .IPC());
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_data_out8_4  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_4_[2]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_648 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_4_net_1 ));
    INV_BA AFLSDF_INV_31 (.A(AFLSDF_INV_31_net_1), .Y(
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/A_BLK_net[1] )
        );
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_87_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB15_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_0__1_sqmuxa ), .ALn(
        AFLSDF_INV_35_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(GND)
        , .Q(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_87_set_net_1 ));
    CFG3 #( .INIT(8'hF2) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_147  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_0_[0]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_645 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_147_i ));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_4_[1]  (.D(
        \CoreAPB3_0_APBmslave5_PWDATA[1] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB17_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_4__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_137_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_4_rs[1] ));
    CFG4 #( .INIT(16'h7530) )  
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_4[4]  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_6_[4]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/mem_3_[4]_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/N_655 ), .D(
        \reg_apb_wrp_0/reg16x8_0/N_652 ), .Y(
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_4[4]_net_1 ));
    IOTRI_OB_EB \GPIO_OUT_1_obuf[3]/U0/U_IOTRI  (.D(\GPIO_OUT_1_c[3] ), 
        .E(VCC), .DOUT(\GPIO_OUT_1_obuf[3]/U0/DOUT1 ), .EOUT(
        \GPIO_OUT_1_obuf[3]/U0/EOUT1 ));
    CFG4 #( .INIT(16'h7530) )  
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_7[5]  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_8_[5]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/mem_5_[5]_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/N_653 ), .D(N_639), .Y(
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_7[5]_net_1 ));
    CFG2_IP_BC 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/CFG_19  
        (.B(\CoreAPB3_0_APBmslave5_PWDATA[28] ), .C(
        \CoreAPB3_0_APBmslave5_PADDR[3] ), .IPB(
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/B_DIN_net[13] )
        , .IPC(
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/B_ADDR_net[8] )
        );
    SLE \COREAPBLSRAM_0/PRDATA_reg[21]  (.D(
        \COREAPBLSRAM_0.lsram_width32_PRDATA[21] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB9_rgbr_net_1 ), .EN(
        \COREAPBLSRAM_0.PRDATA4 ), .ALn(
        \hello_regs_MSS_0/MSS_ADLIB_INST_RNIUO3B/U0_RGB1_RGB1_rgbr_net_1 )
        , .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \COREAPBLSRAM_0.PRDATA_reg[21] ));
    CFG4 #( .INIT(16'hECA0) )  \CoreAPB3_0/u_mux_p_to_b3/PRDATA_0[16]  
        (.A(\CoreAPB3_0/u_mux_p_to_b3/N_636 ), .B(
        \COREAPBLSRAM_0.PRDATA4 ), .C(\COREAPBLSRAM_0.PRDATA_reg[16] ), 
        .D(\COREAPBLSRAM_0.lsram_width32_PRDATA[16] ), .Y(
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[16] ));
    SLE \COREAPBLSRAM_0/PRDATA_reg[1]  (.D(
        \COREAPBLSRAM_0.lsram_width32_PRDATA[1] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB9_rgbr_net_1 ), .EN(
        \COREAPBLSRAM_0.PRDATA4 ), .ALn(
        \hello_regs_MSS_0/MSS_ADLIB_INST_RNIUO3B/U0_RGB1_RGB1_rgbr_net_1 )
        , .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \COREAPBLSRAM_0.PRDATA_reg[1] ));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_6_[1]  (.D(
        \CoreAPB3_0_APBmslave5_PWDATA[1] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB10_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_6__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_205_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_6_rs[1] ));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_13_[5]  (.D(
        \CoreAPB3_0_APBmslave5_PWDATA[5] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB2_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_13__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_213_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_13_rs[5] ));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_271  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[31] ), 
        .IPB(\hello_regs_MSS_0/MSS_ADLIB_INST/FPGA_MDDR_ARESET_N_net ), 
        .IPC());
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_99  (.A(
        VCC), .B(VCC), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/GTX_CLKPF_net ), .IPB(
        \hello_regs_MSS_0/MSS_ADLIB_INST/RCGF_net[6] ), .IPC());
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_141  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F2HCALIB_net ), .IPB(
        \hello_regs_MSS_0/MSS_ADLIB_INST/SPI0_CLK_IN_net ), .IPC());
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_16_set_RNIMO0V  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_16_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_238_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_12_rs[0] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_12_[0]_net_1 ));
    CFG3 #( .INIT(8'h80) )  
        \reg_apb_wrp_0/reg16x8_0/mem_12__1_sqmuxa_0_a2  (.A(
        \reg_apb_wrp_0/reg16x8_0/N_644 ), .B(N_637), .C(N_638), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_12__1_sqmuxa ));
    CFG3 #( .INIT(8'hF2) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_201  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_5_[7]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_653 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_201_i ));
    CFG3 #( .INIT(8'hF2) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_234  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_11_[6]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_649 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_234_i ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_57_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB16_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_15__1_sqmuxa ), .ALn(
        AFLSDF_INV_36_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(GND)
        , .Q(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_57_set_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_15_[7]  (.D(
        \CoreAPB3_0_APBmslave5_PWDATA[7] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB15_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_15__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_254_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_15_rs[7] ));
    CFG3 #( .INIT(8'hF2) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_177  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_6_[7]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_652 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_177_i ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_240_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_17_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_240_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_240_rs_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_206_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_97_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_206_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_206_rs_net_1 ));
    SLE \COREAPBLSRAM_0/PRDATA_reg[25]  (.D(
        \COREAPBLSRAM_0.lsram_width32_PRDATA[25] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB10_rgbr_net_1 ), .EN(
        \COREAPBLSRAM_0.PRDATA4 ), .ALn(
        \hello_regs_MSS_0/MSS_ADLIB_INST_RNIUO3B/U0_RGB1_RGB2_rgbr_net_1 )
        , .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \COREAPBLSRAM_0.PRDATA_reg[25] ));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_12_[5]  (.D(
        \CoreAPB3_0_APBmslave5_PWDATA[5] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB13_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_12__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_245_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_12_rs[5] ));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_186_rs_RNIJQTS  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_70_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_186_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_8_rs[6] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_8_[6]_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_172_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_96_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_172_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_172_rs_net_1 ));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_55  (.A(
        GND), .B(GND), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[9] ), .IPB(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[16] ), .IPC());
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_166  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(), .IPB(
        \hello_regs_MSS_0/MSS_ADLIB_INST/MGPIO11B_F2H_GPIN_net ), .IPC(
        ));
    IP_INTERFACE \FCCC_0/CCC_INST/IP_INTERFACE_7  (.A(VCC), .B(VCC), 
        .C(VCC), .IPA(\FCCC_0/CCC_INST/CLK3_net ), .IPB(), .IPC(
        \FCCC_0/CCC_INST/PWDATA_net[5] ));
    CFG3 #( .INIT(8'h02) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_122  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_6_[7]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_652 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_122_net_1 ));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_97  (.A(
        VCC), .B(VCC), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/COLF_net ), .IPB(), .IPC());
    CFG2_IP_BC 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/CFG_29  
        (.B(\CoreAPB3_0_APBmslave5_PWDATA[23] ), .C(
        \CoreAPB3_0_APBmslave5_PADDR[6] ), .IPB(
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/B_DIN_net[7] )
        , .IPC(
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/B_ADDR_net[11] )
        );
    CFG3 #( .INIT(8'h80) )  
        \reg_apb_wrp_0/reg16x8_0/mem_11__1_sqmuxa_0_a2  (.A(
        \reg_apb_wrp_0/reg16x8_0/N_649 ), .B(N_637), .C(N_638), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_11__1_sqmuxa ));
    SLE \COREAPBLSRAM_0/PRDATA_reg[24]  (.D(
        \COREAPBLSRAM_0.lsram_width32_PRDATA[24] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB10_rgbr_net_1 ), .EN(
        \COREAPBLSRAM_0.PRDATA4 ), .ALn(
        \hello_regs_MSS_0/MSS_ADLIB_INST_RNIUO3B/U0_RGB1_RGB2_rgbr_net_1 )
        , .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \COREAPBLSRAM_0.PRDATA_reg[24] ));
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_data_out8_66  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_8_[3]_net_1 ), .B(N_639), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_66_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_81_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB18_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_0__1_sqmuxa ), .ALn(
        AFLSDF_INV_37_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(GND)
        , .Q(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_81_set_net_1 ));
    CFG3 #( .INIT(8'h80) )  
        \reg_apb_wrp_0/reg16x8_0/mem_9__1_sqmuxa_0_a2_0_a2  (.A(
        \reg_apb_wrp_0/reg16x8_0/N_643 ), .B(N_637), .C(N_638), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_9__1_sqmuxa ));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_127_set_RNIKSKH  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_127_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_131_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_3_rs[3] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_3_[3]_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_205_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_30_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_205_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_205_rs_net_1 ));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/mem_2__RNIVS5M[0]  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_25_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_160_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_2_rs[0] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_2_[0]_net_1 ));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_119  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(), .IPB(
        \hello_regs_MSS_0/MSS_ADLIB_INST/FAB_RXERROR_net ), .IPC());
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_63  (.A(
        GND), .B(GND), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[24] ), .IPB(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[31] ), .IPC());
    SLE \reg_apb_wrp_0/reg16x8_0/mem_14_[5]  (.D(
        \CoreAPB3_0_APBmslave5_PWDATA[5] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB11_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_14__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_221_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_14_rs[5] ));
    CFG4 #( .INIT(16'h7350) )  
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_0_5[6]  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_0_[6]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/mem_7_[6]_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/N_645 ), .D(
        \reg_apb_wrp_0/reg16x8_0/N_641 ), .Y(
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_0_5[6]_net_1 ));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_29  (.A(
        GND), .B(GND), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[5] ), .IPB(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[12] ), .IPC());
    CFG3 #( .INIT(8'h02) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_102  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_10_[5]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_647 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_102_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/data_out[4]  (.D(
        \reg_apb_wrp_0/reg16x8_0/N_41_i_0 ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB10_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/rd_enable ), .ALn(
        \hello_regs_MSS_0/MSS_ADLIB_INST_RNIUO3B/U0_RGB1_RGB2_rgbr_net_1 )
        , .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreAPB3_0_APBmslave5_PRDATA[4] ));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_11  (.A(
        VCC), .B(\hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[16] ), .C(
        VCC), .IPA(), .IPB(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[16] ), .IPC());
    IOTRI_OB_EB \GPIO_OUT_1_obuf[4]/U0/U_IOTRI  (.D(\GPIO_OUT_1_c[4] ), 
        .E(VCC), .DOUT(\GPIO_OUT_1_obuf[4]/U0/DOUT1 ), .EOUT(
        \GPIO_OUT_1_obuf[4]/U0/EOUT1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_51_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB13_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_3__1_sqmuxa ), .ALn(
        AFLSDF_INV_38_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(GND)
        , .Q(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_51_set_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_13_[0]  (.D(
        \CoreAPB3_0_APBmslave5_PWDATA[0] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB2_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_13__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_208_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_13_rs[0] ));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_194  (
        .A(GND), .B(VCC), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_AWID_HSEL0_net[2] ), .IPB(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[10] ), 
        .IPC());
    IOENFF_BYPASS \GPIO_OUT_1_obuf[3]/U0/U_IOENFF  (.A(
        \GPIO_OUT_1_obuf[3]/U0/EOUT1 ), .Y(
        \GPIO_OUT_1_obuf[3]/U0/EOUT ));
    SLE_IP_EN 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/FF_28  
        (.EN(VCC), .IPENn());
    CFG1_IP_B 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/CFG_11  
        (.B(\CoreAPB3_0_APBmslave5_PWDATA[26] ), .IPB(
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/B_DIN_net[11] )
        );
    INV_BA AFLSDF_INV_96 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_61_net_1 ), .Y(
        AFLSDF_INV_96_net_1));
    CFG3 #( .INIT(8'h02) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_117  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_14_[5]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_650 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_117_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_196_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_75_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_196_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_196_rs_net_1 ));
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_data_out8_45  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_5_[5]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_653 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_45_net_1 ));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_192_rs_RNIFTFT  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_73_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_192_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_9_rs[1] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_9_[1]_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_15_[2]  (.D(
        \CoreAPB3_0_APBmslave5_PWDATA[2] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB17_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_15__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_249_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_15_rs[2] ));
    INV_BA AFLSDF_INV_57 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_94_net_1 ), .Y(
        AFLSDF_INV_57_net_1));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_27  (.A(
        GND), .B(GND), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[3] ), .IPB(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[10] ), .IPC());
    CFG4 #( .INIT(16'h7350) )  
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_1[1]  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_15_[1]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/mem_14_[1]_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/N_654 ), .D(
        \reg_apb_wrp_0/reg16x8_0/N_650 ), .Y(
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_1[1]_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_2_[2]  (.D(
        \CoreAPB3_0_APBmslave5_PWDATA[2] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB5_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_2__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_162_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_2_rs[2] ));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_12_[0]  (.D(
        \CoreAPB3_0_APBmslave5_PWDATA[0] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB18_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_12__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_238_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_12_rs[0] ));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/mem_6__RNI0RUI[1]  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_30_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_205_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_6_rs[1] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_6_[1]_net_1 ));
    CFG4 #( .INIT(16'h7350) )  
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_0[3]  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_11_[3]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/mem_10_[3]_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/N_649 ), .D(
        \reg_apb_wrp_0/reg16x8_0/N_647 ), .Y(
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_0[3]_net_1 ));
    SLE_IP_EN 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/FF_4  
        (.EN(VCC), .IPENn());
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_181  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/MMUART0_DCD_F2H_SCP_net ), 
        .IPB(), .IPC());
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/mem_6__RNI5AHT[2]  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_32_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_207_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_6_rs[2] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_6_[2]_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_223_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_119_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_223_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_223_rs_net_1 ));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_200_rs_RNIDCL01  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_77_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_200_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_9_rs[5] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_9_[5]_net_1 ));
    CFG3 #( .INIT(8'h02) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_121  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_3_[0]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_655 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_121_net_1 ));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_174  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/MGPIO25B_F2H_GPIN_net ), .IPB(
        \hello_regs_MSS_0/MSS_ADLIB_INST/MMUART0_DTR_F2H_SCP_net ), 
        .IPC());
    IOENFF_BYPASS \MSS_RESET_N_M2F_obuf/U0/U_IOENFF  (.A(
        \MSS_RESET_N_M2F_obuf/U0/EOUT1 ), .Y(
        \MSS_RESET_N_M2F_obuf/U0/EOUT ));
    CFG4 #( .INIT(16'hECA0) )  \CoreAPB3_0/u_mux_p_to_b3/PRDATA_0[14]  
        (.A(\CoreAPB3_0/u_mux_p_to_b3/N_636 ), .B(
        \COREAPBLSRAM_0.PRDATA4 ), .C(\COREAPBLSRAM_0.PRDATA_reg[14] ), 
        .D(\COREAPBLSRAM_0.lsram_width32_PRDATA[14] ), .Y(
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[14] ));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_10_[3]  (.D(
        \CoreAPB3_0_APBmslave5_PWDATA[3] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB11_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_10__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_172_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_10_rs[3] ));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_62  (.A(
        GND), .B(VCC), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[23] ), .IPB(), 
        .IPC());
    CFG2_IP_BC 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/CFG_21  
        (.B(\CoreAPB3_0_APBmslave5_PWDATA[21] ), .C(
        \COREAPBLSRAM_0/wen ), .IPB(
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/B_DIN_net[5] )
        , .IPC(
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/A_WEN_net[1] )
        );
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_data_out8_58  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_15_[1]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_654 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_58_net_1 ));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_200  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[4] ), 
        .IPB(\hello_regs_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[16] )
        , .IPC());
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_93_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB5_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_11__1_sqmuxa ), .ALn(
        AFLSDF_INV_39_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(GND)
        , .Q(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_93_set_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_214_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_110_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_214_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_214_rs_net_1 ));
    CFG4 #( .INIT(16'h7350) )  
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_2[7]  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_12_[7]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/mem_9_[7]_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/N_644 ), .D(
        \reg_apb_wrp_0/reg16x8_0/N_643 ), .Y(
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_2[7]_net_1 ));
    CFG0 #( .INIT(1'h0) )  CFG0_GND_INST (.Y(CFG0_GND_INST_NET));
    CFG4 #( .INIT(16'hECA0) )  \CoreAPB3_0/u_mux_p_to_b3/PRDATA_0[27]  
        (.A(\CoreAPB3_0/u_mux_p_to_b3/N_636 ), .B(
        \COREAPBLSRAM_0.PRDATA4 ), .C(\COREAPBLSRAM_0.PRDATA_reg[27] ), 
        .D(\COREAPBLSRAM_0.lsram_width32_PRDATA[27] ), .Y(
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[27] ));
    CFG4 #( .INIT(16'hEAC0) )  
        \CoreAPB3_0/u_mux_p_to_b3/PRDATA_0_iv_0_0[5]  (.A(
        \COREAPBLSRAM_0.PRDATA_reg[5] ), .B(
        \CoreAPB3_0/u_mux_p_to_b3/PRDATA_0_iv_0_a2_2_0[5]_net_1 ), .C(
        \CoreAPB3_0.u_mux_p_to_b3.PRDATA_0_iv_0_a2_3_5[1] ), .D(
        \CoreAPB3_0/u_mux_p_to_b3/N_636 ), .Y(
        \CoreAPB3_0/u_mux_p_to_b3/PRDATA_0_iv_0_0[5]_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_14_[0]  (.D(
        \CoreAPB3_0_APBmslave5_PWDATA[0] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB15_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_14__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_216_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_14_rs[0] ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_156_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_40_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_156_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_156_rs_net_1 ));
    SLE \COREAPBLSRAM_0/PRDATA_reg[2]  (.D(
        \COREAPBLSRAM_0.lsram_width32_PRDATA[2] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB8_rgbr_net_1 ), .EN(
        \COREAPBLSRAM_0.PRDATA4 ), .ALn(
        \hello_regs_MSS_0/MSS_ADLIB_INST_RNIUO3B/U0_RGB1_RGB0_rgbr_net_1 )
        , .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \COREAPBLSRAM_0.PRDATA_reg[2] ));
    CFG3 #( .INIT(8'h02) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_101  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_10_[4]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_647 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_101_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_9_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB11_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_1__1_sqmuxa ), .ALn(
        AFLSDF_INV_40_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(GND)
        , .Q(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_9_set_net_1 ));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_156  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/MGPIO9A_F2H_GPIN_net ), .IPB()
        , .IPC());
    SLE \reg_apb_wrp_0/reg16x8_0/mem_9_[1]  (.D(
        \CoreAPB3_0_APBmslave5_PWDATA[1] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB19_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_9__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_192_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_9_rs[1] ));
    INV_BA AFLSDF_INV_59 (.A(AFLSDF_INV_59_net_1), .Y(
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/B_ARST_N_net )
        );
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_88_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB6_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_11__1_sqmuxa ), .ALn(
        AFLSDF_INV_41_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(GND)
        , .Q(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_88_set_net_1 ));
    SLE_IP_EN 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/FF_31  
        (.EN(VCC), .IPENn(AFLSDF_INV_42_net_1));
    CFG2 #( .INIT(4'h8) )  
        \CoreAPB3_0/u_mux_p_to_b3/PRDATA_0_iv_0_a2_2_0[5]  (.A(N_639), 
        .B(\GPIO_OUT_1_c[5] ), .Y(
        \CoreAPB3_0/u_mux_p_to_b3/PRDATA_0_iv_0_a2_2_0[5]_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_191_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_43_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_191_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_191_rs_net_1 ));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_89  (.A(
        VCC), .B(VCC), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[30] ), 
        .IPB(\hello_regs_MSS_0/MSS_ADLIB_INST/RXDF_net[5] ), .IPC());
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_data_out8_94  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_11_[6]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_649 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_94_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_6_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB16_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_4__1_sqmuxa ), .ALn(
        AFLSDF_INV_43_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(GND)
        , .Q(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_6_set_net_1 ));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/mem_11__RNISSFV[0]  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_88_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_182_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_11_rs[0] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_11_[0]_net_1 ));
    INV_BA AFLSDF_INV_40 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_9_net_1 ), .Y(
        AFLSDF_INV_40_net_1));
    INV_BA AFLSDF_INV_123 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_24_net_1 ), .Y(
        AFLSDF_INV_123_net_1));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_163  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/SPI1_SDO_F2H_SCP_net ), .IPB(
        \hello_regs_MSS_0/MSS_ADLIB_INST/SPI1_SS2_F2H_SCP_net ), .IPC()
        );
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_58_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB12_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_15__1_sqmuxa ), .ALn(
        AFLSDF_INV_44_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(GND)
        , .Q(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_58_set_net_1 ));
    CFG3 #( .INIT(8'hF2) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_180  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_10_[7]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_647 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_180_i ));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_87  (.A(
        VCC), .B(VCC), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[28] ), 
        .IPB(\hello_regs_MSS_0/MSS_ADLIB_INST/RXDF_net[3] ), .IPC());
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_253_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_63_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_253_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_253_rs_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_4_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB18_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_4__1_sqmuxa ), .ALn(
        AFLSDF_INV_45_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(GND)
        , .Q(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_4_set_net_1 ));
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_data_out8_97  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_10_[0]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_647 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_97_net_1 ));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_204  (
        .A(VCC), .B(GND), .C(GND), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[22] ), 
        .IPB(\hello_regs_MSS_0/MSS_ADLIB_INST/F_AWLEN_HBURST0_net[0] ), 
        .IPC(\hello_regs_MSS_0/MSS_ADLIB_INST/F_AWVALID_HWRITE0_net ));
    INV_BA AFLSDF_INV_88 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_43_net_1 ), .Y(
        AFLSDF_INV_88_net_1));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_123_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB16_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_3__1_sqmuxa ), .ALn(
        AFLSDF_INV_46_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(GND)
        , .Q(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_123_set_net_1 ));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/mem_10__RNI2KPJ[4]  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_101_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_174_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_10_rs[4] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_10_[4]_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_85_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB13_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_0__1_sqmuxa ), .ALn(
        AFLSDF_INV_47_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(GND)
        , .Q(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_85_set_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_151_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_87_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_151_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_151_rs_net_1 ));
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_data_out8_28  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_6_[0]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_652 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_28_net_1 ));
    CFG3 #( .INIT(8'hF2) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_165  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_2_[5]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_642 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_165_i ));
    RAM1K18 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/INST_RAM1K18_IP  
        (.A_DOUT({nc338, \COREAPBLSRAM_0.lsram_width32_PRDATA[15] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[14] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[13] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[12] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[11] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[10] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[9] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[8] , nc339, 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[7] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[6] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[5] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[4] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[3] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[2] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[1] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[0] }), .B_DOUT({nc340, 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[31] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[30] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[29] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[28] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[27] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[26] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[25] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[24] , nc341, 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[23] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[22] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[21] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[20] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[19] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[18] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[17] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[16] }), .BUSY(), .A_CLK(
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/A_CLK_net )
        , .A_DOUT_CLK(
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/A_DOUT_CLK_net )
        , .A_ARST_N(
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/A_ARST_N_net )
        , .A_DOUT_EN(
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/A_DOUT_EN_net )
        , .A_BLK({
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/A_BLK_net[2] , 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/A_BLK_net[1] , 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/A_BLK_net[0] })
        , .A_DOUT_ARST_N(
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/A_DOUT_ARST_N_net )
        , .A_DOUT_SRST_N(
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/A_DOUT_SRST_N_net )
        , .A_DIN({
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/A_DIN_net[17] , 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/A_DIN_net[16] , 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/A_DIN_net[15] , 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/A_DIN_net[14] , 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/A_DIN_net[13] , 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/A_DIN_net[12] , 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/A_DIN_net[11] , 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/A_DIN_net[10] , 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/A_DIN_net[9] , 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/A_DIN_net[8] , 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/A_DIN_net[7] , 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/A_DIN_net[6] , 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/A_DIN_net[5] , 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/A_DIN_net[4] , 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/A_DIN_net[3] , 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/A_DIN_net[2] , 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/A_DIN_net[1] , 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/A_DIN_net[0] })
        , .A_ADDR({
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/A_ADDR_net[13] , 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/A_ADDR_net[12] , 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/A_ADDR_net[11] , 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/A_ADDR_net[10] , 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/A_ADDR_net[9] , 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/A_ADDR_net[8] , 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/A_ADDR_net[7] , 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/A_ADDR_net[6] , 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/A_ADDR_net[5] , 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/A_ADDR_net[4] , 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/A_ADDR_net[3] , 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/A_ADDR_net[2] , 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/A_ADDR_net[1] , 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/A_ADDR_net[0] })
        , .A_WEN({
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/A_WEN_net[1] , 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/A_WEN_net[0] })
        , .B_CLK(
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/B_CLK_net )
        , .B_DOUT_CLK(
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/B_DOUT_CLK_net )
        , .B_ARST_N(
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/B_ARST_N_net )
        , .B_DOUT_EN(
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/B_DOUT_EN_net )
        , .B_BLK({
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/B_BLK_net[2] , 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/B_BLK_net[1] , 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/B_BLK_net[0] })
        , .B_DOUT_ARST_N(
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/B_DOUT_ARST_N_net )
        , .B_DOUT_SRST_N(
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/B_DOUT_SRST_N_net )
        , .B_DIN({
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/B_DIN_net[17] , 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/B_DIN_net[16] , 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/B_DIN_net[15] , 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/B_DIN_net[14] , 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/B_DIN_net[13] , 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/B_DIN_net[12] , 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/B_DIN_net[11] , 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/B_DIN_net[10] , 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/B_DIN_net[9] , 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/B_DIN_net[8] , 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/B_DIN_net[7] , 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/B_DIN_net[6] , 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/B_DIN_net[5] , 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/B_DIN_net[4] , 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/B_DIN_net[3] , 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/B_DIN_net[2] , 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/B_DIN_net[1] , 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/B_DIN_net[0] })
        , .B_ADDR({
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/B_ADDR_net[13] , 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/B_ADDR_net[12] , 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/B_ADDR_net[11] , 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/B_ADDR_net[10] , 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/B_ADDR_net[9] , 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/B_ADDR_net[8] , 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/B_ADDR_net[7] , 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/B_ADDR_net[6] , 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/B_ADDR_net[5] , 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/B_ADDR_net[4] , 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/B_ADDR_net[3] , 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/B_ADDR_net[2] , 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/B_ADDR_net[1] , 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/B_ADDR_net[0] })
        , .B_WEN({
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/B_WEN_net[1] , 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/B_WEN_net[0] })
        , .A_EN(VCC), .A_DOUT_LAT(VCC), .A_WIDTH({VCC, GND, VCC}), 
        .A_WMODE(GND), .B_EN(VCC), .B_DOUT_LAT(VCC), .B_WIDTH({VCC, 
        GND, VCC}), .B_WMODE(GND), .SII_LOCK(GND));
    CFG4 #( .INIT(16'h35FF) )  
        \CoreAPB3_0/u_mux_p_to_b3/PRDATA_m3_i_0  (.A(
        \COREAPBLSRAM_0.lsram_width32_PRDATA[4] ), .B(
        \COREAPBLSRAM_0.PRDATA_reg[4] ), .C(N_354), .D(
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PADDR[17] ), .Y(
        \CoreAPB3_0/u_mux_p_to_b3/PRDATA_m3_i_0_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_175_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_120_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_175_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_175_rs_net_1 ));
    CFG3 #( .INIT(8'h80) )  
        \reg_apb_wrp_0/reg16x8_0/mem_13__1_sqmuxa_0_a2  (.A(
        \reg_apb_wrp_0/reg16x8_0/N_646 ), .B(N_637), .C(N_638), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_13__1_sqmuxa ));
    IOENFF_BYPASS \GPIO_OUT_1_obuf[5]/U0/U_IOENFF  (.A(
        \GPIO_OUT_1_obuf[5]/U0/EOUT1 ), .Y(
        \GPIO_OUT_1_obuf[5]/U0/EOUT ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_130_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_125_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_130_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_130_rs_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_73_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB19_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_9__1_sqmuxa ), .ALn(
        AFLSDF_INV_48_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(GND)
        , .Q(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_73_set_net_1 ));
    INV_BA AFLSDF_INV_137 (.A(AFLSDF_INV_137_net_1), .Y(
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/A_BLK_net[0] )
        );
    SLE_IP_EN 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/FF_11  
        (.EN(VCC), .IPENn(AFLSDF_INV_49_net_1));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_219  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[3] ), 
        .IPB(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[15] ), 
        .IPC());
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_data_out8_14  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_5_[1]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_653 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_14_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_55_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB13_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_3__1_sqmuxa ), .ALn(
        AFLSDF_INV_50_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(GND)
        , .Q(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_55_set_net_1 ));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_24_set_RNIJI051  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_24_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_199_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_5_rs[6] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_5_[6]_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_249_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_59_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_249_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_249_rs_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_15_[1]  (.D(
        \CoreAPB3_0_APBmslave5_PWDATA[1] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB13_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_15__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_248_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_15_rs[1] ));
    CFG3 #( .INIT(8'hF2) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_163  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_2_[3]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_642 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_163_i ));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_1  (.A(
        GND), .B(VCC), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_HM0_RESP_net ), .IPB(), 
        .IPC());
    RGB \FCCC_0/GL1_INST/U0_RGB1_RGB6  (.An(\FCCC_0/GL1_INST/U0_YNn ), 
        .ENn(GND), .YL(\FCCC_0/GL1_INST/U0_RGB1_RGB6_rgbl_net_1 ), .YR(
        \FCCC_0/GL1_INST/U0_RGB1_RGB6_rgbr_net_1 ));
    CFG4 #( .INIT(16'hFFFE) )  
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_13[7]  (.A(
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_4[7]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_5[7]_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_7[7]_net_1 ), .D(
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_6[7]_net_1 ), .Y(
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_13[7]_net_1 ));
    SLE \COREAPBLSRAM_0/PRDATA_reg[11]  (.D(
        \COREAPBLSRAM_0.lsram_width32_PRDATA[11] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB8_rgbr_net_1 ), .EN(
        \COREAPBLSRAM_0.PRDATA4 ), .ALn(
        \hello_regs_MSS_0/MSS_ADLIB_INST_RNIUO3B/U0_RGB1_RGB0_rgbr_net_1 )
        , .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \COREAPBLSRAM_0.PRDATA_reg[11] ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_60_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB15_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_15__1_sqmuxa ), .ALn(
        AFLSDF_INV_51_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(GND)
        , .Q(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_60_set_net_1 ));
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_data_out8_91  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_11_[3]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_649 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_91_net_1 ));
    sdf_IOPAD_TRI \MSS_RESET_N_M2F_obuf/U0/U_IOPAD  (.PAD(
        MSS_RESET_N_M2F), .D(\MSS_RESET_N_M2F_obuf/U0/DOUT ), .E(
        \MSS_RESET_N_M2F_obuf/U0/EOUT ));
    CFG4 #( .INIT(16'h0002) )  
        \reg_apb_wrp_0/reg16x8_0/WRITE_GEN.mem_1__2_i_a2[3]  (.A(
        \CoreAPB3_0_APBmslave5_PADDR[2] ), .B(
        \CoreAPB3_0_APBmslave5_PADDR[5] ), .C(
        \CoreAPB3_0_APBmslave5_PADDR[4] ), .D(
        \CoreAPB3_0_APBmslave5_PADDR[3] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/N_651 ));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_191_rs_RNI8SLS  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_43_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_191_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_5_rs[2] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_5_[2]_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_2_[5]  (.D(
        \CoreAPB3_0_APBmslave5_PWDATA[5] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB2_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_2__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_165_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_2_rs[5] ));
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_data_out8_59  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_15_[2]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_654 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_59_net_1 ));
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_data_out8_17  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_12_[1]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_644 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_17_net_1 ));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_247  (
        .A(VCC), .B(GND), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[59] ), 
        .IPB(\hello_regs_MSS_0/MSS_ADLIB_INST/F_WSTRB_net[7] ), .IPC());
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_89_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB6_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_11__1_sqmuxa ), .ALn(
        AFLSDF_INV_52_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(GND)
        , .Q(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_89_set_net_1 ));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_218  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[2] ), 
        .IPB(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[14] ), 
        .IPC());
    SLE \COREAPBLSRAM_0/PRDATA_reg[28]  (.D(
        \COREAPBLSRAM_0.lsram_width32_PRDATA[28] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB13_rgbr_net_1 ), .EN(
        \COREAPBLSRAM_0.PRDATA4 ), .ALn(
        \hello_regs_MSS_0/MSS_ADLIB_INST_RNIUO3B/U0_RGB1_RGB5_rgbr_net_1 )
        , .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \COREAPBLSRAM_0.PRDATA_reg[28] ));
    INV_BA AFLSDF_INV_113 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_100_net_1 ), .Y(
        AFLSDF_INV_113_net_1));
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_data_out8_5  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_8_[1]_net_1 ), .B(N_639), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_5_net_1 ));
    SLE \COREAPBLSRAM_0/PRDATA_reg[22]  (.D(
        \COREAPBLSRAM_0.lsram_width32_PRDATA[22] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB14_rgbr_net_1 ), .EN(
        \COREAPBLSRAM_0.PRDATA4 ), .ALn(
        \hello_regs_MSS_0/MSS_ADLIB_INST_RNIUO3B/U0_RGB1_RGB6_rgbr_net_1 )
        , .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \COREAPBLSRAM_0.PRDATA_reg[22] ));
    CFG3 #( .INIT(8'hF2) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_184  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_8_[5]_net_1 ), .B(N_639), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_184_i ));
    CFG3 #( .INIT(8'hF2) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_137  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_4_[1]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_648 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_137_i ));
    SLE \COREAPBLSRAM_0/PRDATA_reg[15]  (.D(
        \COREAPBLSRAM_0.lsram_width32_PRDATA[15] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB9_rgbr_net_1 ), .EN(
        \COREAPBLSRAM_0.PRDATA4 ), .ALn(
        \hello_regs_MSS_0/MSS_ADLIB_INST_RNIUO3B/U0_RGB1_RGB1_rgbr_net_1 )
        , .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \COREAPBLSRAM_0.PRDATA_reg[15] ));
    CFG2 #( .INIT(4'h7) )  
        \CoreAPB3_0/u_mux_p_to_b3/PRDATA_0_iv_0_1_0[5]  (.A(N_637), .B(
        \CoreAPB3_0_APBmslave5_PRDATA[5] ), .Y(
        \CoreAPB3_0/u_mux_p_to_b3/PRDATA_0_iv_0_1_0[5]_net_1 ));
    CFG3 #( .INIT(8'hF2) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_168  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_10_[1]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_647 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_168_i ));
    INV_BA AFLSDF_INV_3 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_29_net_1 ), .Y(
        AFLSDF_INV_3_net_1));
    CFG4 #( .INIT(16'h7530) )  
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_7[7]  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_8_[7]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/mem_5_[7]_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/N_653 ), .D(N_639), .Y(
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_7[7]_net_1 ));
    INV_BA AFLSDF_INV_54 (.A(AFLSDF_INV_54_net_1), .Y(
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/A_CLK_net )
        );
    INV_BA AFLSDF_INV_83 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_64_net_1 ), .Y(
        AFLSDF_INV_83_net_1));
    SLE \COREAPBLSRAM_0/PRDATA_reg[14]  (.D(
        \COREAPBLSRAM_0.lsram_width32_PRDATA[14] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB9_rgbr_net_1 ), .EN(
        \COREAPBLSRAM_0.PRDATA4 ), .ALn(
        \hello_regs_MSS_0/MSS_ADLIB_INST_RNIUO3B/U0_RGB1_RGB1_rgbr_net_1 )
        , .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \COREAPBLSRAM_0.PRDATA_reg[14] ));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_153  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/CAN_RXBUS_F2H_SCP_net ), .IPB(
        \hello_regs_MSS_0/MSS_ADLIB_INST/MGPIO7A_F2H_GPIN_net ), .IPC()
        );
    INV_BA AFLSDF_INV_109 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_92_net_1 ), .Y(
        AFLSDF_INV_109_net_1));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_59_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB17_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_15__1_sqmuxa ), .ALn(
        AFLSDF_INV_53_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(GND)
        , .Q(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_59_set_net_1 ));
    SLE_IP_CLK 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/FF_0  
        (.CLK(\FCCC_0/GL1_INST/U0_RGB1_RGB0_rgbr_net_1 ), .IPCLKn(
        AFLSDF_INV_54_net_1));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_11_[3]  (.D(
        \CoreAPB3_0_APBmslave5_PWDATA[3] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB7_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_11__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_228_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_11_rs[3] ));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_54  (.A(
        GND), .B(GND), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[8] ), .IPB(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[15] ), .IPC());
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_113_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB13_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_14__1_sqmuxa ), .ALn(
        AFLSDF_INV_55_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(GND)
        , .Q(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_113_set_net_1 ));
    RCOSC_25_50MHZ #( .FREQUENCY(50.0) )  \OSC_0/I_RCOSC_25_50MHZ  (
        .CLKOUT(OSC_0_RCOSC_25_50MHZ_CCC_OUT_RCOSC_25_50MHZ_CCC));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_170  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/MMUART1_RI_F2H_SCP_net ), 
        .IPB(), .IPC());
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_data_out8_72  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_9_[0]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_643 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_72_net_1 ));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_169  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/MMUART1_DSR_F2H_SCP_net ), 
        .IPB(), .IPC());
    CFG3 #( .INIT(8'hF2) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_190  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_9_[0]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_643 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_190_i ));
    CFG2_IP_BC 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/CFG_9  
        (.B(\CoreAPB3_0_APBmslave5_PWDATA[18] ), .C(GND), .IPB(
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/B_DIN_net[2] )
        , .IPC(
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/B_ADDR_net[4] )
        );
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_data_out8_11  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_1_[1]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_651 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_11_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_2_[7]  (.D(
        \CoreAPB3_0_APBmslave5_PWDATA[7] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB3_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_2__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_167_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_2_rs[7] ));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_13_[6]  (.D(
        \CoreAPB3_0_APBmslave5_PWDATA[6] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB9_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_13__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_214_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_13_rs[6] ));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/mem_2__RNIAMVL[5]  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_35_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_165_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_2_rs[5] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_2_[5]_net_1 ));
    CFG4 #( .INIT(16'hFFFE) )  
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_12[7]  (.A(
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_1[7]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_3[7]_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_2[7]_net_1 ), .D(
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_0[7]_net_1 ), .Y(
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_12[7]_net_1 ));
    sdf_IOPAD_TRI \GPIO_OUT_1_obuf[5]/U0/U_IOPAD  (.PAD(GPIO_OUT_1[5]), 
        .D(\GPIO_OUT_1_obuf[5]/U0/DOUT ), .E(
        \GPIO_OUT_1_obuf[5]/U0/EOUT ));
    CFG4 #( .INIT(16'h7530) )  
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_4[0]  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_6_[0]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/mem_3_[0]_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/N_655 ), .D(
        \reg_apb_wrp_0/reg16x8_0/N_652 ), .Y(
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_4[0]_net_1 ));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_275  (
        .A(GND), .B(GND), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_ARLEN_HBURST1_net[3] ), 
        .IPB(\hello_regs_MSS_0/MSS_ADLIB_INST/PRESET_N_net ), .IPC());
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_195  (
        .A(GND), .B(VCC), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_AWID_HSEL0_net[3] ), .IPB(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[11] ), 
        .IPC());
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_16  (.A(
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[21] ), .B(
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[28] ), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[21] ), .IPB(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[28] ), .IPC());
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_data_out8_38  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_6_[5]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_652 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_38_net_1 ));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_64_set_RNIHR0S  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_64_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_239_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_8_rs[2] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_8_[2]_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_12_[6]  (.D(
        \CoreAPB3_0_APBmslave5_PWDATA[6] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB16_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_12__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_246_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_12_rs[6] ));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_212  (
        .A(VCC), .B(GND), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[30] ), 
        .IPB(\hello_regs_MSS_0/MSS_ADLIB_INST/F_WID_HREADY01_net[0] ), 
        .IPC());
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_197  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[1] ), 
        .IPB(\hello_regs_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[13] )
        , .IPC());
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_79  (.A(
        VCC), .B(VCC), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[13] ), 
        .IPB(
        \hello_regs_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[20] ), 
        .IPC());
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_213  (
        .A(VCC), .B(GND), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[31] ), 
        .IPB(\hello_regs_MSS_0/MSS_ADLIB_INST/F_WID_HREADY01_net[1] ), 
        .IPC());
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_287  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PADDR_net[10] ), 
        .IPB(
        \hello_regs_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[14] ), 
        .IPC());
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_data_out8_29  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_2_[2]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_642 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_29_net_1 ));
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_data_out8_70  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_8_[6]_net_1 ), .B(N_639), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_70_net_1 ));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_175  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/MMUART1_SCK_F2H_SCP_net ), 
        .IPB(\hello_regs_MSS_0/MSS_ADLIB_INST/MGPIO19B_F2H_GPIN_net ), 
        .IPC());
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_139_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_6_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_139_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_139_rs_net_1 ));
    INV_BA AFLSDF_INV_85 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_78_net_1 ), .Y(
        AFLSDF_INV_85_net_1));
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_data_out8_2  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_4_[1]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_648 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_2_net_1 ));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/mem_2__RNIIEUO[7]  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_39_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_167_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_2_rs[7] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_2_[7]_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_121_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB9_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_3__1_sqmuxa ), .ALn(
        AFLSDF_INV_56_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(GND)
        , .Q(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_121_set_net_1 ));
    RGB \FCCC_0/GL1_INST/U0_RGB1  (.An(\FCCC_0/GL1_INST/U0_YNn ), .ENn(
        GND), .YL(), .YR(\FCCC_0/GL1_INST/U0_RGB1_YR ));
    SLE_IP_EN 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/FF_26  
        (.EN(VCC), .IPENn());
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_228_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_91_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_228_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_228_rs_net_1 ));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_177  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/MMUART1_RXD_F2H_SCP_net ), 
        .IPB(\hello_regs_MSS_0/MSS_ADLIB_INST/MGPIO20B_F2H_GPIN_net ), 
        .IPC());
    INV_BA AFLSDF_INV_90 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_75_net_1 ), .Y(
        AFLSDF_INV_90_net_1));
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_data_out8_55  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_3_[7]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_655 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_55_net_1 ));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_77  (.A(
        VCC), .B(VCC), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[11] ), 
        .IPB(
        \hello_regs_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[18] ), 
        .IPC());
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_242_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_18_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_242_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_242_rs_net_1 ));
    CFG2 #( .INIT(4'h2) )  \reg_apb_wrp_0/rd_enable_0_a2  (.A(N_637), 
        .B(CoreAPB3_0_APBmslave5_PWRITE), .Y(\reg_apb_wrp_0/rd_enable )
        );
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_49  (.A(
        GND), .B(VCC), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[3] ), .IPB(), 
        .IPC());
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_211_rs_RNI2RC71  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_107_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_211_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_13_rs[3] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_13_[3]_net_1 ));
    CFG3 #( .INIT(8'hF2) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_243  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_12_[3]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_644 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_243_i ));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_14_[6]  (.D(
        \CoreAPB3_0_APBmslave5_PWDATA[6] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB13_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_14__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_222_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_14_rs[6] ));
    RGB \FCCC_0/GL1_INST/U0_RGB1_RGB3  (.An(\FCCC_0/GL1_INST/U0_YNn ), 
        .ENn(GND), .YL(), .YR(
        \FCCC_0/GL1_INST/U0_RGB1_RGB3_rgbr_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_10_[7]  (.D(
        \CoreAPB3_0_APBmslave5_PWDATA[7] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB10_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_10__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_180_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_10_rs[7] ));
    CFG3 #( .INIT(8'hF2) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_189  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_5_[1]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_653 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_189_i ));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_58  (.A(
        VCC), .B(GND), .C(VCC), .IPA(), .IPB(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[19] ), .IPC());
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_192  (
        .A(GND), .B(VCC), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_AWID_HSEL0_net[0] ), .IPB(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[8] ), 
        .IPC(\hello_regs_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[20] )
        );
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_26_set_RNI647P  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_26_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_201_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_5_rs[7] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_5_[7]_net_1 ));
    CFG3 #( .INIT(8'hF2) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_222  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_14_[6]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_650 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_222_i ));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_47  (.A(
        VCC), .B(GND), .C(VCC), .IPA(), .IPB(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[1] ), .IPC());
    CFG3 #( .INIT(8'h80) )  
        \reg_apb_wrp_0/reg16x8_0/mem_3__1_sqmuxa_0_a2  (.A(
        \reg_apb_wrp_0/reg16x8_0/N_655 ), .B(N_637), .C(N_638), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_3__1_sqmuxa ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_94_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB5_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_11__1_sqmuxa ), .ALn(
        AFLSDF_INV_57_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(GND)
        , .Q(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_94_set_net_1 ));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_190_rs_RNIBI3N  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_72_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_190_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_9_rs[0] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_9_[0]_net_1 ));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_131  (
        .A(VCC), .B(GND), .C(VCC), .IPA(), .IPB(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[13] ), .IPC(
        ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_234_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_94_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_234_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_234_rs_net_1 ));
    CFG3 #( .INIT(8'hF2) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_194  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_9_[2]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_643 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_194_i ));
    CFG4 #( .INIT(16'h7530) )  
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_4[2]  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_6_[2]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/mem_3_[2]_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/N_655 ), .D(
        \reg_apb_wrp_0/reg16x8_0/N_652 ), .Y(
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_4[2]_net_1 ));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_172  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/MGPIO24B_F2H_GPIN_net ), .IPB(
        \hello_regs_MSS_0/MSS_ADLIB_INST/MMUART0_RTS_F2H_SCP_net ), 
        .IPC());
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_146  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/MGPIO0A_F2H_GPIN_net ), .IPB()
        , .IPC());
    CFG4 #( .INIT(16'h8000) )  
        \reg_apb_wrp_0/reg16x8_0/WRITE_GEN.mem_15__2_i_a2[5]  (.A(
        \CoreAPB3_0_APBmslave5_PADDR[2] ), .B(
        \CoreAPB3_0_APBmslave5_PADDR[5] ), .C(
        \CoreAPB3_0_APBmslave5_PADDR[4] ), .D(
        \CoreAPB3_0_APBmslave5_PADDR[3] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/N_654 ));
    INV_BA AFLSDF_INV_127 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_49_net_1 ), .Y(
        AFLSDF_INV_127_net_1));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_10_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB15_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_4__1_sqmuxa ), .ALn(
        AFLSDF_INV_58_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(GND)
        , .Q(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_10_set_net_1 ));
    CFG3 #( .INIT(8'hF2) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_150  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_0_[6]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_645 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_150_i ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_176_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_102_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_176_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_176_rs_net_1 ));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_159  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/SPI0_SS3_F2H_SCP_net ), .IPB(
        \hello_regs_MSS_0/MSS_ADLIB_INST/SPI0_SS1_F2H_SCP_net ), .IPC()
        );
    CFG3 #( .INIT(8'hF2) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_202  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_9_[6]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_643 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_202_i ));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_138_rs_RNIL15L  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_4_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_138_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_4_rs[2] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_4_[2]_net_1 ));
    CFG4 #( .INIT(16'h7530) )  
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_0_6[6]  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_4_[6]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/mem_1_[6]_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/N_651 ), .D(
        \reg_apb_wrp_0/reg16x8_0/N_648 ), .Y(
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_0_6[6]_net_1 ));
    CFG4 #( .INIT(16'h7530) )  
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_4[5]  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_6_[5]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/mem_3_[5]_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/N_655 ), .D(
        \reg_apb_wrp_0/reg16x8_0/N_652 ), .Y(
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_4[5]_net_1 ));
    INV_BA AFLSDF_INV_28 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_84_net_1 ), .Y(
        AFLSDF_INV_28_net_1));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_15  (.A(
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[20] ), .B(
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[27] ), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[20] ), .IPB(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[27] ), .IPC());
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_data_out8_93  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_11_[5]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_649 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_93_net_1 ));
    SLE_IP_EN 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/FF_29  
        (.EN(\hello_regs_MSS_0/MSS_ADLIB_INST_RNIUO3B/U0_RGB1_YR ), 
        .IPENn(AFLSDF_INV_59_net_1));
    CFG4 #( .INIT(16'h7530) )  
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_4[3]  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_6_[3]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/mem_3_[3]_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/N_655 ), .D(
        \reg_apb_wrp_0/reg16x8_0/N_652 ), .Y(
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_4[3]_net_1 ));
    CFG4 #( .INIT(16'h7530) )  
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_7[3]  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_8_[3]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/mem_5_[3]_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/N_653 ), .D(N_639), .Y(
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_7[3]_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_1_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB16_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_7__1_sqmuxa ), .ALn(
        AFLSDF_INV_60_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(GND)
        , .Q(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_1_set_net_1 ));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_276  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[0] ), 
        .IPB(
        \hello_regs_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[3] ), 
        .IPC(
        \hello_regs_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[15] ));
    CFG3 #( .INIT(8'hF2) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_250  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_15_[3]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_654 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_250_i ));
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_data_out8_25  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_2_[0]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_642 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_25_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_10_[2]  (.D(
        \CoreAPB3_0_APBmslave5_PWDATA[2] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB10_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_10__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_170_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_10_rs[2] ));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/mem_12__RNIL9951[5]  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_21_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_245_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_12_rs[5] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_12_[5]_net_1 ));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/mem_15__RNI16E11[1]  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_58_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_248_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_15_rs[1] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_15_[1]_net_1 ));
    CFG4 #( .INIT(16'hECA0) )  \CoreAPB3_0/u_mux_p_to_b3/PRDATA_0[23]  
        (.A(\CoreAPB3_0/u_mux_p_to_b3/N_636 ), .B(
        \COREAPBLSRAM_0.PRDATA4 ), .C(\COREAPBLSRAM_0.PRDATA_reg[23] ), 
        .D(\COREAPBLSRAM_0.lsram_width32_PRDATA[23] ), .Y(
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[23] ));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_121  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/FAB_AVALID_net ), .IPB(), 
        .IPC());
    INV_BA AFLSDF_INV_37 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_81_net_1 ), .Y(
        AFLSDF_INV_37_net_1));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_111_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB7_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_13__1_sqmuxa ), .ALn(
        AFLSDF_INV_61_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(GND)
        , .Q(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_111_set_net_1 ));
    CFG3 #( .INIT(8'hF2) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_213  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_13_[5]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_646 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_213_i ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_3_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB12_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_7__1_sqmuxa ), .ALn(
        AFLSDF_INV_62_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(GND)
        , .Q(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_3_set_net_1 ));
    SLE_IP_EN 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/FF_18  
        (.EN(VCC), .IPENn());
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_data_out8_39  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_2_[7]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_642 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_39_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_86_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB13_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_0__1_sqmuxa ), .ALn(
        AFLSDF_INV_63_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(GND)
        , .Q(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_86_set_net_1 ));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_198  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[2] ), 
        .IPB(\hello_regs_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[14] )
        , .IPC());
    INV_BA AFLSDF_INV_82 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_116_net_1 ), .Y(
        AFLSDF_INV_82_net_1));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_146_rs_RNI8OGH  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_83_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_146_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_0_rs[3] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_0_[3]_net_1 ));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_269  (
        .A(VCC), .B(GND), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[29] ), 
        .IPB(\hello_regs_MSS_0/MSS_ADLIB_INST/F_ARVALID_HWRITE1_net ), 
        .IPC());
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_data_out8_3  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_7_[6]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_641 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_3_net_1 ));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_210  (
        .A(VCC), .B(GND), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[28] ), 
        .IPB(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_AWLOCK_HMASTLOCK0_net[0] ), 
        .IPC());
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_39  (.A(
        GND), .B(GND), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[22] ), .IPB(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[29] ), .IPC());
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_201  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[5] ), 
        .IPB(\hello_regs_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[17] )
        , .IPC());
    CFG4 #( .INIT(16'h0001) )  
        \reg_apb_wrp_0/reg16x8_0/WRITE_GEN.mem_0__2_i_a2[3]  (.A(
        \CoreAPB3_0_APBmslave5_PADDR[2] ), .B(
        \CoreAPB3_0_APBmslave5_PADDR[5] ), .C(
        \CoreAPB3_0_APBmslave5_PADDR[4] ), .D(
        \CoreAPB3_0_APBmslave5_PADDR[3] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/N_645 ));
    SLE \reg_apb_wrp_0/reg16x8_0/data_out[3]  (.D(
        \reg_apb_wrp_0/reg16x8_0/N_37_i_0 ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB11_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/rd_enable ), .ALn(
        \hello_regs_MSS_0/MSS_ADLIB_INST_RNIUO3B/U0_RGB1_RGB3_rgbr_net_1 )
        , .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreAPB3_0_APBmslave5_PRDATA[3] ));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_42_set_RNI8DHT  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_42_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_157_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_1_rs[5] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_1_[5]_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_171_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_36_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_171_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_171_rs_net_1 ));
    CFG4 #( .INIT(16'h7350) )  
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_2[0]  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_12_[0]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/mem_9_[0]_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/N_644 ), .D(
        \reg_apb_wrp_0/reg16x8_0/N_643 ), .Y(
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_2[0]_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_74_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB19_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_9__1_sqmuxa ), .ALn(
        AFLSDF_INV_64_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(GND)
        , .Q(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_74_set_net_1 ));
    CFG4 #( .INIT(16'hFFB3) )  
        \CoreAPB3_0/u_mux_p_to_b3/PRDATA_0_iv_0[7]  (.A(
        \COREAPBLSRAM_0.lsram_width32_PRDATA[7] ), .B(
        \CoreAPB3_0/u_mux_p_to_b3/PRDATA_0_iv_0_1_0[7]_net_1 ), .C(
        \COREAPBLSRAM_0.PRDATA4 ), .D(
        \CoreAPB3_0/u_mux_p_to_b3/PRDATA_0_iv_0_0[7]_net_1 ), .Y(
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[7] ));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_178  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(), .IPB(
        \hello_regs_MSS_0/MSS_ADLIB_INST/MMUART0_DSR_F2H_SCP_net ), 
        .IPC());
    CFG4 #( .INIT(16'hFFFE) )  
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_12[5]  (.A(
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_1[5]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_3[5]_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_2[5]_net_1 ), .D(
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_0[5]_net_1 ), .Y(
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_12[5]_net_1 ));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_186  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/MGPIO29B_F2H_GPIN_net ), .IPB(
        ), .IPC());
    CFG4 #( .INIT(16'hECA0) )  \CoreAPB3_0/u_mux_p_to_b3/PRDATA_0[19]  
        (.A(\CoreAPB3_0/u_mux_p_to_b3/N_636 ), .B(
        \COREAPBLSRAM_0.PRDATA4 ), .C(\COREAPBLSRAM_0.PRDATA_reg[19] ), 
        .D(\COREAPBLSRAM_0.lsram_width32_PRDATA[19] ), .Y(
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[19] ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_56_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB15_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_15__1_sqmuxa ), .ALn(
        AFLSDF_INV_65_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(GND)
        , .Q(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_56_set_net_1 ));
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_data_out8_13  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_1_[2]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_651 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_13_net_1 ));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_37  (.A(
        GND), .B(VCC), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[20] ), .IPB(), 
        .IPC());
    INV_BA AFLSDF_INV_117 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_34_net_1 ), .Y(
        AFLSDF_INV_117_net_1));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_90  (.A(
        VCC), .B(VCC), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[31] ), 
        .IPB(\hello_regs_MSS_0/MSS_ADLIB_INST/RXDF_net[6] ), .IPC());
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_210_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_106_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_210_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_210_rs_net_1 ));
    SLE \COREAPBLSRAM_0/PRDATA_reg[18]  (.D(
        \COREAPBLSRAM_0.lsram_width32_PRDATA[18] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB8_rgbr_net_1 ), .EN(
        \COREAPBLSRAM_0.PRDATA4 ), .ALn(
        \hello_regs_MSS_0/MSS_ADLIB_INST_RNIUO3B/U0_RGB1_RGB0_rgbr_net_1 )
        , .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \COREAPBLSRAM_0.PRDATA_reg[18] ));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_71_set_RNIN5AJ  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_71_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_188_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_8_rs[7] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_8_[7]_net_1 ));
    CFG3 #( .INIT(8'hF2) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_154  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_1_[2]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_651 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_154_i ));
    CFG4 #( .INIT(16'h7350) )  
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_2[4]  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_12_[4]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/mem_9_[4]_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/N_644 ), .D(
        \reg_apb_wrp_0/reg16x8_0/N_643 ), .Y(
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_2[4]_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/data_out[5]  (.D(
        \reg_apb_wrp_0/reg16x8_0/N_82_i_0 ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB10_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/rd_enable ), .ALn(
        \hello_regs_MSS_0/MSS_ADLIB_INST_RNIUO3B/U0_RGB1_RGB2_rgbr_net_1 )
        , .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreAPB3_0_APBmslave5_PRDATA[5] ));
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_data_out8_42  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_1_[5]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_651 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_42_net_1 ));
    CFG3 #( .INIT(8'hF2) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_255  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_15_[4]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_654 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_255_i ));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_268  (
        .A(VCC), .B(\FCCC_0/GL1_INST/U0_RGB1_YR ), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[28] ), 
        .IPB(\hello_regs_MSS_0/MSS_ADLIB_INST/CLK_BASE_net ), .IPC());
    SLE \COREAPBLSRAM_0/PRDATA_reg[12]  (.D(
        \COREAPBLSRAM_0.lsram_width32_PRDATA[12] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB9_rgbr_net_1 ), .EN(
        \COREAPBLSRAM_0.PRDATA4 ), .ALn(
        \hello_regs_MSS_0/MSS_ADLIB_INST_RNIUO3B/U0_RGB1_RGB1_rgbr_net_1 )
        , .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \COREAPBLSRAM_0.PRDATA_reg[12] ));
    INV_BA AFLSDF_INV_39 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_93_net_1 ), .Y(
        AFLSDF_INV_39_net_1));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_63_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB12_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_15__1_sqmuxa ), .ALn(
        AFLSDF_INV_66_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(GND)
        , .Q(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_63_set_net_1 ));
    CFG3 #( .INIT(8'hF2) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_228  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_11_[3]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_649 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_228_i ));
    CFG4 #( .INIT(16'hFF80) )  
        \CoreAPB3_0/u_mux_p_to_b3/PRDATA_0_iv_0_0[1]  (.A(N_639), .B(
        \GPIO_OUT_1_c[1] ), .C(
        \CoreAPB3_0.u_mux_p_to_b3.PRDATA_0_iv_0_a2_3_5[1] ), .D(
        \CoreAPB3_0/u_mux_p_to_b3/N_584 ), .Y(
        \CoreAPB3_0/u_mux_p_to_b3/PRDATA_0_iv_0_0[1]_net_1 ));
    INV_BA AFLSDF_INV_23 (.A(AFLSDF_INV_23_net_1), .Y(
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/A_DOUT_CLK_net )
        );
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_201_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_26_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_201_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_201_rs_net_1 ));
    CFG4 #( .INIT(16'h7530) )  
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_6[7]  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_4_[7]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/mem_1_[7]_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/N_651 ), .D(
        \reg_apb_wrp_0/reg16x8_0/N_648 ), .Y(
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_6[7]_net_1 ));
    CFG4 #( .INIT(16'hFFB3) )  
        \CoreAPB3_0/u_mux_p_to_b3/PRDATA_0_iv_0[5]  (.A(
        \COREAPBLSRAM_0.lsram_width32_PRDATA[5] ), .B(
        \CoreAPB3_0/u_mux_p_to_b3/PRDATA_0_iv_0_1_0[5]_net_1 ), .C(
        \COREAPBLSRAM_0.PRDATA4 ), .D(
        \CoreAPB3_0/u_mux_p_to_b3/PRDATA_0_iv_0_0[5]_net_1 ), .Y(
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[5] ));
    CFG3 #( .INIT(8'hF2) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_227  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_7_[4]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_641 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_227_i ));
    CFG3 #( .INIT(8'hF2) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_199  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_5_[6]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_653 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_199_i ));
    CFG2_IP_BC 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/CFG_31  
        (.B(\CoreAPB3_0_APBmslave5_PWDATA[31] ), .C(
        \CoreAPB3_0_APBmslave5_PADDR[7] ), .IPB(
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/B_DIN_net[16] )
        , .IPC(
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/B_ADDR_net[12] )
        );
    CFG4 #( .INIT(16'hECA0) )  \CoreAPB3_0/u_mux_p_to_b3/PRDATA_0[26]  
        (.A(\CoreAPB3_0/u_mux_p_to_b3/N_636 ), .B(
        \COREAPBLSRAM_0.PRDATA4 ), .C(\COREAPBLSRAM_0.PRDATA_reg[26] ), 
        .D(\COREAPBLSRAM_0.lsram_width32_PRDATA[26] ), .Y(
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[26] ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_246_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_22_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_246_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_246_rs_net_1 ));
    IP_INTERFACE ip_interface_inst (.A(VCC), .B(ff_to_start_net), .C(
        VCC), .IPA(), .IPB(), .IPC());
    CFG4 #( .INIT(16'h7530) )  
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_3[1]  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_2_[1]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/mem_13_[1]_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/N_646 ), .D(
        \reg_apb_wrp_0/reg16x8_0/N_642 ), .Y(
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_3[1]_net_1 ));
    RGB \FCCC_0/GL1_INST/U0_RGB1_RGB12  (.An(
        \FCCC_0/GL1_INST/U0_YNn_GSouth ), .ENn(GND), .YL(
        \FCCC_0/GL1_INST/U0_RGB1_RGB12_rgbl_net_1 ), .YR(
        \FCCC_0/GL1_INST/U0_RGB1_RGB12_rgbr_net_1 ));
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_data_out8_40  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_1_[4]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_651 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_40_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_160_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_25_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_160_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_160_rs_net_1 ));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_214  (
        .A(GND), .B(GND), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_AWSIZE_HSIZE0_net[0] ), 
        .IPB(\hello_regs_MSS_0/MSS_ADLIB_INST/F_WID_HREADY01_net[2] ), 
        .IPC());
    INV_BA AFLSDF_INV_56 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_121_net_1 ), .Y(
        AFLSDF_INV_56_net_1));
    CFG3 #( .INIT(8'hF2) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_208  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_13_[0]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_646 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_208_i ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_138_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_4_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_138_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_138_rs_net_1 ));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_143  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(), .IPB(
        \hello_regs_MSS_0/MSS_ADLIB_INST/FAB_M3_RESET_N_net ), .IPC());
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_241_rs_RNIDGQV  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_66_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_241_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_8_rs[3] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_8_[3]_net_1 ));
    CFG3 #( .INIT(8'hF2) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_207  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_6_[2]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_652 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_207_i ));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_5_[1]  (.D(
        \CoreAPB3_0_APBmslave5_PWDATA[1] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB9_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_5__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_189_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_5_rs[1] ));
    CFG4 #( .INIT(16'h7530) )  
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_7[0]  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_8_[0]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/mem_5_[0]_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/N_653 ), .D(N_639), .Y(
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_7[0]_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_11_[7]  (.D(
        \CoreAPB3_0_APBmslave5_PWDATA[7] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB5_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_11__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_236_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_11_rs[7] ));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_20  (.A(
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[25] ), .B(GND), .C(
        VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[25] ), .IPB(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_MASTLOCK_net ), .IPC());
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_97_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB7_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_10__1_sqmuxa ), .ALn(
        AFLSDF_INV_67_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(GND)
        , .Q(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_97_set_net_1 ));
    CFG3 #( .INIT(8'hF2) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_167  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_2_[7]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_642 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_167_i ));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_0_[6]  (.D(
        \CoreAPB3_0_APBmslave5_PWDATA[6] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB13_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_0__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_150_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_0_rs[6] ));
    INV_BA AFLSDF_INV_81 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_95_net_1 ), .Y(
        AFLSDF_INV_81_net_1));
    IP_INTERFACE \FCCC_0/CCC_INST/IP_INTERFACE_0  (.A(VCC), .B(VCC), 
        .C(VCC), .IPA(\FCCC_0/CCC_INST/CLK0_net ), .IPB(
        \FCCC_0/CCC_INST/PSEL_net ), .IPC());
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_245_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_21_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_245_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_245_rs_net_1 ));
    CFG4 #( .INIT(16'hECA0) )  \CoreAPB3_0/u_mux_p_to_b3/PRDATA_0[31]  
        (.A(\CoreAPB3_0/u_mux_p_to_b3/N_636 ), .B(
        \COREAPBLSRAM_0.PRDATA4 ), .C(\COREAPBLSRAM_0.PRDATA_reg[31] ), 
        .D(\COREAPBLSRAM_0.lsram_width32_PRDATA[31] ), .Y(
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[31] ));
    SLE \COREAPBLSRAM_0/PRDATA_reg[9]  (.D(
        \COREAPBLSRAM_0.lsram_width32_PRDATA[9] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB11_rgbr_net_1 ), .EN(
        \COREAPBLSRAM_0.PRDATA4 ), .ALn(
        \hello_regs_MSS_0/MSS_ADLIB_INST_RNIUO3B/U0_RGB1_RGB3_rgbr_net_1 )
        , .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \COREAPBLSRAM_0.PRDATA_reg[9] ));
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_data_out8_35  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_2_[5]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_642 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_35_net_1 ));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_104  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/RCGF_net[4] ), .IPB(
        \hello_regs_MSS_0/MSS_ADLIB_INST/FAB_LINESTATE_net[0] ), .IPC()
        );
    CFG3 #( .INIT(8'hF2) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_226  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_11_[2]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_649 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_226_i ));
    sdf_IOPAD_IN \hello_regs_MSS_0/MMUART_0_RXD_PAD/U_IOPAD  (.PAD(
        MMUART_0_RXD), .Y(\hello_regs_MSS_0/MMUART_0_RXD_PAD_Y ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_227_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_52_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_227_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_227_rs_net_1 ));
    CFG1_IP_B 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/CFG_10  
        (.B(\CoreAPB3_0_APBmslave5_PWDATA[10] ), .IPB(
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/A_DIN_net[11] )
        );
    CFG4 #( .INIT(16'hECA0) )  \CoreAPB3_0/u_mux_p_to_b3/PRDATA_0[10]  
        (.A(\CoreAPB3_0/u_mux_p_to_b3/N_636 ), .B(
        \COREAPBLSRAM_0.PRDATA4 ), .C(\COREAPBLSRAM_0.PRDATA_reg[10] ), 
        .D(\COREAPBLSRAM_0.lsram_width32_PRDATA[10] ), .Y(
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[10] ));
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_data_out8_68  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_8_[4]_net_1 ), .B(N_639), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_68_net_1 ));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_262  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[10] ), 
        .IPB(\hello_regs_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[22] )
        , .IPC());
    INV_BA AFLSDF_INV_25 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_119_net_1 ), .Y(
        AFLSDF_INV_25_net_1));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_259  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[7] ), 
        .IPB(\hello_regs_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[19] )
        , .IPC());
    CFG2_IP_BC 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/CFG_0  
        (.B(\CoreAPB3_0_APBmslave5_PWDATA[0] ), .C(GND), .IPB(
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/A_DIN_net[0] )
        , .IPC(
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/A_ADDR_net[0] )
        );
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_263  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[11] ), 
        .IPB(\hello_regs_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[23] )
        , .IPC());
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_40_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB15_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_1__1_sqmuxa ), .ALn(
        AFLSDF_INV_68_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(GND)
        , .Q(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_40_set_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_10_[1]  (.D(
        \CoreAPB3_0_APBmslave5_PWDATA[1] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB10_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_10__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_168_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_10_rs[1] ));
    INV_BA AFLSDF_INV_145 (.A(AFLSDF_INV_145_net_1), .Y(
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/B_DOUT_EN_net )
        );
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_209_rs_RNI55JJ  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_105_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_209_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_13_rs[1] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_13_[1]_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_118_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB13_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_14__1_sqmuxa ), .ALn(
        AFLSDF_INV_69_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(GND)
        , .Q(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_118_set_net_1 ));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_187_rs_RNI7LTR  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_12_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_187_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_5_rs[0] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_5_[0]_net_1 ));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_10_set_RNI9A5D  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_10_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_185_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_4_rs[7] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_4_[7]_net_1 ));
    CFG2_IP_BC 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/CFG_6  
        (.B(\CoreAPB3_0_APBmslave5_PWDATA[9] ), .C(GND), .IPB(
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/A_DIN_net[10] )
        , .IPC(
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/A_ADDR_net[3] )
        );
    IP_INTERFACE \FCCC_0/CCC_INST/IP_INTERFACE_13  (.A(VCC), .B(VCC), 
        .C(VCC), .IPA(\FCCC_0/CCC_INST/NGMUX1_ARST_N_net ), .IPB(), 
        .IPC(\FCCC_0/CCC_INST/PADDR_net[3] ));
    IP_INTERFACE \FCCC_0/CCC_INST/IP_INTERFACE_11  (.A(VCC), .B(VCC), 
        .C(VCC), .IPA(\FCCC_0/CCC_INST/PLL_POWERDOWN_N_net ), .IPB(
        \FCCC_0/CCC_INST/NGMUX3_HOLD_N_net ), .IPC());
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_22_set_RNIOHIQ  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_22_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_246_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_12_rs[6] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_12_[6]_net_1 ));
    CFG3 #( .INIT(8'hF2) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_206  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_10_[0]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_647 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_206_i ));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_3_[6]  (.D(
        \CoreAPB3_0_APBmslave5_PWDATA[6] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB11_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_3__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_134_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_3_rs[6] ));
    CFG2_IP_BC 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/CFG_20  
        (.B(\CoreAPB3_0_APBmslave5_PWDATA[5] ), .C(
        \COREAPBLSRAM_0/wen ), .IPB(
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/A_DIN_net[5] )
        , .IPC(
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/A_WEN_net[0] )
        );
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_91_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB6_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_11__1_sqmuxa ), .ALn(
        AFLSDF_INV_70_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(GND)
        , .Q(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_91_set_net_1 ));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_153_rs_RNIS90M  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_11_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_153_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_1_rs[1] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_1_[1]_net_1 ));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_258  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[6] ), 
        .IPB(\hello_regs_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[18] )
        , .IPC());
    SLE \COREAPBLSRAM_0/PRDATA_reg[27]  (.D(
        \COREAPBLSRAM_0.lsram_width32_PRDATA[27] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB8_rgbr_net_1 ), .EN(
        \COREAPBLSRAM_0.PRDATA4 ), .ALn(
        \hello_regs_MSS_0/MSS_ADLIB_INST_RNIUO3B/U0_RGB1_RGB0_rgbr_net_1 )
        , .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \COREAPBLSRAM_0.PRDATA_reg[27] ));
    SLE_IP_EN 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/FF_6  
        (.EN(VCC), .IPENn(AFLSDF_INV_71_net_1));
    CFG3 #( .INIT(8'hF2) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_159  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_1_[7]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_651 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_159_i ));
    INV_BA AFLSDF_INV_136 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_21_net_1 ), .Y(
        AFLSDF_INV_136_net_1));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_11_[2]  (.D(
        \CoreAPB3_0_APBmslave5_PWDATA[2] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB5_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_11__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_226_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_11_rs[2] ));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_65_set_RNI7LEV  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_65_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_140_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_4_rs[4] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_4_[4]_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_82_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB14_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_0__1_sqmuxa ), .ALn(
        AFLSDF_INV_72_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(GND)
        , .Q(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_82_set_net_1 ));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_183  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/MMUART0_TXD_F2H_SCP_net ), 
        .IPB(\hello_regs_MSS_0/MSS_ADLIB_INST/MMUART0_RI_F2H_SCP_net ), 
        .IPC());
    SLE \reg_apb_wrp_0/reg16x8_0/mem_7_[6]  (.D(
        \CoreAPB3_0_APBmslave5_PWDATA[6] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB12_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_7__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_231_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_7_rs[6] ));
    CFG4 #( .INIT(16'hECA0) )  \CoreAPB3_0/u_mux_p_to_b3/PRDATA_0[24]  
        (.A(\CoreAPB3_0/u_mux_p_to_b3/N_636 ), .B(
        \COREAPBLSRAM_0.PRDATA4 ), .C(\COREAPBLSRAM_0.PRDATA_reg[24] ), 
        .D(\COREAPBLSRAM_0.lsram_width32_PRDATA[24] ), .Y(
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[24] ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_147_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_80_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_147_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_147_rs_net_1 ));
    INV_BA AFLSDF_INV_34 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_104_net_1 ), .Y(
        AFLSDF_INV_34_net_1));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_80  (.A(
        VCC), .B(VCC), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[14] ), 
        .IPB(
        \hello_regs_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[21] ), 
        .IPC());
    CFG3 #( .INIT(8'hF2) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_233  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_7_[7]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_641 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_233_i ));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_237  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[35] ), 
        .IPB(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[47] ), 
        .IPC());
    RGB \hello_regs_MSS_0/MSS_ADLIB_INST_RNIUO3B/U0_RGB1_RGB5  (.An(
        \hello_regs_MSS_0/MSS_ADLIB_INST_RNIUO3B/U0_YNn_GSouth ), .ENn(
        GND), .YL(), .YR(
        \hello_regs_MSS_0/MSS_ADLIB_INST_RNIUO3B/U0_RGB1_RGB5_rgbr_net_1 )
        );
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_152_rs_RNIHTAV  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_9_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_152_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_1_rs[0] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_1_[0]_net_1 ));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_29_set_RNI7L49  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_29_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_162_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_2_rs[2] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_2_[2]_net_1 ));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_156_rs_RNI41241  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_40_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_156_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_1_rs[4] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_1_[4]_net_1 ));
    INV_BA AFLSDF_INV_134 (.A(AFLSDF_INV_134_net_1), .Y(
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/A_DOUT_SRST_N_net )
        );
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_224_rs_RNIRK1N  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_89_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_224_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_11_rs[1] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_11_[1]_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_144_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_81_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_144_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_144_rs_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_77_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB14_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_9__1_sqmuxa ), .ALn(
        AFLSDF_INV_73_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(GND)
        , .Q(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_77_set_net_1 ));
    CFG3 #( .INIT(8'hF2) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_229  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_7_[5]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_641 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_229_i ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[5].APB_8.GPOUT_reg[5]  (.D(
        \CoreAPB3_0_APBmslave5_PWDATA[5] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB12_rgbr_net_1 ), .EN(
        \CoreGPIO_0/GPOUT_reg35 ), .ALn(
        \hello_regs_MSS_0/MSS_ADLIB_INST_RNIUO3B/U0_RGB1_RGB4_rgbr_net_1 )
        , .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \GPIO_OUT_1_c[5] ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_52_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB15_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_7__1_sqmuxa ), .ALn(
        AFLSDF_INV_74_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(GND)
        , .Q(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_52_set_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_8_[6]  (.D(
        \CoreAPB3_0_APBmslave5_PWDATA[6] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB5_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_8__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_186_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_8_rs[6] ));
    CFG3 #( .INIT(8'hF2) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_146  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_0_[3]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_645 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_146_i ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_126_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB16_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_7__1_sqmuxa ), .ALn(
        AFLSDF_INV_75_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(GND)
        , .Q(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_126_set_net_1 ));
    INV_BA AFLSDF_INV_131 (.A(AFLSDF_INV_131_net_1), .Y(
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/B_CLK_net )
        );
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_169_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_34_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_169_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_169_rs_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_13_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB15_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_1__1_sqmuxa ), .ALn(
        AFLSDF_INV_76_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(GND)
        , .Q(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_13_set_net_1 ));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_45_set_RNIJPKR  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_45_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_197_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_5_rs[5] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_5_[5]_net_1 ));
    CFG4 #( .INIT(16'h7350) )  
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_2[1]  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_12_[1]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/mem_9_[1]_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/N_644 ), .D(
        \reg_apb_wrp_0/reg16x8_0/N_643 ), .Y(
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_2[1]_net_1 ));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_53  (.A(
        GND), .B(GND), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[7] ), .IPB(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[14] ), .IPC());
    SLE \reg_apb_wrp_0/reg16x8_0/data_out[0]  (.D(
        \reg_apb_wrp_0/reg16x8_0/N_7_i_0 ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB11_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/rd_enable ), .ALn(
        \hello_regs_MSS_0/MSS_ADLIB_INST_RNIUO3B/U0_RGB1_RGB3_rgbr_net_1 )
        , .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreAPB3_0_APBmslave5_PRDATA[0] ));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_149  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/I2C1_SCL_F2H_SCP_net ), .IPB(
        \hello_regs_MSS_0/MSS_ADLIB_INST/MGPIO5A_F2H_GPIN_net ), .IPC()
        );
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_252  (
        .A(VCC), .B(VCC), .C(GND), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[0] ), 
        .IPB(\hello_regs_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[12] )
        , .IPC(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_ARSIZE_HSIZE1_net[0] ));
    CFG4 #( .INIT(16'h7530) )  
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_6[0]  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_4_[0]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/mem_1_[0]_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/N_651 ), .D(
        \reg_apb_wrp_0/reg16x8_0/N_648 ), .Y(
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_6[0]_net_1 ));
    CFG3 #( .INIT(8'hF2) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_209  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_13_[1]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_646 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_209_i ));
    CFG3 #( .INIT(8'hF2) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_176  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_10_[5]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_647 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_176_i ));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_253  (
        .A(VCC), .B(VCC), .C(GND), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[1] ), 
        .IPB(\hello_regs_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[13] )
        , .IPC(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_ARSIZE_HSIZE1_net[1] ));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_4_[6]  (.D(
        \CoreAPB3_0_APBmslave5_PWDATA[6] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB15_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_4__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_143_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_4_rs[6] ));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_227  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[11] ), 
        .IPB(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[23] ), 
        .IPC());
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_data_out8_84  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_0_[4]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_645 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_84_net_1 ));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_14  (.A(
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[19] ), .B(VCC), .C(
        VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[19] ), .IPB(), 
        .IPC());
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/mem_14__RNIAK9M[3]  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_115_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_219_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_14_rs[3] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_14_[3]_net_1 ));
    INV_BA AFLSDF_INV_22 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_108_net_1 ), .Y(
        AFLSDF_INV_22_net_1));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_219_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_115_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_219_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_219_rs_net_1 ));
    IP_INTERFACE \FCCC_0/CCC_INST/IP_INTERFACE_16  (.A(VCC), .B(VCC), 
        .C(VCC), .IPA(), .IPB(\FCCC_0/CCC_INST/GPD2_ARST_N_net ), .IPC(
        \FCCC_0/CCC_INST/PADDR_net[6] ));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_6_[6]  (.D(
        \CoreAPB3_0_APBmslave5_PWDATA[6] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB12_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_6__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_175_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_6_rs[6] ));
    IOTRI_OB_EB \GPIO_OUT_1_obuf[0]/U0/U_IOTRI  (.D(\GPIO_OUT_1_c[0] ), 
        .E(VCC), .DOUT(\GPIO_OUT_1_obuf[0]/U0/DOUT1 ), .EOUT(
        \GPIO_OUT_1_obuf[0]/U0/EOUT1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_71_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB7_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_8__1_sqmuxa ), .ALn(
        AFLSDF_INV_77_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(GND)
        , .Q(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_71_set_net_1 ));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/mem_3__RNI429V[5]  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_51_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_133_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_3_rs[5] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_3_[5]_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_98_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB10_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_10__1_sqmuxa ), .ALn(
        AFLSDF_INV_78_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(GND)
        , .Q(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_98_set_net_1 ));
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_data_out8_69  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_8_[5]_net_1 ), .B(N_639), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_69_net_1 ));
    CFG4 #( .INIT(16'h7530) )  
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_3[4]  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_2_[4]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/mem_13_[4]_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/N_646 ), .D(
        \reg_apb_wrp_0/reg16x8_0/N_642 ), .Y(
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_3[4]_net_1 ));
    IOENFF_BYPASS \GPIO_OUT_1_obuf[6]/U0/U_IOENFF  (.A(
        \GPIO_OUT_1_obuf[6]/U0/EOUT1 ), .Y(
        \GPIO_OUT_1_obuf[6]/U0/EOUT ));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_1_[1]  (.D(
        \CoreAPB3_0_APBmslave5_PWDATA[1] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB17_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_1__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_153_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_1_rs[1] ));
    CFG4 #( .INIT(16'hFFFE) )  
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_13[0]  (.A(
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_4[0]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_5[0]_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_7[0]_net_1 ), .D(
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_6[0]_net_1 ), .Y(
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_13[0]_net_1 ));
    sdf_IOPAD_TRI \GPIO_OUT_1_obuf[2]/U0/U_IOPAD  (.PAD(GPIO_OUT_1[2]), 
        .D(\GPIO_OUT_1_obuf[2]/U0/DOUT ), .E(
        \GPIO_OUT_1_obuf[2]/U0/EOUT ));
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_data_out8_6  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_4_[3]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_648 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_6_net_1 ));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_260  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[8] ), 
        .IPB(\hello_regs_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[20] )
        , .IPC());
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_data_out8_96  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_10_[3]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_647 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_96_net_1 ));
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_data_out8_87  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_0_[7]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_645 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_87_net_1 ));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/mem_10__RNI19QJ[1]  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_98_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_168_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_10_rs[1] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_10_[1]_net_1 ));
    GB \hello_regs_MSS_0/MSS_ADLIB_INST_RNIUO3B  (.An(
        AFLSDF_INV_79_net_1), .ENn(GND), .YNn(
        \hello_regs_MSS_0/MSS_ADLIB_INST_RNIUO3B/U0_YNn ), .YSn(
        \hello_regs_MSS_0/MSS_ADLIB_INST_RNIUO3B/U0_YNn_GSouth ));
    CFG3 #( .INIT(8'hF2) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_185  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_4_[7]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_648 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_185_i ));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_52  (.A(
        GND), .B(GND), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[6] ), .IPB(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[13] ), .IPC());
    SLE_IP_EN 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/FF_16  
        (.EN(VCC), .IPENn());
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/mem_6__RNIB1OQ[4]  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_36_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_171_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_6_rs[4] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_6_[4]_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_124_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB15_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_7__1_sqmuxa ), .ALn(
        AFLSDF_INV_80_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(GND)
        , .Q(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_124_set_net_1 ));
    SLE \COREAPBLSRAM_0/PRDATA_reg[4]  (.D(
        \COREAPBLSRAM_0.lsram_width32_PRDATA[4] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB10_rgbr_net_1 ), .EN(
        \COREAPBLSRAM_0.PRDATA4 ), .ALn(
        \hello_regs_MSS_0/MSS_ADLIB_INST_RNIUO3B/U0_RGB1_RGB2_rgbr_net_1 )
        , .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \COREAPBLSRAM_0.PRDATA_reg[4] ));
    CFG4 #( .INIT(16'h7530) )  
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_6[5]  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_4_[5]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/mem_1_[5]_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/N_651 ), .D(
        \reg_apb_wrp_0/reg16x8_0/N_648 ), .Y(
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_6[5]_net_1 ));
    INV_BA AFLSDF_INV_78 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_98_net_1 ), .Y(
        AFLSDF_INV_78_net_1));
    CFG3 #( .INIT(8'h02) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_116  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_14_[4]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_650 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_116_net_1 ));
    CFG4 #( .INIT(16'h7350) )  
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_1[5]  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_15_[5]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/mem_14_[5]_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/N_654 ), .D(
        \reg_apb_wrp_0/reg16x8_0/N_650 ), .Y(
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_1[5]_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_143_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_8_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_143_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_143_rs_net_1 ));
    CFG3 #( .INIT(8'h80) )  
        \reg_apb_wrp_0/reg16x8_0/mem_6__1_sqmuxa_0_a2_0_a2  (.A(
        \reg_apb_wrp_0/reg16x8_0/N_652 ), .B(N_637), .C(N_638), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_6__1_sqmuxa ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_95_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB5_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_11__1_sqmuxa ), .ALn(
        AFLSDF_INV_81_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(GND)
        , .Q(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_95_set_net_1 ));
    CFG3 #( .INIT(8'hF2) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_183  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_7_[2]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_641 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_183_i ));
    CFG3 #( .INIT(8'h80) )  
        \reg_apb_wrp_0/reg16x8_0/mem_7__1_sqmuxa_0_a2  (.A(
        \reg_apb_wrp_0/reg16x8_0/N_641 ), .B(N_637), .C(N_638), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_7__1_sqmuxa ));
    CFG2 #( .INIT(4'h1) )  \reg_apb_wrp_0/reg16x8_0/data_out_RNO[3]  (
        .A(\reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_13[3]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_12[3]_net_1 ), .Y(
        \reg_apb_wrp_0/reg16x8_0/N_37_i_0 ));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_69  (.A(
        GND), .B(VCC), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[30] ), .IPB(
        \hello_regs_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[3] ), 
        .IPC());
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_203_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_28_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_203_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_203_rs_net_1 ));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_106_set_RNIVI321  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_106_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_210_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_13_rs[2] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_13_[2]_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_11_[1]  (.D(
        \CoreAPB3_0_APBmslave5_PWDATA[1] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB5_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_11__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_224_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_11_rs[1] ));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_100  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/RCGF_net[0] ), .IPB(
        \hello_regs_MSS_0/MSS_ADLIB_INST/RCGF_net[7] ), .IPC());
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_116_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB11_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_14__1_sqmuxa ), .ALn(
        AFLSDF_INV_82_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(GND)
        , .Q(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_116_set_net_1 ));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_189  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/I2C0_SDA_F2H_SCP_net ), .IPB()
        , .IPC());
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_64_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB7_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_8__1_sqmuxa ), .ALn(
        AFLSDF_INV_83_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(GND)
        , .Q(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_64_set_net_1 ));
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_data_out8_52  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_7_[4]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_641 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_52_net_1 ));
    CFG3 #( .INIT(8'hF2) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_241  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_8_[3]_net_1 ), .B(N_639), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_241_i ));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_109_set_RNI8BV11  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_109_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_213_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_13_rs[5] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_13_[5]_net_1 ));
    CFG3 #( .INIT(8'h80) )  
        \reg_apb_wrp_0/reg16x8_0/mem_1__1_sqmuxa_0_a2  (.A(
        \reg_apb_wrp_0/reg16x8_0/N_651 ), .B(N_637), .C(N_638), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_1__1_sqmuxa ));
    CFG4 #( .INIT(16'h7530) )  
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_7[2]  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_8_[2]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/mem_5_[2]_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/N_653 ), .D(N_639), .Y(
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_7[2]_net_1 ));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/mem_6__RNIRB1M[6]  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_120_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_175_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_6_rs[6] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_6_[6]_net_1 ));
    CFG4 #( .INIT(16'h0200) )  
        \reg_apb_wrp_0/reg16x8_0/WRITE_GEN.mem_3__2_i_a2[1]  (.A(
        \CoreAPB3_0_APBmslave5_PADDR[2] ), .B(
        \CoreAPB3_0_APBmslave5_PADDR[5] ), .C(
        \CoreAPB3_0_APBmslave5_PADDR[4] ), .D(
        \CoreAPB3_0_APBmslave5_PADDR[3] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/N_655 ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_230_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_92_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_230_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_230_rs_net_1 ));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_225_rs_RNI7J5K  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_50_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_225_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_7_rs[3] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_7_[3]_net_1 ));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_18  (.A(
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[23] ), .B(
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[30] ), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[23] ), .IPB(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[30] ), .IPC());
    CFG4 #( .INIT(16'h7350) )  
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_1[3]  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_15_[3]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/mem_14_[3]_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/N_654 ), .D(
        \reg_apb_wrp_0/reg16x8_0/N_650 ), .Y(
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_1[3]_net_1 ));
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_data_out8_81  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_0_[1]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_645 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_81_net_1 ));
    CFG2 #( .INIT(4'h7) )  
        \CoreAPB3_0/u_mux_p_to_b3/PRDATA_0_iv_0_1_0[2]  (.A(N_637), .B(
        \CoreAPB3_0_APBmslave5_PRDATA[2] ), .Y(
        \CoreAPB3_0/u_mux_p_to_b3/PRDATA_0_iv_0_1_0[2]_net_1 ));
    INV_BA AFLSDF_INV_132 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_27_net_1 ), .Y(
        AFLSDF_INV_132_net_1));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_67  (.A(
        GND), .B(VCC), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[28] ), .IPB(
        \hello_regs_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[1] ), 
        .IPC());
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_205  (
        .A(VCC), .B(GND), .C(GND), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[23] ), 
        .IPB(\hello_regs_MSS_0/MSS_ADLIB_INST/F_AWLEN_HBURST0_net[1] ), 
        .IPC(\hello_regs_MSS_0/MSS_ADLIB_INST/F_WLAST_net ));
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_data_out8_16  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_12_[0]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_644 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_16_net_1 ));
    CFG4 #( .INIT(16'hFFFE) )  
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_13[5]  (.A(
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_4[5]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_5[5]_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_7[5]_net_1 ), .D(
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_6[5]_net_1 ), .Y(
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_13[5]_net_1 ));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_264  (
        .A(VCC), .B(GND), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[24] ), 
        .IPB(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_ARBURST_HTRANS1_net[0] ), 
        .IPC(\hello_regs_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PENABLE_net )
        );
    INV_BA AFLSDF_INV_21 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_22_net_1 ), .Y(
        AFLSDF_INV_21_net_1));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_136  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/SMBSUS_NI0_net ), .IPB(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_DMAREADY_net[0] ), .IPC());
    CFG3 #( .INIT(8'hF2) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_188  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_8_[7]_net_1 ), .B(N_639), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_188_i ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_30_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB10_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_6__1_sqmuxa ), .ALn(
        AFLSDF_INV_84_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(GND)
        , .Q(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_30_set_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_187_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_12_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_187_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_187_rs_net_1 ));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_41_set_RNI9RFM  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_41_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_193_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_5_rs[3] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_5_[3]_net_1 ));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_105  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/RCGF_net[5] ), .IPB(
        \hello_regs_MSS_0/MSS_ADLIB_INST/FAB_LINESTATE_net[1] ), .IPC()
        );
    INV_BA AFLSDF_INV_126 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_37_net_1 ), .Y(
        AFLSDF_INV_126_net_1));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_78_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB16_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_9__1_sqmuxa ), .ALn(
        AFLSDF_INV_85_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(GND)
        , .Q(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_78_set_net_1 ));
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_data_out8_50  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_7_[3]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_641 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_50_net_1 ));
    INV_BA AFLSDF_INV_50 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_55_net_1 ), .Y(
        AFLSDF_INV_50_net_1));
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_data_out8_65  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_4_[4]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_648 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_65_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_184_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_69_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_184_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_184_rs_net_1 ));
    SLE_IP_EN 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/FF_19  
        (.EN(VCC), .IPENn());
    CFG2 #( .INIT(4'h1) )  \reg_apb_wrp_0/reg16x8_0/data_out_RNO[0]  (
        .A(\reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_13[0]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_12[0]_net_1 ), .Y(
        \reg_apb_wrp_0/reg16x8_0/N_7_i_0 ));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_107  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(), .IPB(
        \hello_regs_MSS_0/MSS_ADLIB_INST/FAB_RXVALID_net ), .IPC());
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB12_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_4__1_sqmuxa ), .ALn(
        AFLSDF_INV_86_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(GND)
        , .Q(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_set_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_99_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB11_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_10__1_sqmuxa ), .ALn(
        AFLSDF_INV_87_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(GND)
        , .Q(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_99_set_net_1 ));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_70  (.A(
        VCC), .B(VCC), .C(VCC), .IPA(), .IPB(
        \hello_regs_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[4] ), 
        .IPC());
    CFG4 #( .INIT(16'h8000) )  
        \CoreAPB3_0/u_mux_p_to_b3/PRDATA_0_iv_0_a2_3_5[1]  (.A(
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PADDR[18] ), .B(
        hello_regs_MSS_0_FIC_0_APB_MASTER_PSELx), .C(
        \CoreAPB3_0/u_mux_p_to_b3/PRDATA_0_iv_0_a2_3_5_4[1]_net_1 ), 
        .D(\CoreAPB3_0/u_mux_p_to_b3/PRDATA_0_iv_0_a2_3_5_3[1]_net_1 ), 
        .Y(\CoreAPB3_0.u_mux_p_to_b3.PRDATA_0_iv_0_a2_3_5[1] ));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_250  (
        .A(VCC), .B(GND), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[62] ), 
        .IPB(\hello_regs_MSS_0/MSS_ADLIB_INST/F_ARID_HSEL1_net[2] ), 
        .IPC());
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_211  (
        .A(VCC), .B(GND), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[29] ), 
        .IPB(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_AWLOCK_HMASTLOCK0_net[1] ), 
        .IPC());
    INV_BA AFLSDF_INV_18 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_101_net_1 ), .Y(
        AFLSDF_INV_18_net_1));
    CFG3 #( .INIT(8'hF2) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_142  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_8_[4]_net_1 ), .B(N_639), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_142_i ));
    CFG3 #( .INIT(8'h02) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_120  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_6_[6]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_652 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_120_net_1 ));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/mem_2__RNI39LF[1]  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_27_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_161_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_2_rs[1] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_2_[1]_net_1 ));
    RGB \FCCC_0/GL1_INST/U0_RGB1_RGB8  (.An(\FCCC_0/GL1_INST/U0_YNn ), 
        .ENn(GND), .YL(\FCCC_0/GL1_INST/U0_RGB1_RGB8_rgbl_net_1 ), .YR(
        \FCCC_0/GL1_INST/U0_RGB1_RGB8_rgbr_net_1 ));
    INV_BA AFLSDF_INV_73 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_77_net_1 ), .Y(
        AFLSDF_INV_73_net_1));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_212_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_108_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_212_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_212_rs_net_1 ));
    INV_BA AFLSDF_INV_8 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_36_net_1 ), .Y(
        AFLSDF_INV_8_net_1));
    INV_BA AFLSDF_INV_124 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_5_net_1 ), .Y(
        AFLSDF_INV_124_net_1));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_240_rs_RNIH9KU  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_17_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_240_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_12_rs[1] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_12_[1]_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_9_[6]  (.D(
        \CoreAPB3_0_APBmslave5_PWDATA[6] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB16_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_9__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_202_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_9_rs[6] ));
    INV_BA AFLSDF_INV_138 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_7_net_1 ), .Y(
        AFLSDF_INV_138_net_1));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_142_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_68_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_142_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_142_rs_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_43_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB5_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_5__1_sqmuxa ), .ALn(
        AFLSDF_INV_88_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(GND)
        , .Q(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_43_set_net_1 ));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_126  (
        .A(GND), .B(GND), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[1] ), .IPB(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[8] ), .IPC()
        );
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_249  (
        .A(VCC), .B(GND), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[61] ), 
        .IPB(\hello_regs_MSS_0/MSS_ADLIB_INST/F_ARID_HSEL1_net[1] ), 
        .IPC());
    CFG4 #( .INIT(16'h0BFF) )  
        \CoreAPB3_0/u_mux_p_to_b3/PRDATA_0_iv_0_1[3]  (.A(
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PADDR[17] ), .B(
        \CoreAPB3_0_APBmslave5_PRDATA[3] ), .C(
        \CoreAPB3_0/u_mux_p_to_b3/PRDATA_0_iv_0_s_0_0[3]_net_1 ), .D(
        N_625), .Y(\CoreAPB3_0/u_mux_p_to_b3/PRDATA_0_iv_0_1[3]_net_1 )
        );
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_114_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB16_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_14__1_sqmuxa ), .ALn(
        AFLSDF_INV_89_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(GND)
        , .Q(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_114_set_net_1 ));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_40  (.A(
        GND), .B(GND), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[23] ), .IPB(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[30] ), .IPC());
    INV_BA AFLSDF_INV_68 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_40_net_1 ), .Y(
        AFLSDF_INV_68_net_1));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_91  (.A(
        VCC), .B(VCC), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/TX_CLKPF_net ), .IPB(
        \hello_regs_MSS_0/MSS_ADLIB_INST/RXDF_net[7] ), .IPC());
    CFG4 #( .INIT(16'hF8F0) )  
        \CoreAPB3_0/u_mux_p_to_b3/PRDATA_0_iv_0[0]  (.A(N_639), .B(
        \GPIO_OUT_1_c[0] ), .C(
        \CoreAPB3_0/u_mux_p_to_b3/PRDATA_0_iv_0_0[0]_net_1 ), .D(
        \CoreAPB3_0.u_mux_p_to_b3.PRDATA_0_iv_0_a2_3_5[1] ), .Y(
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[0] ));
    SLE \COREAPBLSRAM_0/PRDATA_reg[17]  (.D(
        \COREAPBLSRAM_0.lsram_width32_PRDATA[17] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB8_rgbr_net_1 ), .EN(
        \COREAPBLSRAM_0.PRDATA4 ), .ALn(
        \hello_regs_MSS_0/MSS_ADLIB_INST_RNIUO3B/U0_RGB1_RGB0_rgbr_net_1 )
        , .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \COREAPBLSRAM_0.PRDATA_reg[17] ));
    CFG4 #( .INIT(16'h7530) )  
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_3[2]  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_2_[2]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/mem_13_[2]_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/N_646 ), .D(
        \reg_apb_wrp_0/reg16x8_0/N_642 ), .Y(
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_3[2]_net_1 ));
    INV_BA AFLSDF_INV_121 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_48_net_1 ), .Y(
        AFLSDF_INV_121_net_1));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_232_rs_RNIP37Q  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_93_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_232_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_11_rs[5] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_11_[5]_net_1 ));
    IOTRI_OB_EB \GPIO_OUT_1_obuf[2]/U0/U_IOTRI  (.D(\GPIO_OUT_1_c[2] ), 
        .E(VCC), .DOUT(\GPIO_OUT_1_obuf[2]/U0/DOUT1 ), .EOUT(
        \GPIO_OUT_1_obuf[2]/U0/EOUT1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_75_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB16_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_9__1_sqmuxa ), .ALn(
        AFLSDF_INV_90_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(GND)
        , .Q(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_75_set_net_1 ));
    CFG3 #( .INIT(8'hF2) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_220  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_14_[4]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_650 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_220_i ));
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_data_out8_22  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_12_[6]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_644 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_22_net_1 ));
    CFG3 #( .INIT(8'hF2) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_172  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_10_[3]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_647 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_172_i ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_190_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_72_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_190_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_190_rs_net_1 ));
    CFG3 #( .INIT(8'hF2) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_211  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_13_[3]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_646 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_211_i ));
    CFG4 #( .INIT(16'h0800) )  
        \reg_apb_wrp_0/reg16x8_0/WRITE_GEN.mem_11__2_i_a2[5]  (.A(
        \CoreAPB3_0_APBmslave5_PADDR[2] ), .B(
        \CoreAPB3_0_APBmslave5_PADDR[5] ), .C(
        \CoreAPB3_0_APBmslave5_PADDR[4] ), .D(
        \CoreAPB3_0_APBmslave5_PADDR[3] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/N_649 ));
    CFG3 #( .INIT(8'h02) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_100  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_10_[7]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_647 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_100_net_1 ));
    CFG3 #( .INIT(8'hF2) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_195  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_5_[4]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_653 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_195_i ));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_102  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/RCGF_net[2] ), .IPB(
        \hello_regs_MSS_0/MSS_ADLIB_INST/RCGF_net[9] ), .IPC());
    SLE \reg_apb_wrp_0/reg16x8_0/mem_13_[3]  (.D(
        \CoreAPB3_0_APBmslave5_PWDATA[3] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB8_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_13__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_211_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_13_rs[3] ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_168_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_98_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_168_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_168_rs_net_1 ));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_184_rs_RNIOI4M  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_69_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_184_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_8_rs[5] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_8_[5]_net_1 ));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_248  (
        .A(VCC), .B(GND), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[60] ), 
        .IPB(\hello_regs_MSS_0/MSS_ADLIB_INST/F_ARID_HSEL1_net[0] ), 
        .IPC());
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/mem_10__RNISK1P[3]  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_96_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_172_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_10_rs[3] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_10_[3]_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_12_[3]  (.D(
        \CoreAPB3_0_APBmslave5_PWDATA[3] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB13_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_12__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_243_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_12_rs[3] ));
    CFG3 #( .INIT(8'hF2) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_200  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_9_[5]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_643 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_200_i ));
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_data_out8_20  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_12_[4]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_644 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_20_net_1 ));
    INV_BA AFLSDF_INV_116 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_15_net_1 ), .Y(
        AFLSDF_INV_116_net_1));
    CFG3 #( .INIT(8'hF2) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_141  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_4_[5]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_648 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_141_i ));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_254  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[2] ), 
        .IPB(\hello_regs_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[14] )
        , .IPC());
    INV_BA AFLSDF_INV_75 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_126_net_1 ), .Y(
        AFLSDF_INV_75_net_1));
    CFG3 #( .INIT(8'hF2) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_193  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_5_[3]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_653 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_193_i ));
    IOTRI_OB_EB \MSS_RESET_N_M2F_obuf/U0/U_IOTRI  (.D(
        \hello_regs_MSS_0/FPGA_RESET_N ), .E(VCC), .DOUT(
        \MSS_RESET_N_M2F_obuf/U0/DOUT1 ), .EOUT(
        \MSS_RESET_N_M2F_obuf/U0/EOUT1 ));
    IP_INTERFACE \FCCC_0/CCC_INST/IP_INTERFACE_8  (.A(VCC), .B(GND), 
        .C(VCC), .IPA(\FCCC_0/CCC_INST/PWRITE_net ), .IPB(
        \FCCC_0/CCC_INST/NGMUX2_SEL_net ), .IPC(
        \FCCC_0/CCC_INST/PWDATA_net[6] ));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_206  (
        .A(VCC), .B(GND), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[24] ), 
        .IPB(\hello_regs_MSS_0/MSS_ADLIB_INST/F_AWLEN_HBURST0_net[2] ), 
        .IPC());
    SLE \COREAPBLSRAM_0/PRDATA_reg[26]  (.D(
        \COREAPBLSRAM_0.lsram_width32_PRDATA[26] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB10_rgbr_net_1 ), .EN(
        \COREAPBLSRAM_0.PRDATA4 ), .ALn(
        \hello_regs_MSS_0/MSS_ADLIB_INST_RNIUO3B/U0_RGB1_RGB2_rgbr_net_1 )
        , .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \COREAPBLSRAM_0.PRDATA_reg[26] ));
    INV_BA AFLSDF_INV_36 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_57_net_1 ), .Y(
        AFLSDF_INV_36_net_1));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/mem_6__RNIFCUM[3]  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_34_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_169_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_6_rs[3] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_6_[3]_net_1 ));
    IOTRI_OB_EB \hello_regs_MSS_0/MMUART_0_TXD_PAD/U_IOOUT  (.D(VCC), 
        .E(VCC), .DOUT(), .EOUT());
    INV_BA AFLSDF_INV_143 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_28_net_1 ), .Y(
        AFLSDF_INV_143_net_1));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_21  (.A(
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[26] ), .B(GND), .C(
        VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[26] ), .IPB(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_SIZE_net[0] ), .IPC());
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_150_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_86_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_150_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_150_rs_net_1 ));
    INV_BA AFLSDF_INV_13 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_120_net_1 ), .Y(
        AFLSDF_INV_13_net_1));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_183_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_48_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_183_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_183_rs_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_79_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB19_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_9__1_sqmuxa ), .ALn(
        AFLSDF_INV_91_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(GND)
        , .Q(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_79_set_net_1 ));
    CFG3 #( .INIT(8'h02) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_112  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_14_[0]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_650 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_112_net_1 ));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/mem_10__RNIAAIG[6]  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_103_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_178_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_10_rs[6] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_10_[6]_net_1 ));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_114  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/FAB_XDATAIN_net[6] ), .IPB(
        \hello_regs_MSS_0/MSS_ADLIB_INST/FAB_VSTATUS_net[3] ), .IPC());
    IP_INTERFACE \FCCC_0/CCC_INST/IP_INTERFACE_12  (.A(VCC), .B(VCC), 
        .C(VCC), .IPA(\FCCC_0/CCC_INST/NGMUX0_ARST_N_net ), .IPB(), 
        .IPC(\FCCC_0/CCC_INST/PADDR_net[2] ));
    CFG3 #( .INIT(8'h02) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_124  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_7_[0]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_641 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_124_net_1 ));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/mem_3__RNICQ721[7]  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_55_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_135_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_3_rs[7] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_3_[7]_net_1 ));
    CFG3 #( .INIT(8'hF2) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_225  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_7_[3]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_641 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_225_i ));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/mem_7__RNIHHAP[5]  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_54_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_229_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_7_rs[5] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_7_[5]_net_1 ));
    INV_BA AFLSDF_INV_114 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_47_net_1 ), .Y(
        AFLSDF_INV_114_net_1));
    CFG3 #( .INIT(8'hF2) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_171  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_6_[4]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_652 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_171_i ));
    CFG3 #( .INIT(8'h80) )  
        \reg_apb_wrp_0/reg16x8_0/mem_5__1_sqmuxa_0_a2  (.A(
        \reg_apb_wrp_0/reg16x8_0/N_653 ), .B(N_637), .C(N_638), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_5__1_sqmuxa ));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_14_[3]  (.D(
        \CoreAPB3_0_APBmslave5_PWDATA[3] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB16_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_14__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_219_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_14_rs[3] ));
    CFG3 #( .INIT(8'hF2) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_136  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_4_[0]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_648 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_136_i ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_20_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB12_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_12__1_sqmuxa ), .ALn(
        AFLSDF_INV_92_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(GND)
        , .Q(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_20_set_net_1 ));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_49_set_RNI9PCL  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_49_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_132_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_3_rs[4] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_3_[4]_net_1 ));
    CFG3 #( .INIT(8'hF2) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_198  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_9_[4]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_643 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_198_i ));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_133  (
        .A(GND), .B(VCC), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[15] ), .IPB(
        ), .IPC());
    SLE_IP_EN 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/FF_5  
        (.EN(\hello_regs_MSS_0/MSS_ADLIB_INST_RNIUO3B/U0_RGB1_YR ), 
        .IPENn(AFLSDF_INV_93_net_1));
    INV_BA AFLSDF_INV_63 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_86_net_1 ), .Y(
        AFLSDF_INV_63_net_1));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_14_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB9_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_5__1_sqmuxa ), .ALn(
        AFLSDF_INV_94_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(GND)
        , .Q(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_14_set_net_1 ));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_137_rs_RNIHLLB  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_2_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_137_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_4_rs[1] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_4_[1]_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_67_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB13_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_4__1_sqmuxa ), .ALn(
        AFLSDF_INV_95_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(GND)
        , .Q(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_67_set_net_1 ));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_149_rs_RNIFB6T  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_85_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_149_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_0_rs[5] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_0_[5]_net_1 ));
    INV_BA AFLSDF_INV_111 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_69_net_1 ), .Y(
        AFLSDF_INV_111_net_1));
    RGB \hello_regs_MSS_0/MSS_ADLIB_INST_RNIUO3B/U0_RGB1_RGB4  (.An(
        \hello_regs_MSS_0/MSS_ADLIB_INST_RNIUO3B/U0_YNn_GSouth ), .ENn(
        GND), .YL(), .YR(
        \hello_regs_MSS_0/MSS_ADLIB_INST_RNIUO3B/U0_RGB1_RGB4_rgbr_net_1 )
        );
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_242  (
        .A(VCC), .B(GND), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[54] ), 
        .IPB(\hello_regs_MSS_0/MSS_ADLIB_INST/F_WSTRB_net[2] ), .IPC());
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_108  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/FAB_XDATAIN_net[0] ), .IPB(), 
        .IPC());
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_243  (
        .A(VCC), .B(GND), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[55] ), 
        .IPB(\hello_regs_MSS_0/MSS_ADLIB_INST/F_WSTRB_net[3] ), .IPC());
    CFG3 #( .INIT(8'h02) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_104  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_13_[0]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_646 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_104_net_1 ));
    CFG3 #( .INIT(8'hF2) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_205  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_6_[1]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_652 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_205_i ));
    CFG4 #( .INIT(16'hFFFE) )  
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_12[3]  (.A(
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_1[3]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_3[3]_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_2[3]_net_1 ), .D(
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_0[3]_net_1 ), .Y(
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_12[3]_net_1 ));
    SLE \COREAPBLSRAM_0/PRDATA_reg[6]  (.D(
        \COREAPBLSRAM_0.lsram_width32_PRDATA[6] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB10_rgbr_net_1 ), .EN(
        \COREAPBLSRAM_0.PRDATA4 ), .ALn(
        \hello_regs_MSS_0/MSS_ADLIB_INST_RNIUO3B/U0_RGB1_RGB2_rgbr_net_1 )
        , .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \COREAPBLSRAM_0.PRDATA_reg[6] ));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_30  (.A(
        GND), .B(GND), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[6] ), .IPB(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[13] ), .IPC());
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_129_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_123_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_129_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_129_rs_net_1 ));
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_data_out8_83  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_0_[3]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_645 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_83_net_1 ));
    sdf_IOPAD_TRI \GPIO_OUT_1_obuf[0]/U0/U_IOPAD  (.PAD(GPIO_OUT_1[0]), 
        .D(\GPIO_OUT_1_obuf[0]/U0/DOUT ), .E(
        \GPIO_OUT_1_obuf[0]/U0/EOUT ));
    CFG3 #( .INIT(8'hF2) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_155  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_1_[3]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_651 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_155_i ));
    INV_BA AFLSDF_INV_122 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_109_net_1 ), .Y(
        AFLSDF_INV_122_net_1));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_119_set_RNIDQL4  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_119_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_223_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_14_rs[7] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_14_[7]_net_1 ));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/mem_11__RNI1QVM[7]  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_95_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_236_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_11_rs[7] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_11_[7]_net_1 ));
    CFG4 #( .INIT(16'h0010) )  
        \CoreAPB3_0/u_mux_p_to_b3/PRDATA_0_iv_0_a2_3_5_4[1]  (.A(
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PADDR[16] ), .B(
        \CoreAPB3_0_APBmslave5_PADDR[0] ), .C(
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PADDR[17] ), .D(
        \CoreAPB3_0_APBmslave5_PADDR[6] ), .Y(
        \CoreAPB3_0/u_mux_p_to_b3/PRDATA_0_iv_0_a2_3_5_4[1]_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_239_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_64_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_239_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_239_rs_net_1 ));
    INV_BA AFLSDF_INV_15 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_26_net_1 ), .Y(
        AFLSDF_INV_15_net_1));
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_data_out8_32  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_6_[2]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_652 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_32_net_1 ));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_123  (
        .A(VCC), .B(GND), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/FAB_HOSTDISCON_net ), .IPB(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[5] ), .IPC()
        );
    CFG3 #( .INIT(8'h02) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_111  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_13_[7]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_646 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_111_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_199_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_24_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_199_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_199_rs_net_1 ));
    sdf_IOPAD_TRI \GPIO_OUT_1_obuf[7]/U0/U_IOPAD  (.PAD(GPIO_OUT_1[7]), 
        .D(\GPIO_OUT_1_obuf[7]/U0/DOUT ), .E(
        \GPIO_OUT_1_obuf[7]/U0/EOUT ));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_81  (.A(
        VCC), .B(VCC), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[15] ), 
        .IPB(
        \hello_regs_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[22] ), 
        .IPC());
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_61_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB14_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_15__1_sqmuxa ), .ALn(
        AFLSDF_INV_96_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(GND)
        , .Q(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_61_set_net_1 ));
    CFG3 #( .INIT(8'hF2) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_153  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_1_[1]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_651 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_153_i ));
    INV_BA AFLSDF_INV_65 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_56_net_1 ), .Y(
        AFLSDF_INV_65_net_1));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_216_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_112_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_216_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_216_rs_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_182_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_88_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_182_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_182_rs_net_1 ));
    IOOUTFF_BYPASS \GPIO_OUT_1_obuf[0]/U0/U_IOOUTFF  (.A(
        \GPIO_OUT_1_obuf[0]/U0/DOUT1 ), .Y(
        \GPIO_OUT_1_obuf[0]/U0/DOUT ));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_9  (.A(
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[7] ), .B(
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[14] ), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[7] ), .IPB(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[14] ), .IPC());
    CFG4 #( .INIT(16'hEAC0) )  
        \CoreAPB3_0/u_mux_p_to_b3/PRDATA_0_iv_0_0[6]  (.A(
        \COREAPBLSRAM_0.PRDATA_reg[6] ), .B(
        \CoreAPB3_0/u_mux_p_to_b3/PRDATA_0_iv_0_a2_2_0[6]_net_1 ), .C(
        \CoreAPB3_0.u_mux_p_to_b3.PRDATA_0_iv_0_a2_3_5[1] ), .D(
        \CoreAPB3_0/u_mux_p_to_b3/N_636 ), .Y(
        \CoreAPB3_0/u_mux_p_to_b3/PRDATA_0_iv_0_0[6]_net_1 ));
    CFG4 #( .INIT(16'hECA0) )  \CoreAPB3_0/u_mux_p_to_b3/PRDATA_0[29]  
        (.A(\CoreAPB3_0/u_mux_p_to_b3/N_636 ), .B(
        \COREAPBLSRAM_0.PRDATA4 ), .C(\COREAPBLSRAM_0.PRDATA_reg[29] ), 
        .D(\COREAPBLSRAM_0.lsram_width32_PRDATA[29] ), .Y(
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[29] ));
    CFG2_IP_BC 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/CFG_30  
        (.B(\CoreAPB3_0_APBmslave5_PWDATA[15] ), .C(
        \CoreAPB3_0_APBmslave5_PADDR[7] ), .IPB(
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/A_DIN_net[16] )
        , .IPC(
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/A_ADDR_net[12] )
        );
    INV_BA AFLSDF_INV_87 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_99_net_1 ), .Y(
        AFLSDF_INV_87_net_1));
    CFG4 #( .INIT(16'h7350) )  
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_0[0]  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_11_[0]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/mem_10_[0]_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/N_649 ), .D(
        \reg_apb_wrp_0/reg16x8_0/N_647 ), .Y(
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_0[0]_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_241_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_66_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_241_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_241_rs_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_208_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_104_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_208_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_208_rs_net_1 ));
    INV_BA AFLSDF_INV_72 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_82_net_1 ), .Y(
        AFLSDF_INV_72_net_1));
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_data_out8_30  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_6_[1]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_652 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_30_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_224_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_89_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_224_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_224_rs_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_145_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_82_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_145_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_145_rs_net_1 ));
    IOTRI_OB_EB \GPIO_OUT_1_obuf[5]/U0/U_IOTRI  (.D(\GPIO_OUT_1_c[5] ), 
        .E(VCC), .DOUT(\GPIO_OUT_1_obuf[5]/U0/DOUT1 ), .EOUT(
        \GPIO_OUT_1_obuf[5]/U0/EOUT1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_102_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB8_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_10__1_sqmuxa ), .ALn(
        AFLSDF_INV_97_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(GND)
        , .Q(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_102_set_net_1 ));
    IP_INTERFACE \FCCC_0/CCC_INST/IP_INTERFACE_4  (.A(VCC), .B(VCC), 
        .C(VCC), .IPA(), .IPB(\FCCC_0/CCC_INST/NGMUX0_HOLD_N_net ), 
        .IPC(\FCCC_0/CCC_INST/PWDATA_net[2] ));
    INV_BA AFLSDF_INV_128 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_31_net_1 ), .Y(
        AFLSDF_INV_128_net_1));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_96_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB11_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_10__1_sqmuxa ), .ALn(
        AFLSDF_INV_98_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(GND)
        , .Q(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_96_set_net_1 ));
    SLE \COREAPBLSRAM_0/PRDATA_reg[23]  (.D(
        \COREAPBLSRAM_0.lsram_width32_PRDATA[23] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB9_rgbr_net_1 ), .EN(
        \COREAPBLSRAM_0.PRDATA4 ), .ALn(
        \hello_regs_MSS_0/MSS_ADLIB_INST_RNIUO3B/U0_RGB1_RGB1_rgbr_net_1 )
        , .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \COREAPBLSRAM_0.PRDATA_reg[23] ));
    CFG3 #( .INIT(8'hF2) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_129  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_3_[1]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_655 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_129_i ));
    CFG3 #( .INIT(8'hF2) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_158  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_1_[6]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_651 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_158_i ));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_282  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PADDR_net[5] ), 
        .IPB(
        \hello_regs_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[9] ), 
        .IPC());
    IOENFF_BYPASS \GPIO_OUT_1_obuf[4]/U0/U_IOENFF  (.A(
        \GPIO_OUT_1_obuf[4]/U0/EOUT1 ), .Y(
        \GPIO_OUT_1_obuf[4]/U0/EOUT ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_215_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_111_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_215_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_215_rs_net_1 ));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_283  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PADDR_net[6] ), 
        .IPB(
        \hello_regs_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[10] ), 
        .IPC());
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_159_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_46_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_159_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_159_rs_net_1 ));
    IOIN_IB \hello_regs_MSS_0/MMUART_0_RXD_PAD/U_IOIN  (.YIN(
        \hello_regs_MSS_0/MMUART_0_RXD_PAD/YIN ), .E(GND), .Y());
    CFG3 #( .INIT(8'hF2) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_231  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_7_[6]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_641 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_231_i ));
    SLE_IP_EN 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/FF_8  
        (.EN(VCC), .IPENn(AFLSDF_INV_99_net_1));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_23_set_RNIRPRV  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_23_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_247_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_12_rs[7] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_12_[7]_net_1 ));
    INV_BA AFLSDF_INV_130 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_16_net_1 ), .Y(
        AFLSDF_INV_130_net_1));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_2_[1]  (.D(
        \CoreAPB3_0_APBmslave5_PWDATA[1] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB0_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_2__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_161_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_2_rs[1] ));
    CFG4 #( .INIT(16'hFFFE) )  
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_13[2]  (.A(
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_4[2]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_5[2]_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_7[2]_net_1 ), .D(
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_6[2]_net_1 ), .Y(
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_13[2]_net_1 ));
    CFG4 #( .INIT(16'h7530) )  
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_6[4]  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_4_[4]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/mem_1_[4]_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/N_651 ), .D(
        \reg_apb_wrp_0/reg16x8_0/N_648 ), .Y(
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_6[4]_net_1 ));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_82_set_RNI5G7C  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_82_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_145_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_0_rs[2] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_0_[2]_net_1 ));
    CFG4 #( .INIT(16'h0004) )  
        \reg_apb_wrp_0/reg16x8_0/WRITE_GEN.mem_8__2_i_0_0_a2[6]  (.A(
        \CoreAPB3_0_APBmslave5_PADDR[2] ), .B(
        \CoreAPB3_0_APBmslave5_PADDR[5] ), .C(
        \CoreAPB3_0_APBmslave5_PADDR[4] ), .D(
        \CoreAPB3_0_APBmslave5_PADDR[3] ), .Y(N_639));
    INV_BA AFLSDF_INV_112 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_18_net_1 ), .Y(
        AFLSDF_INV_112_net_1));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_33_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB1_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_2__1_sqmuxa ), .ALn(
        AFLSDF_INV_100_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_33_set_net_1 ));
    CFG4 #( .INIT(16'hECA0) )  \CoreAPB3_0/u_mux_p_to_b3/PRDATA_0[12]  
        (.A(\CoreAPB3_0/u_mux_p_to_b3/N_636 ), .B(
        \COREAPBLSRAM_0.PRDATA4 ), .C(\COREAPBLSRAM_0.PRDATA_reg[12] ), 
        .D(\COREAPBLSRAM_0.lsram_width32_PRDATA[12] ), .Y(
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[12] ));
    INV_BA AFLSDF_INV_2 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_112_net_1 ), .Y(
        AFLSDF_INV_2_net_1));
    CFG2 #( .INIT(4'h1) )  \reg_apb_wrp_0/reg16x8_0/data_out_RNO[4]  (
        .A(\reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_13[4]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_12[4]_net_1 ), .Y(
        \reg_apb_wrp_0/reg16x8_0/N_41_i_0 ));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_2  (.A(
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[0] ), .B(VCC), .C(
        VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[0] ), .IPB(), 
        .IPC());
    INV_BA AFLSDF_INV_89 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_114_net_1 ), .Y(
        AFLSDF_INV_89_net_1));
    CFG3 #( .INIT(8'h02) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_109  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_13_[5]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_646 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_109_net_1 ));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_176_rs_RNI6V5A  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_102_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_176_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_10_rs[5] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_10_[5]_net_1 ));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_139  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/SMBSUS_NI1_net ), .IPB(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F2_DMAREADY_net[1] ), .IPC());
    CFG3 #( .INIT(8'hF2) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_254  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_15_[7]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_654 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_254_i ));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_261  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[9] ), 
        .IPB(\hello_regs_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[21] )
        , .IPC());
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_13  (.A(
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[18] ), .B(VCC), .C(
        VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[18] ), .IPB(), 
        .IPC());
    CFG3 #( .INIT(8'hF2) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_187  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_5_[0]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_653 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_187_i ));
    RGB \FCCC_0/GL1_INST/U0_RGB1_RGB4  (.An(\FCCC_0/GL1_INST/U0_YNn ), 
        .ENn(GND), .YL(), .YR(
        \FCCC_0/GL1_INST/U0_RGB1_RGB4_rgbr_net_1 ));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_240  (
        .A(VCC), .B(GND), .C(GND), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[52] ), 
        .IPB(\hello_regs_MSS_0/MSS_ADLIB_INST/F_WSTRB_net[0] ), .IPC(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WVALID_net ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_68_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB7_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_8__1_sqmuxa ), .ALn(
        AFLSDF_INV_101_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_68_set_net_1 ));
    CFG4 #( .INIT(16'hECA0) )  \CoreAPB3_0/u_mux_p_to_b3/PRDATA_0[20]  
        (.A(\CoreAPB3_0/u_mux_p_to_b3/N_636 ), .B(
        \COREAPBLSRAM_0.PRDATA4 ), .C(\COREAPBLSRAM_0.PRDATA_reg[20] ), 
        .D(\COREAPBLSRAM_0.lsram_width32_PRDATA[20] ), .Y(
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[20] ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_254_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_60_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_254_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_254_rs_net_1 ));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_96  (.A(
        VCC), .B(VCC), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/CRSF_net ), .IPB(), .IPC());
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_data_out8_74  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_9_[2]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_643 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_74_net_1 ));
    CFG3 #( .INIT(8'hF2) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_132  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_3_[4]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_655 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_132_i ));
    INV_BA AFLSDF_INV_12 (.A(AFLSDF_INV_12_net_1), .Y(
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/B_DOUT_CLK_net )
        );
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_17_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB18_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_12__1_sqmuxa ), .ALn(
        AFLSDF_INV_102_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_17_set_net_1 ));
    CFG4 #( .INIT(16'hFFFE) )  
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_13[1]  (.A(
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_4[1]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_5[1]_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_7[1]_net_1 ), .D(
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_6[1]_net_1 ), .Y(
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_13[1]_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_44_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB14_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_1__1_sqmuxa ), .ALn(
        AFLSDF_INV_103_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_44_set_net_1 ));
    INV_BA AFLSDF_INV_71 (.A(AFLSDF_INV_71_net_1), .Y(
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/A_DOUT_ARST_N_net )
        );
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_232_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_93_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_232_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_232_rs_net_1 ));
    CFG4 #( .INIT(16'hF8F0) )  
        \CoreAPB3_0/u_mux_p_to_b3/PRDATA_0_iv_0[4]  (.A(N_639), .B(
        \GPIO_OUT_1_c[4] ), .C(
        \CoreAPB3_0/u_mux_p_to_b3/PRDATA_0_iv_0_1[4]_net_1 ), .D(
        \CoreAPB3_0.u_mux_p_to_b3.PRDATA_0_iv_0_a2_3_5[1] ), .Y(
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[4] ));
    CFG4 #( .INIT(16'hFFB3) )  
        \CoreAPB3_0/u_mux_p_to_b3/PRDATA_0_iv_0[2]  (.A(
        \COREAPBLSRAM_0.lsram_width32_PRDATA[2] ), .B(
        \CoreAPB3_0/u_mux_p_to_b3/PRDATA_0_iv_0_1_0[2]_net_1 ), .C(
        \COREAPBLSRAM_0.PRDATA4 ), .D(
        \CoreAPB3_0/u_mux_p_to_b3/PRDATA_0_iv_0_0[2]_net_1 ), .Y(
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[2] ));
    IP_INTERFACE \FCCC_0/CCC_INST/IP_INTERFACE_1  (.A(VCC), .B(VCC), 
        .C(VCC), .IPA(\FCCC_0/CCC_INST/CLK1_net ), .IPB(
        \FCCC_0/CCC_INST/PENABLE_net ), .IPC());
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_171  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/MMUART1_DCD_F2H_SCP_net ), 
        .IPB(\hello_regs_MSS_0/MSS_ADLIB_INST/MGPIO17B_F2H_GPIN_net ), 
        .IPC());
    INV_BA AFLSDF_INV_118 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_41_net_1 ), .Y(
        AFLSDF_INV_118_net_1));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_110  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/FAB_XDATAIN_net[2] ), .IPB(), 
        .IPC());
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_75_set_RNINJ8Q  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_75_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_196_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_9_rs[3] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_9_[3]_net_1 ));
    CFG4 #( .INIT(16'h7350) )  
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_1[4]  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_15_[4]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/mem_14_[4]_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/N_654 ), .D(
        \reg_apb_wrp_0/reg16x8_0/N_650 ), .Y(
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_1[4]_net_1 ));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_129  (
        .A(GND), .B(GND), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[4] ), .IPB(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[11] ), .IPC(
        ));
    INV_BA AFLSDF_INV_105 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_65_net_1 ), .Y(
        AFLSDF_INV_105_net_1));
    INV_BA AFLSDF_INV_62 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_3_net_1 ), .Y(
        AFLSDF_INV_62_net_1));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_76_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB14_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_9__1_sqmuxa ), .ALn(
        AFLSDF_INV_104_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_76_set_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_13_[7]  (.D(
        \CoreAPB3_0_APBmslave5_PWDATA[7] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB8_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_13__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_215_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_13_rs[7] ));
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_data_out8_77  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_9_[5]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_643 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_77_net_1 ));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_12  (.A(
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[17] ), .B(VCC), .C(
        VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[17] ), .IPB(), 
        .IPC());
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_150_rs_RNI9PMB  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_86_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_150_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_0_rs[6] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_0_[6]_net_1 ));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_215  (
        .A(GND), .B(GND), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_AWSIZE_HSIZE0_net[1] ), 
        .IPB(\hello_regs_MSS_0/MSS_ADLIB_INST/F_WID_HREADY01_net[3] ), 
        .IPC());
    INV_BA AFLSDF_INV_147 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_25_net_1 ), .Y(
        AFLSDF_INV_147_net_1));
    SLE \COREAPBLSRAM_0/PRDATA_reg[16]  (.D(
        \COREAPBLSRAM_0.lsram_width32_PRDATA[16] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB8_rgbr_net_1 ), .EN(
        \COREAPBLSRAM_0.PRDATA4 ), .ALn(
        \hello_regs_MSS_0/MSS_ADLIB_INST_RNIUO3B/U0_RGB1_RGB0_rgbr_net_1 )
        , .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \COREAPBLSRAM_0.PRDATA_reg[16] ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_65_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB13_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_4__1_sqmuxa ), .ALn(
        AFLSDF_INV_105_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_65_set_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_12_[7]  (.D(
        \CoreAPB3_0_APBmslave5_PWDATA[7] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB17_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_12__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_247_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_12_rs[7] ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_105_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB9_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_13__1_sqmuxa ), .ALn(
        AFLSDF_INV_106_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_105_set_net_1 )
        );
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_255_rs_RNISCAF  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_61_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_255_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_15_rs[4] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_15_[4]_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_107_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB7_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_13__1_sqmuxa ), .ALn(
        AFLSDF_INV_107_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_107_set_net_1 )
        );
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_8  (.A(
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[6] ), .B(
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[13] ), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[6] ), .IPB(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[13] ), .IPC());
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_26  (.A(
        GND), .B(VCC), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[2] ), .IPB(), 
        .IPC());
    CFG4 #( .INIT(16'h7350) )  
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_1[0]  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_15_[0]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/mem_14_[0]_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/N_654 ), .D(
        \reg_apb_wrp_0/reg16x8_0/N_650 ), .Y(
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_1[0]_net_1 ));
    CFG4 #( .INIT(16'hEAC0) )  
        \CoreAPB3_0/u_mux_p_to_b3/PRDATA_0_iv_0_0[2]  (.A(
        \COREAPBLSRAM_0.PRDATA_reg[2] ), .B(
        \CoreAPB3_0/u_mux_p_to_b3/PRDATA_0_iv_0_a2_2_0[2]_net_1 ), .C(
        \CoreAPB3_0.u_mux_p_to_b3.PRDATA_0_iv_0_a2_3_5[1] ), .D(
        \CoreAPB3_0/u_mux_p_to_b3/N_636 ), .Y(
        \CoreAPB3_0/u_mux_p_to_b3/PRDATA_0_iv_0_0[2]_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_11_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB17_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_1__1_sqmuxa ), .ALn(
        AFLSDF_INV_108_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_11_set_net_1 ));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_115  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/FAB_XDATAIN_net[7] ), .IPB(
        \hello_regs_MSS_0/MSS_ADLIB_INST/FAB_VSTATUS_net[4] ), .IPC());
    INV_BA AFLSDF_INV_48 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_73_net_1 ), .Y(
        AFLSDF_INV_48_net_1));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/mem_11__RNIQ77K[3]  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_91_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_228_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_11_rs[3] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_11_[3]_net_1 ));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_244  (
        .A(VCC), .B(GND), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[56] ), 
        .IPB(\hello_regs_MSS_0/MSS_ADLIB_INST/F_WSTRB_net[4] ), .IPC());
    IP_INTERFACE \FCCC_0/CCC_INST/IP_INTERFACE_15  (.A(VCC), .B(VCC), 
        .C(VCC), .IPA(\FCCC_0/CCC_INST/NGMUX3_ARST_N_net ), .IPB(
        \FCCC_0/CCC_INST/GPD1_ARST_N_net ), .IPC(
        \FCCC_0/CCC_INST/PADDR_net[5] ));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_164  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/MGPIO13A_F2H_GPIN_net ), .IPB(
        \hello_regs_MSS_0/MSS_ADLIB_INST/MGPIO16A_F2H_GPIN_net ), .IPC(
        ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_128_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_121_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_128_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_128_rs_net_1 ));
    CFG2 #( .INIT(4'h1) )  \reg_apb_wrp_0/reg16x8_0/data_out_RNO[2]  (
        .A(\reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_13[2]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_12[2]_net_1 ), .Y(
        \reg_apb_wrp_0/reg16x8_0/N_15_i_0 ));
    CFG3 #( .INIT(8'hF2) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_131  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_3_[3]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_655 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_131_i ));
    CFG4 #( .INIT(16'h7350) )  
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_2[2]  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_12_[2]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/mem_9_[2]_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/N_644 ), .D(
        \reg_apb_wrp_0/reg16x8_0/N_643 ), .Y(
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_2[2]_net_1 ));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_117  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/FAB_RXACTIVE_net ), .IPB(
        \hello_regs_MSS_0/MSS_ADLIB_INST/FAB_VSTATUS_net[6] ), .IPC());
    sdf_IOPAD_TRI \GPIO_OUT_1_obuf[4]/U0/U_IOPAD  (.PAD(GPIO_OUT_1[4]), 
        .D(\GPIO_OUT_1_obuf[4]/U0/DOUT ), .E(
        \GPIO_OUT_1_obuf[4]/U0/EOUT ));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_71  (.A(
        VCC), .B(VCC), .C(VCC), .IPA(), .IPB(
        \hello_regs_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[5] ), 
        .IPC());
    INV_BA AFLSDF_INV_30 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_90_net_1 ), .Y(
        AFLSDF_INV_30_net_1));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_280  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PADDR_net[3] ), 
        .IPB(
        \hello_regs_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[7] ), 
        .IPC());
    CFG3 #( .INIT(8'hF2) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_242  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_12_[2]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_644 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_242_i ));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_15_[4]  (.D(
        \CoreAPB3_0_APBmslave5_PWDATA[4] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB14_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_15__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_255_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_15_rs[4] ));
    SLE \reg_apb_wrp_0/reg16x8_0/data_out[1]  (.D(
        \reg_apb_wrp_0/reg16x8_0/N_13_i_0 ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB11_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/rd_enable ), .ALn(
        \hello_regs_MSS_0/MSS_ADLIB_INST_RNIUO3B/U0_RGB1_RGB3_rgbr_net_1 )
        , .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreAPB3_0_APBmslave5_PRDATA[1] ));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_251  (
        .A(VCC), .B(GND), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[63] ), 
        .IPB(\hello_regs_MSS_0/MSS_ADLIB_INST/F_ARID_HSEL1_net[3] ), 
        .IPC());
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_185_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_10_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_185_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_185_rs_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_14_[7]  (.D(
        \CoreAPB3_0_APBmslave5_PWDATA[7] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB15_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_14__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_223_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_14_rs[7] ));
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_data_out8_71  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_8_[7]_net_1 ), .B(N_639), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_71_net_1 ));
    INV_BA AFLSDF_INV_11 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_117_net_1 ), .Y(
        AFLSDF_INV_11_net_1));
    INV_BA AFLSDF_INV_0 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_80_net_1 ), .Y(
        AFLSDF_INV_0_net_1));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_170_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_99_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_170_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_170_rs_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_92_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB5_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_11__1_sqmuxa ), .ALn(
        AFLSDF_INV_109_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_92_set_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_23_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB17_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_12__1_sqmuxa ), .ALn(
        AFLSDF_INV_110_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_23_set_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_198_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_76_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_198_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_198_rs_net_1 ));
    SLE \COREAPBLSRAM_0/PRDATA_reg[3]  (.D(
        \COREAPBLSRAM_0.lsram_width32_PRDATA[3] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB10_rgbr_net_1 ), .EN(
        \COREAPBLSRAM_0.PRDATA4 ), .ALn(
        \hello_regs_MSS_0/MSS_ADLIB_INST_RNIUO3B/U0_RGB1_RGB2_rgbr_net_1 )
        , .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \COREAPBLSRAM_0.PRDATA_reg[3] ));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_13_[2]  (.D(
        \CoreAPB3_0_APBmslave5_PWDATA[2] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB4_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_13__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_210_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_13_rs[2] ));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_60_set_RNIT81Q  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_60_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_254_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_15_rs[7] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_15_[7]_net_1 ));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_41  (.A(
        GND), .B(GND), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[24] ), .IPB(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[31] ), .IPC());
    INV_BA AFLSDF_INV_84 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_30_net_1 ), .Y(
        AFLSDF_INV_84_net_1));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_69_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB7_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_8__1_sqmuxa ), .ALn(
        AFLSDF_INV_111_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_69_set_net_1 ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[4].APB_8.GPOUT_reg[4]  (.D(
        \CoreAPB3_0_APBmslave5_PWDATA[4] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB8_rgbr_net_1 ), .EN(
        \CoreGPIO_0/GPOUT_reg35 ), .ALn(
        \hello_regs_MSS_0/MSS_ADLIB_INST_RNIUO3B/U0_RGB1_RGB0_rgbr_net_1 )
        , .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \GPIO_OUT_1_c[4] ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[1].APB_8.GPOUT_reg[1]  (.D(
        \CoreAPB3_0_APBmslave5_PWDATA[1] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB12_rgbr_net_1 ), .EN(
        \CoreGPIO_0/GPOUT_reg35 ), .ALn(
        \hello_regs_MSS_0/MSS_ADLIB_INST_RNIUO3B/U0_RGB1_RGB4_rgbr_net_1 )
        , .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \GPIO_OUT_1_c[1] ));
    INV_BA AFLSDF_INV_61 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_111_net_1 ), .Y(
        AFLSDF_INV_61_net_1));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_12_[2]  (.D(
        \CoreAPB3_0_APBmslave5_PWDATA[2] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB17_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_12__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_242_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_12_rs[2] ));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_0_[3]  (.D(
        \CoreAPB3_0_APBmslave5_PWDATA[3] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB15_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_0__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_146_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_0_rs[3] ));
    CFG4 #( .INIT(16'h0010) )  
        \reg_apb_wrp_0/reg16x8_0/WRITE_GEN.mem_4__2_i_a2[3]  (.A(
        \CoreAPB3_0_APBmslave5_PADDR[2] ), .B(
        \CoreAPB3_0_APBmslave5_PADDR[5] ), .C(
        \CoreAPB3_0_APBmslave5_PADDR[4] ), .D(
        \CoreAPB3_0_APBmslave5_PADDR[3] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/N_648 ));
    CFG3 #( .INIT(8'hF2) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_197  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_5_[5]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_653 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_197_i ));
    CFG3 #( .INIT(8'hF2) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_166  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_2_[6]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_642 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_166_i ));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_112  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/FAB_XDATAIN_net[4] ), .IPB(
        \hello_regs_MSS_0/MSS_ADLIB_INST/FAB_VSTATUS_net[1] ), .IPC());
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/mem_14__RNI7A3Q[5]  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_117_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_221_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_14_rs[5] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_14_[5]_net_1 ));
    CFG4 #( .INIT(16'hFFB3) )  
        \CoreAPB3_0/u_mux_p_to_b3/PRDATA_0_iv_0[6]  (.A(
        \COREAPBLSRAM_0.lsram_width32_PRDATA[6] ), .B(
        \CoreAPB3_0/u_mux_p_to_b3/PRDATA_0_iv_0_1_0[6]_net_1 ), .C(
        \COREAPBLSRAM_0.PRDATA4 ), .D(
        \CoreAPB3_0/u_mux_p_to_b3/PRDATA_0_iv_0_0[6]_net_1 ), .Y(
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[6] ));
    CFG4 #( .INIT(16'h0100) )  
        \reg_apb_wrp_0/reg16x8_0/WRITE_GEN.mem_2__2_i_a2[3]  (.A(
        \CoreAPB3_0_APBmslave5_PADDR[2] ), .B(
        \CoreAPB3_0_APBmslave5_PADDR[5] ), .C(
        \CoreAPB3_0_APBmslave5_PADDR[4] ), .D(
        \CoreAPB3_0_APBmslave5_PADDR[3] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/N_642 ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_146_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_83_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_146_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_146_rs_net_1 ));
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_data_out8_62  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_15_[5]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_654 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_62_net_1 ));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_239  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[37] ), 
        .IPB(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[49] ), 
        .IPC());
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_177_rs_RNI0RJG  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_122_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_177_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_6_rs[7] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_6_[7]_net_1 ));
    INV_BA AFLSDF_INV_120 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_66_net_1 ), .Y(
        AFLSDF_INV_120_net_1));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_207_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_32_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_207_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_207_rs_net_1 ));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_195_rs_RNIIQQ11  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_47_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_195_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_5_rs[4] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_5_[4]_net_1 ));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_86  (.A(
        VCC), .B(VCC), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[27] ), 
        .IPB(\hello_regs_MSS_0/MSS_ADLIB_INST/RXDF_net[2] ), .IPC());
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_158_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_44_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_158_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_158_rs_net_1 ));
    INV_BA AFLSDF_INV_43 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_6_net_1 ), .Y(
        AFLSDF_INV_43_net_1));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_284  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PADDR_net[7] ), 
        .IPB(
        \hello_regs_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[11] ), 
        .IPC());
    INV_BA AFLSDF_INV_27 (.A(AFLSDF_INV_27_net_1), .Y(
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/B_DOUT_ARST_N_net )
        );
    SLE \reg_apb_wrp_0/reg16x8_0/mem_5_[6]  (.D(
        \CoreAPB3_0_APBmslave5_PWDATA[6] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB5_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_5__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_199_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_5_rs[6] ));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/mem_2__RNI2U0J[3]  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_31_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_163_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_2_rs[3] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_2_[3]_net_1 ));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_60  (.A(
        GND), .B(VCC), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[21] ), .IPB(), 
        .IPC());
    RGB \FCCC_0/GL1_INST/U0_RGB1_RGB18  (.An(
        \FCCC_0/GL1_INST/U0_YNn_GSouth ), .ENn(GND), .YL(
        \FCCC_0/GL1_INST/U0_RGB1_RGB18_rgbl_net_1 ), .YR(
        \FCCC_0/GL1_INST/U0_RGB1_RGB18_rgbr_net_1 ));
    CFG2_IP_BC 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/CFG_15  
        (.B(\CoreAPB3_0_APBmslave5_PWDATA[27] ), .C(
        \CoreAPB3_0_APBmslave5_PADDR[1] ), .IPB(
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/B_DIN_net[12] )
        , .IPC(
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/B_ADDR_net[6] )
        );
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_data_out8_98  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_10_[1]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_647 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_98_net_1 ));
    RGB \FCCC_0/GL1_INST/U0_RGB1_RGB1  (.An(\FCCC_0/GL1_INST/U0_YNn ), 
        .ENn(GND), .YL(), .YR(
        \FCCC_0/GL1_INST/U0_RGB1_RGB1_rgbr_net_1 ));
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_data_out8_86  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_0_[6]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_645 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_86_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_14_[2]  (.D(
        \CoreAPB3_0_APBmslave5_PWDATA[2] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB15_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_14__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_218_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_14_rs[2] ));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_0_[4]  (.D(
        \CoreAPB3_0_APBmslave5_PWDATA[4] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB14_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_0__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_148_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_0_rs[4] ));
    RGB \hello_regs_MSS_0/MSS_ADLIB_INST_RNIUO3B/U0_RGB1_RGB6  (.An(
        \hello_regs_MSS_0/MSS_ADLIB_INST_RNIUO3B/U0_YNn_GSouth ), .ENn(
        GND), .YL(), .YR(
        \hello_regs_MSS_0/MSS_ADLIB_INST_RNIUO3B/U0_RGB1_RGB6_rgbr_net_1 )
        );
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_216  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[0] ), 
        .IPB(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[12] ), 
        .IPC(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[24] ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_18_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB17_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_12__1_sqmuxa ), .ALn(
        AFLSDF_INV_112_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_18_set_net_1 ));
    RGB \FCCC_0/GL1_INST/U0_RGB1_RGB10  (.An(\FCCC_0/GL1_INST/U0_YNn ), 
        .ENn(GND), .YL(\FCCC_0/GL1_INST/U0_RGB1_RGB10_rgbl_net_1 ), 
        .YR(\FCCC_0/GL1_INST/U0_RGB1_RGB10_rgbr_net_1 ));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_25  (.A(
        GND), .B(VCC), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[1] ), .IPB(), 
        .IPC());
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_238  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[36] ), 
        .IPB(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[48] ), 
        .IPC());
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_data_out8_60  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_15_[7]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_654 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_60_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_243_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_19_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_243_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_243_rs_net_1 ));
    CFG3 #( .INIT(8'hF2) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_212  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_13_[4]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_646 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_212_i ));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_3_[3]  (.D(
        \CoreAPB3_0_APBmslave5_PWDATA[3] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB16_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_3__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_131_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_3_rs[3] ));
    SLE \COREAPBLSRAM_0/PRDATA_reg[13]  (.D(
        \COREAPBLSRAM_0.lsram_width32_PRDATA[13] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB8_rgbr_net_1 ), .EN(
        \COREAPBLSRAM_0.PRDATA4 ), .ALn(
        \hello_regs_MSS_0/MSS_ADLIB_INST_RNIUO3B/U0_RGB1_RGB0_rgbr_net_1 )
        , .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \COREAPBLSRAM_0.PRDATA_reg[13] ));
    CFG2 #( .INIT(4'h7) )  
        \CoreAPB3_0/u_mux_p_to_b3/PRDATA_0_iv_0_1_0[7]  (.A(N_637), .B(
        \CoreAPB3_0_APBmslave5_PRDATA[7] ), .Y(
        \CoreAPB3_0/u_mux_p_to_b3/PRDATA_0_iv_0_1_0[7]_net_1 ));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/mem_2__RNI6AGC[4]  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_33_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_164_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_2_rs[4] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_2_[4]_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_100_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB11_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_10__1_sqmuxa ), .ALn(
        AFLSDF_INV_113_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_100_set_net_1 )
        );
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_154  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(), .IPB(
        \hello_regs_MSS_0/MSS_ADLIB_INST/SPI0_SS0_F2H_SCP_net ), .IPC()
        );
    RGB \FCCC_0/GL1_INST/U0_RGB1_RGB5  (.An(\FCCC_0/GL1_INST/U0_YNn ), 
        .ENn(GND), .YL(\FCCC_0/GL1_INST/U0_RGB1_RGB5_rgbl_net_1 ), .YR(
        \FCCC_0/GL1_INST/U0_RGB1_RGB5_rgbr_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_47_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB8_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_5__1_sqmuxa ), .ALn(
        AFLSDF_INV_114_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_47_set_net_1 ));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_229  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[27] ), 
        .IPB(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[39] ), 
        .IPC(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[51] ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_236_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_95_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_236_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_236_rs_net_1 ));
    IOTRI_OB_EB \GPIO_OUT_1_obuf[7]/U0/U_IOTRI  (.D(\GPIO_OUT_1_c[7] ), 
        .E(VCC), .DOUT(\GPIO_OUT_1_obuf[7]/U0/DOUT1 ), .EOUT(
        \GPIO_OUT_1_obuf[7]/U0/EOUT1 ));
    CFG2_IP_BC 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/CFG_25  
        (.B(\CoreAPB3_0_APBmslave5_PWDATA[22] ), .C(
        \CoreAPB3_0_APBmslave5_PADDR[4] ), .IPB(
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/B_DIN_net[6] )
        , .IPC(
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/B_ADDR_net[9] )
        );
    SLE \reg_apb_wrp_0/reg16x8_0/data_out[6]  (.D(
        \reg_apb_wrp_0/reg16x8_0/N_22_i_0 ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB10_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/rd_enable ), .ALn(
        \hello_regs_MSS_0/MSS_ADLIB_INST_RNIUO3B/U0_RGB1_RGB2_rgbr_net_1 )
        , .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreAPB3_0_APBmslave5_PRDATA[6] ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_72_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB19_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_9__1_sqmuxa ), .ALn(
        AFLSDF_INV_115_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_72_set_net_1 ));
    CFG4 #( .INIT(16'hFFFE) )  
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_13[3]  (.A(
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_4[3]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_5[3]_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_7[3]_net_1 ), .D(
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_6[3]_net_1 ), .Y(
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_13[3]_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_141_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_67_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_141_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_141_rs_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_7_[3]  (.D(
        \CoreAPB3_0_APBmslave5_PWDATA[3] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB15_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_7__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_225_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_7_rs[3] ));
    CFG4 #( .INIT(16'hFFFE) )  
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_13[4]  (.A(
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_4[4]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_5[4]_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_7[4]_net_1 ), .D(
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_6[4]_net_1 ), .Y(
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_13[4]_net_1 ));
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_data_out8_44  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_1_[6]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_651 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_44_net_1 ));
    INV_BA AFLSDF_INV_29 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_54_net_1 ), .Y(
        AFLSDF_INV_29_net_1));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_0_[0]  (.D(
        \CoreAPB3_0_APBmslave5_PWDATA[0] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB13_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_0__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_147_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_0_rs[0] ));
    IP_INTERFACE \FCCC_0/CCC_INST/IP_INTERFACE_6  (.A(VCC), .B(VCC), 
        .C(VCC), .IPA(\FCCC_0/CCC_INST/CLK2_net ), .IPB(), .IPC(
        \FCCC_0/CCC_INST/PWDATA_net[4] ));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_118  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(), .IPB(
        \hello_regs_MSS_0/MSS_ADLIB_INST/FAB_VSTATUS_net[7] ), .IPC());
    CFG3 #( .INIT(8'hF2) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_248  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_15_[1]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_654 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_248_i ));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_3_[4]  (.D(
        \CoreAPB3_0_APBmslave5_PWDATA[4] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB13_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_3__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_132_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_3_rs[4] ));
    CFG3 #( .INIT(8'hF2) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_247  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_12_[7]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_644 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_247_i ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_15_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB17_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_1__1_sqmuxa ), .ALn(
        AFLSDF_INV_116_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_15_set_net_1 ));
    INV_BA AFLSDF_INV_45 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_4_net_1 ), .Y(
        AFLSDF_INV_45_net_1));
    CFG3 #( .INIT(8'h10) )  
        \CoreAPB3_0/u_mux_p_to_b3/PRDATA_0_iv_0_a2_3_5_3[1]  (.A(
        \CoreAPB3_0_APBmslave5_PADDR[1] ), .B(
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PADDR[19] ), .C(
        \CoreAPB3_0_APBmslave5_PADDR[7] ), .Y(
        \CoreAPB3_0/u_mux_p_to_b3/PRDATA_0_iv_0_a2_3_5_3[1]_net_1 ));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_31  (.A(
        GND), .B(GND), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[7] ), .IPB(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[14] ), .IPC());
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[0].APB_8.GPOUT_reg[0]  (.D(
        \CoreAPB3_0_APBmslave5_PWDATA[0] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB8_rgbr_net_1 ), .EN(
        \CoreGPIO_0/GPOUT_reg35 ), .ALn(
        \hello_regs_MSS_0/MSS_ADLIB_INST_RNIUO3B/U0_RGB1_RGB0_rgbr_net_1 )
        , .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \GPIO_OUT_1_c[0] ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_235_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_7_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_235_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_235_rs_net_1 ));
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_data_out8_18  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_12_[2]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_644 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_18_net_1 ));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_228  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[26] ), 
        .IPB(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[38] ), 
        .IPC(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[50] ));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_48_set_RNIGQ08  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_48_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_183_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_7_rs[2] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_7_[2]_net_1 ));
    CFG2 #( .INIT(4'h4) )  \COREAPBLSRAM_0/PREADY_reg6_0_a2_0  (.A(
        CoreAPB3_0_APBmslave5_PWRITE), .B(CoreAPB3_0_APBmslave7_PREADY)
        , .Y(\COREAPBLSRAM_0/PREADY_reg6_0_a2_0_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_179_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_124_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_179_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_179_rs_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_8_[3]  (.D(
        \CoreAPB3_0_APBmslave5_PWDATA[3] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB8_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_8__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_241_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_8_rs[3] ));
    CFG3 #( .INIT(8'hF2) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_157  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_1_[5]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_651 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_157_i ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_34_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB17_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_6__1_sqmuxa ), .ALn(
        AFLSDF_INV_117_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_34_set_net_1 ));
    INV_BA AFLSDF_INV_110 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_23_net_1 ), .Y(
        AFLSDF_INV_110_net_1));
    IOENFF_BYPASS \GPIO_OUT_1_obuf[7]/U0/U_IOENFF  (.A(
        \GPIO_OUT_1_obuf[7]/U0/EOUT1 ), .Y(
        \GPIO_OUT_1_obuf[7]/U0/EOUT ));
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_data_out8_47  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_5_[4]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_653 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_47_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_41_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB8_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_5__1_sqmuxa ), .ALn(
        AFLSDF_INV_118_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_41_set_net_1 ));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_7  (.A(
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[5] ), .B(
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[12] ), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[5] ), .IPB(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[12] ), .IPC());
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_143_rs_RNIPAKK  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_8_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_143_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_4_rs[6] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_4_[6]_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_7_[4]  (.D(
        \CoreAPB3_0_APBmslave5_PWDATA[4] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB15_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_7__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_227_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_7_rs[4] ));
    CFG4 #( .INIT(16'hCA00) )  
        \CoreAPB3_0/u_mux_p_to_b3/PRDATA_0_iv_0_s_0_0[3]  (.A(
        \COREAPBLSRAM_0.lsram_width32_PRDATA[3] ), .B(
        \COREAPBLSRAM_0.PRDATA_reg[3] ), .C(N_354), .D(
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PADDR[17] ), .Y(
        \CoreAPB3_0/u_mux_p_to_b3/PRDATA_0_iv_0_s_0_0[3]_net_1 ));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_232  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[30] ), 
        .IPB(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[42] ), 
        .IPC());
    SLE \reg_apb_wrp_0/reg16x8_0/mem_13_[1]  (.D(
        \CoreAPB3_0_APBmslave5_PWDATA[1] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB9_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_13__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_209_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_13_rs[1] ));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_233  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[31] ), 
        .IPB(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[43] ), 
        .IPC());
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_100_set_RNI1BDF  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_100_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_180_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_10_rs[7] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_10_[7]_net_1 ));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_85  (.A(
        VCC), .B(VCC), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[26] ), 
        .IPB(\hello_regs_MSS_0/MSS_ADLIB_INST/RXDF_net[1] ), .IPC());
    IOTRI_OB_EB \GPIO_OUT_1_obuf[1]/U0/U_IOTRI  (.D(\GPIO_OUT_1_c[1] ), 
        .E(VCC), .DOUT(\GPIO_OUT_1_obuf[1]/U0/DOUT1 ), .EOUT(
        \GPIO_OUT_1_obuf[1]/U0/EOUT1 ));
    INV_BA AFLSDF_INV_98 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_96_net_1 ), .Y(
        AFLSDF_INV_98_net_1));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_4_[3]  (.D(
        \CoreAPB3_0_APBmslave5_PWDATA[3] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB17_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_4__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_139_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_4_rs[3] ));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_8_[4]  (.D(
        \CoreAPB3_0_APBmslave5_PWDATA[4] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB7_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_8__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_142_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_8_rs[4] ));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_3_[0]  (.D(
        \CoreAPB3_0_APBmslave5_PWDATA[0] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB9_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_3__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_128_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_3_rs[0] ));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_12_[1]  (.D(
        \CoreAPB3_0_APBmslave5_PWDATA[1] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB18_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_12__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_240_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_12_rs[1] ));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_277  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[1] ), 
        .IPB(
        \hello_regs_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[4] ), 
        .IPC());
    SLE \COREAPBLSRAM_0/PRDATA_reg[0]  (.D(
        \COREAPBLSRAM_0.lsram_width32_PRDATA[0] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB9_rgbr_net_1 ), .EN(
        \COREAPBLSRAM_0.PRDATA4 ), .ALn(
        \hello_regs_MSS_0/MSS_ADLIB_INST_RNIUO3B/U0_RGB1_RGB1_rgbr_net_1 )
        , .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \COREAPBLSRAM_0.PRDATA_reg[0] ));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_4  (.A(
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[2] ), .B(
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[9] ), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[2] ), .IPB(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[9] ), .IPC());
    SLE \reg_apb_wrp_0/reg16x8_0/mem_6_[3]  (.D(
        \CoreAPB3_0_APBmslave5_PWDATA[3] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB17_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_6__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_169_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_6_rs[3] ));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_160  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/MGPIO11A_F2H_GPIN_net ), .IPB(
        \hello_regs_MSS_0/MSS_ADLIB_INST/MGPIO14A_F2H_GPIN_net ), .IPC(
        ));
    CFG3 #( .INIT(8'hF2) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_246  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_12_[6]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_644 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_246_i ));
    CFG4 #( .INIT(16'h7530) )  
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_0_3[6]  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_2_[6]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/mem_13_[6]_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/N_646 ), .D(
        \reg_apb_wrp_0/reg16x8_0/N_642 ), .Y(
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_0_3[6]_net_1 ));
    INV_BA AFLSDF_INV_139 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_35_net_1 ), .Y(
        AFLSDF_INV_139_net_1));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_19_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB12_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_12__1_sqmuxa ), .ALn(
        AFLSDF_INV_119_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_19_set_net_1 ));
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_data_out8_73  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_9_[1]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_643 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_73_net_1 ));
    CFG4 #( .INIT(16'h7530) )  
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_6[2]  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_4_[2]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/mem_1_[2]_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/N_651 ), .D(
        \reg_apb_wrp_0/reg16x8_0/N_648 ), .Y(
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_6[2]_net_1 ));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_59  (.A(
        VCC), .B(GND), .C(VCC), .IPA(), .IPB(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[20] ), .IPC());
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_7_set_RNIONGP  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_7_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_235_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_8_rs[0] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_8_[0]_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_7_[0]  (.D(
        \CoreAPB3_0_APBmslave5_PWDATA[0] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB15_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_7__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_179_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_7_rs[0] ));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_265  (
        .A(VCC), .B(GND), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[25] ), 
        .IPB(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_ARBURST_HTRANS1_net[1] ), 
        .IPC(\hello_regs_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWRITE_net ));
    INV_BA AFLSDF_INV_7 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_127_net_1 ), .Y(
        AFLSDF_INV_7_net_1));
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_data_out8_99  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_10_[2]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_647 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_99_net_1 ));
    CFG3 #( .INIT(8'h02) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_125  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_3_[2]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_655 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_125_net_1 ));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_222  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[6] ), 
        .IPB(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[18] ), 
        .IPC());
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_data_out8_41  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_5_[3]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_653 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_41_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_4_[4]  (.D(
        \CoreAPB3_0_APBmslave5_PWDATA[4] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB14_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_4__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_140_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_4_rs[4] ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_186_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_70_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_186_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_186_rs_net_1 ));
    CFG3 #( .INIT(8'hF2) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_162  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_2_[2]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_642 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_162_i ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_137_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_2_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_137_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_137_rs_net_1 ));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_223  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[7] ), 
        .IPB(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[19] ), 
        .IPC());
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_data_out8_9  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_1_[0]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_651 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_9_net_1 ));
    CFG3 #( .INIT(8'hF2) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_218  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_14_[2]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_650 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_218_i ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_220_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_116_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_220_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_220_rs_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_14_[1]  (.D(
        \CoreAPB3_0_APBmslave5_PWDATA[1] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB12_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_14__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_217_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_14_rs[1] ));
    IP_INTERFACE \FCCC_0/CCC_INST/IP_INTERFACE_14  (.A(VCC), .B(VCC), 
        .C(VCC), .IPA(\FCCC_0/CCC_INST/NGMUX2_ARST_N_net ), .IPB(
        \FCCC_0/CCC_INST/GPD0_ARST_N_net ), .IPC(
        \FCCC_0/CCC_INST/PADDR_net[4] ));
    CFG3 #( .INIT(8'hF2) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_217  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_14_[1]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_650 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_217_i ));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_57  (.A(
        GND), .B(GND), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[11] ), .IPB(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[18] ), .IPC());
    SLE \reg_apb_wrp_0/reg16x8_0/mem_6_[4]  (.D(
        \CoreAPB3_0_APBmslave5_PWDATA[4] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB10_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_6__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_171_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_6_rs[4] ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_134_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_53_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_134_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_134_rs_net_1 ));
    CFG2 #( .INIT(4'h1) )  \reg_apb_wrp_0/reg16x8_0/data_out_RNO[1]  (
        .A(\reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_13[1]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_12[1]_net_1 ), .Y(
        \reg_apb_wrp_0/reg16x8_0/N_13_i_0 ));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_8_[0]  (.D(
        \CoreAPB3_0_APBmslave5_PWDATA[0] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB8_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_8__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_235_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_8_rs[0] ));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_165  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/SPI1_SS0_F2H_SCP_net ), .IPB(
        \hello_regs_MSS_0/MSS_ADLIB_INST/SPI1_SS3_F2H_SCP_net ), .IPC()
        );
    RGB \hello_regs_MSS_0/MSS_ADLIB_INST_RNIUO3B/U0_RGB1  (.An(
        \hello_regs_MSS_0/MSS_ADLIB_INST_RNIUO3B/U0_YNn ), .ENn(GND), 
        .YL(), .YR(
        \hello_regs_MSS_0/MSS_ADLIB_INST_RNIUO3B/U0_RGB1_YR ));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_1_[6]  (.D(
        \CoreAPB3_0_APBmslave5_PWDATA[6] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB14_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_1__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_158_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_1_rs[6] ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_66_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB9_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_8__1_sqmuxa ), .ALn(
        AFLSDF_INV_120_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_66_set_net_1 ));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_167  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(), .IPB(
        \hello_regs_MSS_0/MSS_ADLIB_INST/MMUART1_RTS_F2H_SCP_net ), 
        .IPC());
    CFG3 #( .INIT(8'hDF) )  \CoreAPB3_0/u_mux_p_to_b3/N_537_i  (.A(
        N_625), .B(CoreAPB3_0_APBmslave7_PREADY), .C(
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PADDR[17] ), .Y(N_537_i_0));
    CFG3 #( .INIT(8'h02) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_123  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_3_[1]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_655 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_123_net_1 ));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_76  (.A(
        VCC), .B(VCC), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[10] ), 
        .IPB(
        \hello_regs_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[17] ), 
        .IPC());
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_67_set_RNIB1UO  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_67_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_141_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_4_rs[5] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_4_[5]_net_1 ));
    CFG3 #( .INIT(8'h02) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_105  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_13_[1]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_646 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_105_net_1 ));
    CFG2_IP_BC 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/CFG_5  
        (.B(\CoreAPB3_0_APBmslave5_PWDATA[17] ), .C(GND), .IPB(
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/B_DIN_net[1] )
        , .IPC(
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/B_ADDR_net[2] )
        );
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_48_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB12_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_7__1_sqmuxa ), .ALn(
        AFLSDF_INV_121_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_48_set_net_1 ));
    INV_BA AFLSDF_INV_42 (.A(AFLSDF_INV_42_net_1), .Y(
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/B_DOUT_SRST_N_net )
        );
    INV_BA AFLSDF_INV_24 (.A(AFLSDF_INV_24_net_1), .Y(
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/B_BLK_net[0] )
        );
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[6].APB_8.GPOUT_reg[6]  (.D(
        \CoreAPB3_0_APBmslave5_PWDATA[6] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB12_rgbr_net_1 ), .EN(
        \CoreGPIO_0/GPOUT_reg35 ), .ALn(
        \hello_regs_MSS_0/MSS_ADLIB_INST_RNIUO3B/U0_RGB1_RGB4_rgbr_net_1 )
        , .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \GPIO_OUT_1_c[6] ));
    INV_BA AFLSDF_INV_93 (.A(AFLSDF_INV_93_net_1), .Y(
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/A_ARST_N_net )
        );
    SLE \reg_apb_wrp_0/reg16x8_0/mem_4_[0]  (.D(
        \CoreAPB3_0_APBmslave5_PWDATA[0] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB12_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_4__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_136_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_4_rs[0] ));
    RGB \FCCC_0/GL1_INST/U0_RGB1_RGB11  (.An(\FCCC_0/GL1_INST/U0_YNn ), 
        .ENn(GND), .YL(\FCCC_0/GL1_INST/U0_RGB1_RGB11_rgbl_net_1 ), 
        .YR(\FCCC_0/GL1_INST/U0_RGB1_RGB11_rgbr_net_1 ));
    INV_BA AFLSDF_INV_103 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_44_net_1 ), .Y(
        AFLSDF_INV_103_net_1));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_15_[5]  (.D(
        \CoreAPB3_0_APBmslave5_PWDATA[5] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB14_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_15__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_252_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_15_rs[5] ));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_0_[2]  (.D(
        \CoreAPB3_0_APBmslave5_PWDATA[2] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB14_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_0__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_145_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_0_rs[2] ));
    CFG3 #( .INIT(8'h80) )  
        \reg_apb_wrp_0/reg16x8_0/mem_0__1_sqmuxa_0_a2  (.A(
        \reg_apb_wrp_0/reg16x8_0/N_645 ), .B(N_637), .C(N_638), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_0__1_sqmuxa ));
    CFG2 #( .INIT(4'h1) )  \reg_apb_wrp_0/reg16x8_0/data_out_RNO[7]  (
        .A(\reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_13[7]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_12[7]_net_1 ), .Y(
        \reg_apb_wrp_0/reg16x8_0/N_84_i_0 ));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_179_rs_RNIU5CF  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_124_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_179_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_7_rs[0] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_7_[0]_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_109_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB2_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_13__1_sqmuxa ), .ALn(
        AFLSDF_INV_122_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_109_set_net_1 )
        );
    CFG3 #( .INIT(8'hF2) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_249  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_15_[2]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_654 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_249_i ));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_46  (.A(
        VCC), .B(GND), .C(VCC), .IPA(), .IPB(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[0] ), .IPC());
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_241  (
        .A(VCC), .B(GND), .C(GND), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[53] ), 
        .IPB(\hello_regs_MSS_0/MSS_ADLIB_INST/F_WSTRB_net[1] ), .IPC(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_BREADY_net ));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_6_[0]  (.D(
        \CoreAPB3_0_APBmslave5_PWDATA[0] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB10_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_6__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_203_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_6_rs[0] ));
    CFG3 #( .INIT(8'hF2) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_232  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_11_[5]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_649 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_232_i ));
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_data_out8_19  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_12_[3]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_644 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_19_net_1 ));
    CFG3 #( .INIT(8'hF2) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_128  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_3_[0]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_655 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_128_i ));
    CFG3 #( .INIT(8'h02) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_103  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_10_[6]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_647 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_103_net_1 ));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_46_set_RNIG5G01  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_46_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_159_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_1_rs[7] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_1_[7]_net_1 ));
    CFG3 #( .INIT(8'hF2) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_216  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_14_[0]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_650 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_216_i ));
    CFG4 #( .INIT(16'h0020) )  
        \reg_apb_wrp_0/reg16x8_0/WRITE_GEN.mem_5__2_i_a2[4]  (.A(
        \CoreAPB3_0_APBmslave5_PADDR[2] ), .B(
        \CoreAPB3_0_APBmslave5_PADDR[5] ), .C(
        \CoreAPB3_0_APBmslave5_PADDR[4] ), .D(
        \CoreAPB3_0_APBmslave5_PADDR[3] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/N_653 ));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_202_rs_RNIHN171  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_78_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_202_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_9_rs[6] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_9_[6]_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_181_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_126_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_181_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_181_rs_net_1 ));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/mem_14__RNI7C0H[2]  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_114_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_218_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_14_rs[2] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_14_[2]_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_24_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB6_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_5__1_sqmuxa ), .ALn(
        AFLSDF_INV_123_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_24_set_net_1 ));
    CFG3 #( .INIT(8'hF2) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_161  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_2_[1]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_642 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_161_i ));
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_data_out8_1  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_7_[7]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_641 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_1_net_1 ));
    CFG2 #( .INIT(4'h1) )  \reg_apb_wrp_0/reg16x8_0/data_out_RNO[5]  (
        .A(\reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_13[5]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_12[5]_net_1 ), .Y(
        \reg_apb_wrp_0/reg16x8_0/N_82_i_0 ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_5_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB7_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_8__1_sqmuxa ), .ALn(
        AFLSDF_INV_124_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_5_set_net_1 ));
    INV_BA AFLSDF_INV_86 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_net_1 ), .Y(
        AFLSDF_INV_86_net_1));
    INV_BA AFLSDF_INV_1 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_50_net_1 ), .Y(
        AFLSDF_INV_1_net_1));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_162  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/MGPIO12A_F2H_GPIN_net ), .IPB(
        \hello_regs_MSS_0/MSS_ADLIB_INST/MGPIO15A_F2H_GPIN_net ), .IPC(
        ));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_3  (.A(
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[1] ), .B(
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[8] ), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[1] ), .IPB(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[8] ), .IPC());
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_150  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/MGPIO2A_F2H_GPIN_net ), .IPB(
        \hello_regs_MSS_0/MSS_ADLIB_INST/SPI0_SDI_F2H_SCP_net ), .IPC()
        );
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_250_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_56_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_250_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_250_rs_net_1 ));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_230  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[28] ), 
        .IPB(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[40] ), 
        .IPC());
    CFG2 #( .INIT(4'h8) )  \COREAPBLSRAM_0/wen_0_a2_0  (.A(
        CoreAPB3_0_APBmslave5_PENABLE), .B(
        CoreAPB3_0_APBmslave5_PWRITE), .Y(N_638));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_45_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB9_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_5__1_sqmuxa ), .ALn(
        AFLSDF_INV_125_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_45_set_net_1 ));
    CFG4 #( .INIT(16'h7350) )  
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_5[3]  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_0_[3]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/mem_7_[3]_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/N_645 ), .D(
        \reg_apb_wrp_0/reg16x8_0/N_641 ), .Y(
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_5[3]_net_1 ));
    CFG3 #( .INIT(8'hAC) )  
        \CoreAPB3_0/u_mux_p_to_b3/PRDATA_m3_i_m3_0  (.A(
        \COREAPBLSRAM_0.PRDATA_reg[0] ), .B(
        \COREAPBLSRAM_0.lsram_width32_PRDATA[0] ), .C(N_354), .Y(
        \CoreAPB3_0/u_mux_p_to_b3/PRDATA_N_8_0 ));
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_data_out8_95  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_11_[7]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_649 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_95_net_1 ));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_196  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[0] ), 
        .IPB(\hello_regs_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[12] )
        , .IPC());
    INV_BA AFLSDF_INV_6 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_42_net_1 ), .Y(
        AFLSDF_INV_6_net_1));
    CFG3 #( .INIT(8'h02) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_108  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_13_[4]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_646 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_108_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_211_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_107_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_211_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_211_rs_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_37_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB4_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_2__1_sqmuxa ), .ALn(
        AFLSDF_INV_126_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_37_set_net_1 ));
    CFG3 #( .INIT(8'hF2) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_224  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_11_[1]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_649 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_224_i ));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_255  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[3] ), 
        .IPB(\hello_regs_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[15] )
        , .IPC());
    IOENFF_BYPASS \GPIO_OUT_1_obuf[1]/U0/U_IOENFF  (.A(
        \GPIO_OUT_1_obuf[1]/U0/EOUT1 ), .Y(
        \GPIO_OUT_1_obuf[1]/U0/EOUT ));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/mem_3__RNIGG5O[2]  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_125_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_130_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_3_rs[2] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_3_[2]_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_3_[2]  (.D(
        \CoreAPB3_0_APBmslave5_PWDATA[2] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB12_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_3__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_130_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_3_rs[2] ));
    SLE_IP_EN 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/FF_22  
        (.EN(VCC), .IPENn());
    SLE \reg_apb_wrp_0/reg16x8_0/mem_9_[3]  (.D(
        \CoreAPB3_0_APBmslave5_PWDATA[3] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB16_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_9__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_196_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_9_rs[3] ));
    INV_BA AFLSDF_INV_95 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_67_net_1 ), .Y(
        AFLSDF_INV_95_net_1));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_266  (
        .A(VCC), .B(GND), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[26] ), 
        .IPB(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_ARLOCK_HMASTLOCK1_net[0] ), 
        .IPC());
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_133_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_51_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_133_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_133_rs_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_15_[0]  (.D(
        \CoreAPB3_0_APBmslave5_PWDATA[0] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB16_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_15__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_251_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_15_rs[0] ));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_176  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/MGPIO26B_F2H_GPIN_net ), .IPB(
        \hello_regs_MSS_0/MSS_ADLIB_INST/MMUART0_CTS_F2H_SCP_net ), 
        .IPC());
    CFG4 #( .INIT(16'h7350) )  
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_0[4]  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_11_[4]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/mem_10_[4]_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/N_649 ), .D(
        \reg_apb_wrp_0/reg16x8_0/N_647 ), .Y(
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_0[4]_net_1 ));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_155  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(), .IPB(
        \hello_regs_MSS_0/MSS_ADLIB_INST/MGPIO8A_F2H_GPIN_net ), .IPC()
        );
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/mem_2__RNIE2FF[6]  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_37_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_166_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_2_rs[6] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_2_[6]_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_248_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_58_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_248_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_248_rs_net_1 ));
    INV_BA AFLSDF_INV_41 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_88_net_1 ), .Y(
        AFLSDF_INV_41_net_1));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_7_[2]  (.D(
        \CoreAPB3_0_APBmslave5_PWDATA[2] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB12_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_7__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_183_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_7_rs[2] ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_178_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_103_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_178_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_178_rs_net_1 ));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/mem_15__RNIPFOP[0]  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_57_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_251_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_15_rs[0] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_15_[0]_net_1 ));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_157  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/SPI0_SS2_F2H_SCP_net ), .IPB()
        , .IPC());
    CFG4 #( .INIT(16'h7530) )  
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_4[7]  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_6_[7]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/mem_3_[7]_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/N_655 ), .D(
        \reg_apb_wrp_0/reg16x8_0/N_652 ), .Y(
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_4[7]_net_1 ));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_75  (.A(
        VCC), .B(VCC), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[9] ), 
        .IPB(
        \hello_regs_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[16] ), 
        .IPC());
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_24  (.A(
        GND), .B(VCC), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[0] ), .IPB(), 
        .IPC());
    CFG3 #( .INIT(8'hF2) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_204  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_9_[7]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_643 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_204_i ));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_220  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[4] ), 
        .IPB(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[16] ), 
        .IPC());
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/mem_8__RNIPMA31[1]  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_5_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_237_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_8_rs[1] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_8_[1]_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_10_[4]  (.D(
        \CoreAPB3_0_APBmslave5_PWDATA[4] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB7_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_10__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_174_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_10_rs[4] ));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_281  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PADDR_net[4] ), 
        .IPB(
        \hello_regs_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[8] ), 
        .IPC());
    CFG4 #( .INIT(16'h7350) )  
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_5[7]  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_0_[7]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/mem_7_[7]_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/N_645 ), .D(
        \reg_apb_wrp_0/reg16x8_0/N_641 ), .Y(
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_5[7]_net_1 ));
    CFG3 #( .INIT(8'hF2) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_219  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_14_[3]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_650 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_219_i ));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_9_[4]  (.D(
        \CoreAPB3_0_APBmslave5_PWDATA[4] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB18_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_9__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_198_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_9_rs[4] ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_49_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB13_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_3__1_sqmuxa ), .ALn(
        AFLSDF_INV_127_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_49_set_net_1 ));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_144  (
        .A(FCCC_0_LOCK), .B(VCC), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/FAB_PLL_LOCK_net ), .IPB(), 
        .IPC());
    INV_BA AFLSDF_INV_146 (.A(\FCCC_0/GL1_net ), .Y(
        AFLSDF_INV_146_net_1));
    RGB \FCCC_0/GL1_INST/U0_RGB1_RGB13  (.An(
        \FCCC_0/GL1_INST/U0_YNn_GSouth ), .ENn(GND), .YL(
        \FCCC_0/GL1_INST/U0_RGB1_RGB13_rgbl_net_1 ), .YR(
        \FCCC_0/GL1_INST/U0_RGB1_RGB13_rgbr_net_1 ));
    CFG2_IP_BC 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/CFG_14  
        (.B(\CoreAPB3_0_APBmslave5_PWDATA[11] ), .C(
        \CoreAPB3_0_APBmslave5_PADDR[1] ), .IPB(
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/A_DIN_net[12] )
        , .IPC(
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/A_ADDR_net[6] )
        );
    SLE \reg_apb_wrp_0/reg16x8_0/mem_8_[2]  (.D(
        \CoreAPB3_0_APBmslave5_PWDATA[2] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB5_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_8__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_239_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_8_rs[2] ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_31_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB4_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_2__1_sqmuxa ), .ALn(
        AFLSDF_INV_128_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_31_set_net_1 ));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_234  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[32] ), 
        .IPB(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[44] ), 
        .IPC());
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_data_out8_15  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_1_[3]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_651 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_15_net_1 ));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_168  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/MMUART1_CTS_F2H_SCP_net ), 
        .IPB(), .IPC());
    CFG2 #( .INIT(4'h8) )  
        \CoreAPB3_0/u_mux_p_to_b3/PRDATA_0_iv_0_a2_2_0[2]  (.A(N_639), 
        .B(\GPIO_OUT_1_c[2] ), .Y(
        \CoreAPB3_0/u_mux_p_to_b3/PRDATA_0_iv_0_a2_2_0[2]_net_1 ));
    INV_BA AFLSDF_INV_129 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_62_net_1 ), .Y(
        AFLSDF_INV_129_net_1));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_98  (.A(
        VCC), .B(VCC), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/MDIF_net ), .IPB(), .IPC());
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_45  (.A(
        GND), .B(GND), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[28] ), .IPB(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_ENABLE_net ), .IPC());
    CFG4 #( .INIT(16'h7530) )  
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_7[1]  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_8_[1]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/mem_5_[1]_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/N_653 ), .D(N_639), .Y(
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_7[1]_net_1 ));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_36  (.A(
        GND), .B(VCC), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[19] ), .IPB(), 
        .IPC());
    CFG4 #( .INIT(16'hECA0) )  \CoreAPB3_0/u_mux_p_to_b3/PRDATA_0[18]  
        (.A(\CoreAPB3_0/u_mux_p_to_b3/N_636 ), .B(
        \COREAPBLSRAM_0.PRDATA4 ), .C(\COREAPBLSRAM_0.PRDATA_reg[18] ), 
        .D(\COREAPBLSRAM_0.lsram_width32_PRDATA[18] ), .Y(
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[18] ));
    INV_BA AFLSDF_INV_77 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_71_net_1 ), .Y(
        AFLSDF_INV_77_net_1));
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_data_out8_54  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_7_[5]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_641 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_54_net_1 ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[3].APB_8.GPOUT_reg[3]  (.D(
        \CoreAPB3_0_APBmslave5_PWDATA[3] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB12_rgbr_net_1 ), .EN(
        \CoreGPIO_0/GPOUT_reg35 ), .ALn(
        \hello_regs_MSS_0/MSS_ADLIB_INST_RNIUO3B/U0_RGB1_RGB4_rgbr_net_1 )
        , .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \GPIO_OUT_1_c[3] ));
    CFG4 #( .INIT(16'hFEFA) )  
        \CoreAPB3_0/u_mux_p_to_b3/PRDATA_0_iv_0[1]  (.A(
        \CoreAPB3_0/u_mux_p_to_b3/N_585 ), .B(
        \COREAPBLSRAM_0.PRDATA_reg[1] ), .C(
        \CoreAPB3_0/u_mux_p_to_b3/PRDATA_0_iv_0_0[1]_net_1 ), .D(
        \CoreAPB3_0/u_mux_p_to_b3/N_636 ), .Y(
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[1] ));
    INV_BA AFLSDF_INV_144 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_122_net_1 ), .Y(
        AFLSDF_INV_144_net_1));
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_data_out8_43  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_5_[2]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_653 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_43_net_1 ));
    CFG4 #( .INIT(16'hEAC0) )  
        \CoreAPB3_0/u_mux_p_to_b3/PRDATA_0_iv_0_0[7]  (.A(
        \COREAPBLSRAM_0.PRDATA_reg[7] ), .B(
        \CoreAPB3_0/u_mux_p_to_b3/PRDATA_0_iv_0_a2_2_0[7]_net_1 ), .C(
        \CoreAPB3_0.u_mux_p_to_b3.PRDATA_0_iv_0_a2_3_5[1] ), .D(
        \CoreAPB3_0/u_mux_p_to_b3/N_636 ), .Y(
        \CoreAPB3_0/u_mux_p_to_b3/PRDATA_0_iv_0_0[7]_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_62_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB14_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_15__1_sqmuxa ), .ALn(
        AFLSDF_INV_129_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_62_set_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_16_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB18_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_12__1_sqmuxa ), .ALn(
        AFLSDF_INV_130_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_16_set_net_1 ));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_152  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/MGPIO3A_F2H_GPIN_net ), .IPB(
        \hello_regs_MSS_0/MSS_ADLIB_INST/SPI0_SDO_F2H_SCP_net ), .IPC()
        );
    CFG3 #( .INIT(8'hF2) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_238  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_12_[0]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_644 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_238_i ));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_4_[2]  (.D(
        \CoreAPB3_0_APBmslave5_PWDATA[2] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB18_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_4__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_138_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_4_rs[2] ));
    CFG2_IP_BC 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/CFG_24  
        (.B(\CoreAPB3_0_APBmslave5_PWDATA[6] ), .C(
        \CoreAPB3_0_APBmslave5_PADDR[4] ), .IPB(
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/A_DIN_net[6] )
        , .IPC(
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/A_ADDR_net[9] )
        );
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_101  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/RCGF_net[1] ), .IPB(
        \hello_regs_MSS_0/MSS_ADLIB_INST/RCGF_net[8] ), .IPC());
    CFG3 #( .INIT(8'hF2) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_237  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_8_[1]_net_1 ), .B(N_639), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_237_i ));
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_data_out8  (
        .A(\reg_apb_wrp_0/reg16x8_0/mem_4_[0]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_648 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_net_1 ));
    RGB \FCCC_0/GL1_INST/U0_RGB1_RGB19  (.An(
        \FCCC_0/GL1_INST/U0_YNn_GSouth ), .ENn(GND), .YL(), .YR(
        \FCCC_0/GL1_INST/U0_RGB1_RGB19_rgbr_net_1 ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[7].APB_8.GPOUT_reg[7]  (.D(
        \CoreAPB3_0_APBmslave5_PWDATA[7] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB12_rgbr_net_1 ), .EN(
        \CoreGPIO_0/GPOUT_reg35 ), .ALn(
        \hello_regs_MSS_0/MSS_ADLIB_INST_RNIUO3B/U0_RGB1_RGB4_rgbr_net_1 )
        , .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \GPIO_OUT_1_c[7] ));
    CFG4 #( .INIT(16'hECA0) )  \CoreAPB3_0/u_mux_p_to_b3/PRDATA_0[22]  
        (.A(\CoreAPB3_0/u_mux_p_to_b3/N_636 ), .B(
        \COREAPBLSRAM_0.PRDATA4 ), .C(\COREAPBLSRAM_0.PRDATA_reg[22] ), 
        .D(\COREAPBLSRAM_0.lsram_width32_PRDATA[22] ), .Y(
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[22] ));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_144_rs_RNI28UM  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_81_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_144_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_0_rs[1] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_0_[1]_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_9_[0]  (.D(
        \CoreAPB3_0_APBmslave5_PWDATA[0] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB19_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_9__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_190_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_9_rs[0] ));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_6_[2]  (.D(
        \CoreAPB3_0_APBmslave5_PWDATA[2] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB11_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_6__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_207_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_6_rs[2] ));
    INV_BA AFLSDF_INV_141 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_46_net_1 ), .Y(
        AFLSDF_INV_141_net_1));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_132_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_49_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_132_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_132_rs_net_1 ));
    SLE_IP_CLK 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/FF_24  
        (.CLK(\FCCC_0/GL1_INST/U0_RGB1_RGB0_rgbr_net_1 ), .IPCLKn(
        AFLSDF_INV_131_net_1));
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_data_out8_57  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_15_[0]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_654 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_57_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_229_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_54_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_229_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_229_rs_net_1 ));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_224  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[8] ), 
        .IPB(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[20] ), 
        .IPC());
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_18_set_RNILK0L  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_18_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_242_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_12_rs[2] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_12_[2]_net_1 ));
    CFG4 #( .INIT(16'h7530) )  
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_4[1]  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_6_[1]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/mem_3_[1]_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/N_655 ), .D(
        \reg_apb_wrp_0/reg16x8_0/N_652 ), .Y(
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_4[1]_net_1 ));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_61  (.A(
        GND), .B(VCC), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[22] ), .IPB(), 
        .IPC());
    SLE \reg_apb_wrp_0/reg16x8_0/mem_0_[5]  (.D(
        \CoreAPB3_0_APBmslave5_PWDATA[5] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB13_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_0__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_149_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_0_rs[5] ));
    SLE \COREAPBLSRAM_0/PRDATA_reg[29]  (.D(
        \COREAPBLSRAM_0.lsram_width32_PRDATA[29] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB10_rgbr_net_1 ), .EN(
        \COREAPBLSRAM_0.PRDATA4 ), .ALn(
        \hello_regs_MSS_0/MSS_ADLIB_INST_RNIUO3B/U0_RGB1_RGB2_rgbr_net_1 )
        , .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \COREAPBLSRAM_0.PRDATA_reg[29] ));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_28  (.A(
        GND), .B(GND), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[4] ), .IPB(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[11] ), .IPC());
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_256  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[4] ), 
        .IPB(\hello_regs_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[16] )
        , .IPC());
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_84  (.A(
        VCC), .B(VCC), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[25] ), 
        .IPB(\hello_regs_MSS_0/MSS_ADLIB_INST/RXDF_net[0] ), .IPC());
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_147_rs_RNI3C1M  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_80_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_147_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_0_rs[0] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_0_[0]_net_1 ));
    INV_BA AFLSDF_INV_79 (.A(\hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        AFLSDF_INV_79_net_1));
    CFG4 #( .INIT(16'h2000) )  
        \CoreAPB3_0/u_mux_p_to_b3/PREADY_0_i_a2_1  (.A(
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PADDR[18] ), .B(
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PADDR[19] ), .C(
        hello_regs_MSS_0_FIC_0_APB_MASTER_PSELx), .D(
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PADDR[16] ), .Y(N_625));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_184  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/MGPIO28B_F2H_GPIN_net ), .IPB(
        \hello_regs_MSS_0/MSS_ADLIB_INST/MGPIO31B_F2H_GPIN_net ), .IPC(
        ));
    INV_BA AFLSDF_INV_92 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_20_net_1 ), .Y(
        AFLSDF_INV_92_net_1));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_27_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB1_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_2__1_sqmuxa ), .ALn(
        AFLSDF_INV_132_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_27_set_net_1 ));
    CFG3 #( .INIT(8'hF2) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_140  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_4_[4]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_648 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_140_i ));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_193  (
        .A(GND), .B(VCC), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_AWID_HSEL0_net[1] ), .IPB(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[9] ), 
        .IPC(\hello_regs_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[21] )
        );
    CFG4 #( .INIT(16'h7530) )  
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_0_7[6]  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_8_[6]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/mem_5_[6]_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/N_653 ), .D(N_639), .Y(
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_0_7[6]_net_1 ));
    CFG3 #( .INIT(8'hF2) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_236  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_11_[7]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_649 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_236_i ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_8_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB15_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_4__1_sqmuxa ), .ALn(
        AFLSDF_INV_133_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_8_set_net_1 ));
    SLE_IP_EN 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/FF_7  
        (.EN(VCC), .IPENn(AFLSDF_INV_134_net_1));
    INV_BA AFLSDF_INV_119 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_19_net_1 ), .Y(
        AFLSDF_INV_119_net_1));
    RGB \FCCC_0/GL1_INST/U0_RGB1_RGB14  (.An(
        \FCCC_0/GL1_INST/U0_YNn_GSouth ), .ENn(GND), .YL(
        \FCCC_0/GL1_INST/U0_RGB1_RGB14_rgbl_net_1 ), .YR(
        \FCCC_0/GL1_INST/U0_RGB1_RGB14_rgbr_net_1 ));
    CFG2_IP_BC 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/CFG_7  
        (.B(\CoreAPB3_0_APBmslave5_PWDATA[25] ), .C(GND), .IPB(
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/B_DIN_net[10] )
        , .IPC(
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/B_ADDR_net[3] )
        );
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_38_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB9_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_6__1_sqmuxa ), .ALn(
        AFLSDF_INV_135_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_38_set_net_1 ));
    INV_BA AFLSDF_INV_17 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_53_net_1 ), .Y(
        AFLSDF_INV_17_net_1));
    CFG4 #( .INIT(16'h7350) )  
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_5[0]  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_0_[0]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/mem_7_[0]_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/N_645 ), .D(
        \reg_apb_wrp_0/reg16x8_0/N_641 ), .Y(
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_5[0]_net_1 ));
    CFG4 #( .INIT(16'h7350) )  
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_5[2]  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_0_[2]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/mem_7_[2]_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/N_645 ), .D(
        \reg_apb_wrp_0/reg16x8_0/N_641 ), .Y(
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_5[2]_net_1 ));
    RGB \hello_regs_MSS_0/MSS_ADLIB_INST_RNIUO3B/U0_RGB1_RGB3  (.An(
        \hello_regs_MSS_0/MSS_ADLIB_INST_RNIUO3B/U0_YNn ), .ENn(GND), 
        .YL(), .YR(
        \hello_regs_MSS_0/MSS_ADLIB_INST_RNIUO3B/U0_RGB1_RGB3_rgbr_net_1 )
        );
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_173  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/MMUART1_TXD_F2H_SCP_net ), 
        .IPB(\hello_regs_MSS_0/MSS_ADLIB_INST/MGPIO18B_F2H_GPIN_net ), 
        .IPC());
    CFG3 #( .INIT(8'hF2) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_240  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_12_[1]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_644 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_240_i ));
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_data_out8_24  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_5_[6]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_653 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_24_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_3_[5]  (.D(
        \CoreAPB3_0_APBmslave5_PWDATA[5] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB13_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_3__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_133_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_3_rs[5] ));
    CFG3 #( .INIT(8'h08) )  \COREAPBLSRAM_0/g0_0  (.A(
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PADDR[17] ), .B(
        CoreAPB3_0_APBmslave5_PENABLE), .C(
        CoreAPB3_0_APBmslave5_PWRITE), .Y(
        \COREAPBLSRAM_0.PRDATA4_0_a2_0 ));
    CFG3 #( .INIT(8'hF2) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_170  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_10_[2]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_647 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_170_i ));
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_data_out8_51  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_3_[5]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_655 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_51_net_1 ));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_158  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/MGPIO10A_F2H_GPIN_net ), .IPB(
        ), .IPC());
    SLE \COREAPBLSRAM_0/PRDATA_reg[30]  (.D(
        \COREAPBLSRAM_0.lsram_width32_PRDATA[30] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB9_rgbr_net_1 ), .EN(
        \COREAPBLSRAM_0.PRDATA4 ), .ALn(
        \hello_regs_MSS_0/MSS_ADLIB_INST_RNIUO3B/U0_RGB1_RGB1_rgbr_net_1 )
        , .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \COREAPBLSRAM_0.PRDATA_reg[30] ));
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_data_out8_76  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_9_[4]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_643 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_76_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_0_[7]  (.D(
        \CoreAPB3_0_APBmslave5_PWDATA[7] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB17_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_0__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_151_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_0_rs[7] ));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_35  (.A(
        VCC), .B(GND), .C(VCC), .IPA(), .IPB(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[18] ), .IPC());
    INV_BA AFLSDF_INV_67 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_97_net_1 ), .Y(
        AFLSDF_INV_67_net_1));
    CFG3 #( .INIT(8'h80) )  
        \reg_apb_wrp_0/reg16x8_0/mem_14__1_sqmuxa_0_a2_0_a2  (.A(
        \reg_apb_wrp_0/reg16x8_0/N_650 ), .B(N_637), .C(N_638), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_14__1_sqmuxa ));
    CFG3 #( .INIT(8'h80) )  
        \reg_apb_wrp_0/reg16x8_0/mem_8__1_sqmuxa_0_a2_0_a2  (.A(N_639), 
        .B(N_637), .C(N_638), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_8__1_sqmuxa ));
    CFG2 #( .INIT(4'h2) )  \reg_apb_wrp_0/rd_enable_0_a2_0  (.A(N_625), 
        .B(\hello_regs_MSS_0_FIC_0_APB_MASTER_PADDR[17] ), .Y(N_637));
    INV_BA AFLSDF_INV_107 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_107_net_1 ), .Y(
        AFLSDF_INV_107_net_1));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_21_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB14_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_12__1_sqmuxa ), .ALn(
        AFLSDF_INV_136_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_21_set_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_7_[5]  (.D(
        \CoreAPB3_0_APBmslave5_PWDATA[5] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB15_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_7__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_229_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_7_rs[5] ));
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_data_out8_27  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_2_[1]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_642 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_27_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_204_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_79_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_204_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_204_rs_net_1 ));
    CFG1_IP_B 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/CFG_35  
        (.B(GND), .IPB(
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/B_DIN_net[17] )
        );
    SLE_IP_EN 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/FF_9  
        (.EN(VCC), .IPENn(AFLSDF_INV_137_net_1));
    CFG4 #( .INIT(16'h7530) )  
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_6[3]  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_4_[3]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/mem_1_[3]_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/N_651 ), .D(
        \reg_apb_wrp_0/reg16x8_0/N_648 ), .Y(
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_6[3]_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_7_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB8_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_8__1_sqmuxa ), .ALn(
        AFLSDF_INV_138_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_7_set_net_1 ));
    CFG3 #( .INIT(8'hF2) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_253  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_15_[6]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_654 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_253_i ));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_88  (.A(
        VCC), .B(VCC), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[29] ), 
        .IPB(\hello_regs_MSS_0/MSS_ADLIB_INST/RXDF_net[4] ), .IPC());
    sdf_IOPAD_TRI \GPIO_OUT_1_obuf[3]/U0/U_IOPAD  (.PAD(GPIO_OUT_1[3]), 
        .D(\GPIO_OUT_1_obuf[3]/U0/DOUT ), .E(
        \GPIO_OUT_1_obuf[3]/U0/EOUT ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_35_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB2_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_2__1_sqmuxa ), .ALn(
        AFLSDF_INV_139_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_35_set_net_1 ));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_108_set_RNI53MS  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_108_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_212_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_13_rs[4] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_13_[4]_net_1 ));
    INV_BA AFLSDF_INV_26 (.A(AFLSDF_INV_26_net_1), .Y(
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/B_BLK_net[2] )
        );
    INV_BA AFLSDF_INV_19 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_32_net_1 ), .Y(
        AFLSDF_INV_19_net_1));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_8_[5]  (.D(
        \CoreAPB3_0_APBmslave5_PWDATA[5] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB8_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_8__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_184_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_8_rs[5] ));
    INV_BA AFLSDF_INV_142 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_39_net_1 ), .Y(
        AFLSDF_INV_142_net_1));
    INV_BA AFLSDF_INV_91 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_79_net_1 ), .Y(
        AFLSDF_INV_91_net_1));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_11_[4]  (.D(
        \CoreAPB3_0_APBmslave5_PWDATA[4] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB4_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_11__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_230_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_11_rs[4] ));
    IOOUTFF_BYPASS \MSS_RESET_N_M2F_obuf/U0/U_IOOUTFF  (.A(
        \MSS_RESET_N_M2F_obuf/U0/DOUT1 ), .Y(
        \MSS_RESET_N_M2F_obuf/U0/DOUT ));
    CFG3 #( .INIT(8'h02) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_110  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_13_[6]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_646 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_110_net_1 ));
    IP_INTERFACE \FCCC_0/CCC_INST/IP_INTERFACE_17  (.A(VCC), .B(VCC), 
        .C(VCC), .IPA(), .IPB(\FCCC_0/CCC_INST/GPD3_ARST_N_net ), .IPC(
        \FCCC_0/CCC_INST/PADDR_net[7] ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_167_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_39_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_167_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_167_rs_net_1 ));
    CFG3 #( .INIT(8'hF2) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_144  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_0_[1]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_645 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_144_i ));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_3_[7]  (.D(
        \CoreAPB3_0_APBmslave5_PWDATA[7] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB13_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_3__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_135_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_3_rs[7] ));
    CFG3 #( .INIT(8'hF2) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_245  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_12_[5]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_644 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_245_i ));
    CFG3 #( .INIT(8'hF2) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_239  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_8_[2]_net_1 ), .B(N_639), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_239_i ));
    CFG4 #( .INIT(16'hBFFF) )  \COREAPBLSRAM_0/PREADY_reg6_i  (.A(
        CoreAPB3_0_APBmslave5_PENABLE), .B(
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PADDR[17] ), .C(N_625), .D(
        \COREAPBLSRAM_0/PREADY_reg6_0_a2_0_net_1 ), .Y(
        \COREAPBLSRAM_0/PREADY_reg6_i_0 ));
    INV_BA AFLSDF_INV_69 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_118_net_1 ), .Y(
        AFLSDF_INV_69_net_1));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_9_[2]  (.D(
        \CoreAPB3_0_APBmslave5_PWDATA[2] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB18_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_9__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_194_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_9_rs[2] ));
    CFG4 #( .INIT(16'hFFFE) )  
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_0_12[6]  (.A(
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_0_1[6]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_0_3[6]_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_0_2[6]_net_1 ), .D(
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_0_0[6]_net_1 ), .Y(
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_0_12[6]_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_222_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_118_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_222_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_222_rs_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_164_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_33_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_164_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_164_rs_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_4_[5]  (.D(
        \CoreAPB3_0_APBmslave5_PWDATA[5] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB14_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_4__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_141_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_4_rs[5] ));
    INV_BA AFLSDF_INV_80 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_124_net_1 ), .Y(
        AFLSDF_INV_80_net_1));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_140  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/RX_EV_net ), .IPB(
        \hello_regs_MSS_0/MSS_ADLIB_INST/USER_MSS_GPIO_RESET_N_net ), 
        .IPC());
    CFG3 #( .INIT(8'h02) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_127  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_3_[3]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_655 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_127_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_12_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB9_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_5__1_sqmuxa ), .ALn(
        AFLSDF_INV_140_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_12_set_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_247_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_23_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_247_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_247_rs_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_213_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_109_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_213_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_213_rs_net_1 ));
    CFG3 #( .INIT(8'hF2) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_210  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_13_[2]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_646 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_210_i ));
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_data_out8_21  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_12_[5]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_644 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_21_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_7_[7]  (.D(
        \CoreAPB3_0_APBmslave5_PWDATA[7] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB16_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_7__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_233_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_7_rs[7] ));
    CFG3 #( .INIT(8'hF2) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_174  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_10_[4]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_647 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_174_i ));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_2_[6]  (.D(
        \CoreAPB3_0_APBmslave5_PWDATA[6] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB5_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_2__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_166_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_2_rs[6] ));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_15_[6]  (.D(
        \CoreAPB3_0_APBmslave5_PWDATA[6] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB12_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_15__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_253_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_15_rs[6] ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_46_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB16_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_1__1_sqmuxa ), .ALn(
        AFLSDF_INV_141_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_46_set_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_6_[5]  (.D(
        \CoreAPB3_0_APBmslave5_PWDATA[5] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB9_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_6__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_173_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_6_rs[5] ));
    SLE \reg_apb_wrp_0/reg16x8_0/data_out[2]  (.D(
        \reg_apb_wrp_0/reg16x8_0/N_15_i_0 ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB11_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/rd_enable ), .ALn(
        \hello_regs_MSS_0/MSS_ADLIB_INST_RNIUO3B/U0_RGB1_RGB3_rgbr_net_1 )
        , .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreAPB3_0_APBmslave5_PRDATA[2] ));
    IOOUTFF_BYPASS \GPIO_OUT_1_obuf[1]/U0/U_IOOUTFF  (.A(
        \GPIO_OUT_1_obuf[1]/U0/DOUT1 ), .Y(
        \GPIO_OUT_1_obuf[1]/U0/DOUT ));
    CFG3 #( .INIT(8'hF2) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_186  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_8_[6]_net_1 ), .B(N_639), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_186_i ));
    INV_BA AFLSDF_INV_74 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_52_net_1 ), .Y(
        AFLSDF_INV_74_net_1));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_39_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB3_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_2__1_sqmuxa ), .ALn(
        AFLSDF_INV_142_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_39_set_net_1 ));
    CFG4 #( .INIT(16'hFFFE) )  
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_12[2]  (.A(
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_1[2]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_3[2]_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_2[2]_net_1 ), .D(
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_0[2]_net_1 ), .Y(
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_12[2]_net_1 ));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_245  (
        .A(VCC), .B(GND), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[57] ), 
        .IPB(\hello_regs_MSS_0/MSS_ADLIB_INST/F_WSTRB_net[5] ), .IPC());
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_6  (.A(
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[4] ), .B(
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[11] ), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[4] ), .IPB(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[11] ), .IPC());
    SLE \reg_apb_wrp_0/reg16x8_0/mem_8_[7]  (.D(
        \CoreAPB3_0_APBmslave5_PWDATA[7] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB7_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_8__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_188_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_8_rs[7] ));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_199  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[3] ), 
        .IPB(\hello_regs_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[15] )
        , .IPC());
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_231_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_3_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_231_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_231_rs_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_135_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_55_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_135_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_135_rs_net_1 ));
    CFG3 #( .INIT(8'h02) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_107  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_13_[3]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_646 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_107_net_1 ));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_19  (.A(
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[24] ), .B(
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[31] ), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[24] ), .IPB(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[31] ), .IPC());
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_data_out8_34  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_6_[3]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_652 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_34_net_1 ));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_145  (
        .A(GND), .B(VCC), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/SLEEPHOLDREQ_net ), .IPB(), 
        .IPC());
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_28_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB10_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_6__1_sqmuxa ), .ALn(
        AFLSDF_INV_143_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_28_set_net_1 ));
    CFG4 #( .INIT(16'h7350) )  
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_0[5]  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_11_[5]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/mem_10_[5]_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/N_649 ), .D(
        \reg_apb_wrp_0/reg16x8_0/N_647 ), .Y(
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_0[5]_net_1 ));
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_data_out8_88  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_11_[0]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_649 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_88_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_122_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB18_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_6__1_sqmuxa ), .ALn(
        AFLSDF_INV_144_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_122_set_net_1 )
        );
    RGB \hello_regs_MSS_0/MSS_ADLIB_INST_RNIUO3B/U0_RGB1_RGB0  (.An(
        \hello_regs_MSS_0/MSS_ADLIB_INST_RNIUO3B/U0_YNn ), .ENn(GND), 
        .YL(), .YR(
        \hello_regs_MSS_0/MSS_ADLIB_INST_RNIUO3B/U0_RGB1_RGB0_rgbr_net_1 )
        );
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_179  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(), .IPB(
        \hello_regs_MSS_0/MSS_ADLIB_INST/MGPIO21B_F2H_GPIN_net ), .IPC(
        ));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_147  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/I2C1_SDA_F2H_SCP_net ), .IPB(
        \hello_regs_MSS_0/MSS_ADLIB_INST/MGPIO4A_F2H_GPIN_net ), .IPC()
        );
    RGB \FCCC_0/GL1_INST/U0_RGB1_RGB16  (.An(
        \FCCC_0/GL1_INST/U0_YNn_GSouth ), .ENn(GND), .YL(
        \FCCC_0/GL1_INST/U0_RGB1_RGB16_rgbl_net_1 ), .YR(
        \FCCC_0/GL1_INST/U0_RGB1_RGB16_rgbr_net_1 ));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_74  (.A(
        VCC), .B(VCC), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[8] ), 
        .IPB(), .IPC());
    SLE_IP_EN 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/FF_27  
        (.EN(VCC), .IPENn());
    SLE \reg_apb_wrp_0/reg16x8_0/mem_10_[5]  (.D(
        \CoreAPB3_0_APBmslave5_PWDATA[5] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB7_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_10__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_176_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_10_rs[5] ));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_17  (.A(
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[22] ), .B(
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[29] ), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[22] ), .IPB(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[29] ), .IPC());
    INV_BA AFLSDF_INV_4 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_125_net_1 ), .Y(
        AFLSDF_INV_4_net_1));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_4_[7]  (.D(
        \CoreAPB3_0_APBmslave5_PWDATA[7] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB15_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_4__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_185_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_4_rs[7] ));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_222_rs_RNIAICF  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_118_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_222_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_14_rs[6] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_14_[6]_net_1 ));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_6_set_RNIPDKE  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_6_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_139_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_4_rs[3] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_4_[3]_net_1 ));
    CFG3 #( .INIT(8'h02) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_114  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_14_[2]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_650 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_114_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_252_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_62_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_252_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_252_rs_net_1 ));
    CFG3 #( .INIT(8'hF2) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_215  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_13_[7]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_646 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_215_i ));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_123_set_RNILUEL  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_123_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_129_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_3_rs[1] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_3_[1]_net_1 ));
    CFG3 #( .INIT(8'h08) )  
        \CoreAPB3_0/u_mux_p_to_b3/PRDATA_0_iv_0_a2_0[1]  (.A(N_625), 
        .B(\CoreAPB3_0_APBmslave5_PRDATA[1] ), .C(
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PADDR[17] ), .Y(
        \CoreAPB3_0/u_mux_p_to_b3/N_584 ));
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_data_out8_37  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_2_[6]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_642 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_37_net_1 ));
    INV_BA AFLSDF_INV_58 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_10_net_1 ), .Y(
        AFLSDF_INV_58_net_1));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_6_[7]  (.D(
        \CoreAPB3_0_APBmslave5_PWDATA[7] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB18_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_6__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_177_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_6_rs[7] ));
    SLE_IP_EN 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/FF_32  
        (.EN(VCC), .IPENn(AFLSDF_INV_145_net_1));
    IOOUTFF_BYPASS \GPIO_OUT_1_obuf[4]/U0/U_IOOUTFF  (.A(
        \GPIO_OUT_1_obuf[4]/U0/DOUT1 ), .Y(
        \GPIO_OUT_1_obuf[4]/U0/DOUT ));
    CFG2_IP_BC 
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/CFG_13  
        (.B(\CoreAPB3_0_APBmslave5_PWDATA[19] ), .C(
        \CoreAPB3_0_APBmslave5_PADDR[0] ), .IPB(
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/B_DIN_net[3] )
        , .IPC(
        \COREAPBLSRAM_0/genblk1.genblk1.lsram_512to35328x32_block0/block0/B_ADDR_net[5] )
        );
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_154_rs_RNI0MFV  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_13_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_154_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_1_rs[2] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_1_[2]_net_1 ));
    IOOUTFF_BYPASS \GPIO_OUT_1_obuf[7]/U0/U_IOOUTFF  (.A(
        \GPIO_OUT_1_obuf[7]/U0/DOUT1 ), .Y(
        \GPIO_OUT_1_obuf[7]/U0/DOUT ));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_44  (.A(
        GND), .B(VCC), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[27] ), .IPB(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_FM0_READY_net ), .IPC());
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_207  (
        .A(VCC), .B(GND), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[25] ), 
        .IPB(\hello_regs_MSS_0/MSS_ADLIB_INST/F_AWLEN_HBURST0_net[3] ), 
        .IPC());
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_180  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/MGPIO22B_F2H_GPIN_net ), .IPB(
        ), .IPC());
    CFG4 #( .INIT(16'h7350) )  
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_1[7]  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_15_[7]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/mem_14_[7]_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/N_654 ), .D(
        \reg_apb_wrp_0/reg16x8_0/N_650 ), .Y(
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_1[7]_net_1 ));
    GB \FCCC_0/GL1_INST  (.An(AFLSDF_INV_146_net_1), .ENn(GND), .YNn(
        \FCCC_0/GL1_INST/U0_YNn ), .YSn(
        \FCCC_0/GL1_INST/U0_YNn_GSouth ));
    CFG3 #( .INIT(8'hF2) )  
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_149  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_0_[5]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_645 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_149_i ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_163_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_31_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_163_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_163_rs_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_data_out8_25_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB6_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_2__1_sqmuxa ), .ALn(
        AFLSDF_INV_147_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(\reg_apb_wrp_0/reg16x8_0/un1_data_out8_25_set_net_1 ));
    IP_INTERFACE \hello_regs_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_231  (
        .A(VCC), .B(VCC), .C(VCC), .IPA(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[29] ), 
        .IPB(
        \hello_regs_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[41] ), 
        .IPC());
    INV_BA AFLSDF_INV_14 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_2_net_1 ), .Y(
        AFLSDF_INV_14_net_1));
    CFG4 #( .INIT(16'h7350) )  
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_0_1[6]  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_15_[6]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/mem_14_[6]_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/N_654 ), .D(
        \reg_apb_wrp_0/reg16x8_0/N_650 ), .Y(
        \reg_apb_wrp_0/reg16x8_0/data_out_2_15_i_0_1[6]_net_1 ));
    CFG4 #( .INIT(16'hECA0) )  \CoreAPB3_0/u_mux_p_to_b3/PRDATA_0[11]  
        (.A(\CoreAPB3_0/u_mux_p_to_b3/N_636 ), .B(
        \COREAPBLSRAM_0.PRDATA4 ), .C(\COREAPBLSRAM_0.PRDATA_reg[11] ), 
        .D(\COREAPBLSRAM_0.lsram_width32_PRDATA[11] ), .Y(
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[11] ));
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_data_out8_53  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_3_[6]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_655 ), .C(
        \hello_regs_MSS_0/FPGA_RESET_N ), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_data_out8_53_net_1 ));
    CFG4 #( .INIT(16'hECA0) )  \CoreAPB3_0/u_mux_p_to_b3/PRDATA_0[30]  
        (.A(\CoreAPB3_0/u_mux_p_to_b3/N_636 ), .B(
        \COREAPBLSRAM_0.PRDATA4 ), .C(\COREAPBLSRAM_0.PRDATA_reg[30] ), 
        .D(\COREAPBLSRAM_0.lsram_width32_PRDATA[30] ), .Y(
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[30] ));
    GND GND_power_inst1 (.Y(GND_power_net1));
    VCC VCC_power_inst1 (.Y(VCC_power_net1));
    
endmodule
