`timescale 1 ns/100 ps
// Version: v11.5 SP3 11.5.3.10


module RCOSC_25_50MHZ(
       CLKOUT
    );
output CLKOUT;

    parameter FREQUENCY = 50.0 ;
    
endmodule


module MSS_010(
       CAN_RXBUS_MGPIO3A_H2F_A,
       CAN_RXBUS_MGPIO3A_H2F_B,
       CAN_TX_EBL_MGPIO4A_H2F_A,
       CAN_TX_EBL_MGPIO4A_H2F_B,
       CAN_TXBUS_MGPIO2A_H2F_A,
       CAN_TXBUS_MGPIO2A_H2F_B,
       CLK_CONFIG_APB,
       COMMS_INT,
       CONFIG_PRESET_N,
       EDAC_ERROR,
       F_FM0_RDATA,
       F_FM0_READYOUT,
       F_FM0_RESP,
       F_HM0_ADDR,
       F_HM0_ENABLE,
       F_HM0_SEL,
       F_HM0_SIZE,
       F_HM0_TRANS1,
       F_HM0_WDATA,
       F_HM0_WRITE,
       FAB_CHRGVBUS,
       FAB_DISCHRGVBUS,
       FAB_DMPULLDOWN,
       FAB_DPPULLDOWN,
       FAB_DRVVBUS,
       FAB_IDPULLUP,
       FAB_OPMODE,
       FAB_SUSPENDM,
       FAB_TERMSEL,
       FAB_TXVALID,
       FAB_VCONTROL,
       FAB_VCONTROLLOADM,
       FAB_XCVRSEL,
       FAB_XDATAOUT,
       FACC_GLMUX_SEL,
       FIC32_0_MASTER,
       FIC32_1_MASTER,
       FPGA_RESET_N,
       GTX_CLK,
       H2F_INTERRUPT,
       H2F_NMI,
       H2FCALIB,
       I2C0_SCL_MGPIO31B_H2F_A,
       I2C0_SCL_MGPIO31B_H2F_B,
       I2C0_SDA_MGPIO30B_H2F_A,
       I2C0_SDA_MGPIO30B_H2F_B,
       I2C1_SCL_MGPIO1A_H2F_A,
       I2C1_SCL_MGPIO1A_H2F_B,
       I2C1_SDA_MGPIO0A_H2F_A,
       I2C1_SDA_MGPIO0A_H2F_B,
       MDCF,
       MDOENF,
       MDOF,
       MMUART0_CTS_MGPIO19B_H2F_A,
       MMUART0_CTS_MGPIO19B_H2F_B,
       MMUART0_DCD_MGPIO22B_H2F_A,
       MMUART0_DCD_MGPIO22B_H2F_B,
       MMUART0_DSR_MGPIO20B_H2F_A,
       MMUART0_DSR_MGPIO20B_H2F_B,
       MMUART0_DTR_MGPIO18B_H2F_A,
       MMUART0_DTR_MGPIO18B_H2F_B,
       MMUART0_RI_MGPIO21B_H2F_A,
       MMUART0_RI_MGPIO21B_H2F_B,
       MMUART0_RTS_MGPIO17B_H2F_A,
       MMUART0_RTS_MGPIO17B_H2F_B,
       MMUART0_RXD_MGPIO28B_H2F_A,
       MMUART0_RXD_MGPIO28B_H2F_B,
       MMUART0_SCK_MGPIO29B_H2F_A,
       MMUART0_SCK_MGPIO29B_H2F_B,
       MMUART0_TXD_MGPIO27B_H2F_A,
       MMUART0_TXD_MGPIO27B_H2F_B,
       MMUART1_DTR_MGPIO12B_H2F_A,
       MMUART1_RTS_MGPIO11B_H2F_A,
       MMUART1_RTS_MGPIO11B_H2F_B,
       MMUART1_RXD_MGPIO26B_H2F_A,
       MMUART1_RXD_MGPIO26B_H2F_B,
       MMUART1_SCK_MGPIO25B_H2F_A,
       MMUART1_SCK_MGPIO25B_H2F_B,
       MMUART1_TXD_MGPIO24B_H2F_A,
       MMUART1_TXD_MGPIO24B_H2F_B,
       MPLL_LOCK,
       PER2_FABRIC_PADDR,
       PER2_FABRIC_PENABLE,
       PER2_FABRIC_PSEL,
       PER2_FABRIC_PWDATA,
       PER2_FABRIC_PWRITE,
       RTC_MATCH,
       SLEEPDEEP,
       SLEEPHOLDACK,
       SLEEPING,
       SMBALERT_NO0,
       SMBALERT_NO1,
       SMBSUS_NO0,
       SMBSUS_NO1,
       SPI0_CLK_OUT,
       SPI0_SDI_MGPIO5A_H2F_A,
       SPI0_SDI_MGPIO5A_H2F_B,
       SPI0_SDO_MGPIO6A_H2F_A,
       SPI0_SDO_MGPIO6A_H2F_B,
       SPI0_SS0_MGPIO7A_H2F_A,
       SPI0_SS0_MGPIO7A_H2F_B,
       SPI0_SS1_MGPIO8A_H2F_A,
       SPI0_SS1_MGPIO8A_H2F_B,
       SPI0_SS2_MGPIO9A_H2F_A,
       SPI0_SS2_MGPIO9A_H2F_B,
       SPI0_SS3_MGPIO10A_H2F_A,
       SPI0_SS3_MGPIO10A_H2F_B,
       SPI0_SS4_MGPIO19A_H2F_A,
       SPI0_SS5_MGPIO20A_H2F_A,
       SPI0_SS6_MGPIO21A_H2F_A,
       SPI0_SS7_MGPIO22A_H2F_A,
       SPI1_CLK_OUT,
       SPI1_SDI_MGPIO11A_H2F_A,
       SPI1_SDI_MGPIO11A_H2F_B,
       SPI1_SDO_MGPIO12A_H2F_A,
       SPI1_SDO_MGPIO12A_H2F_B,
       SPI1_SS0_MGPIO13A_H2F_A,
       SPI1_SS0_MGPIO13A_H2F_B,
       SPI1_SS1_MGPIO14A_H2F_A,
       SPI1_SS1_MGPIO14A_H2F_B,
       SPI1_SS2_MGPIO15A_H2F_A,
       SPI1_SS2_MGPIO15A_H2F_B,
       SPI1_SS3_MGPIO16A_H2F_A,
       SPI1_SS3_MGPIO16A_H2F_B,
       SPI1_SS4_MGPIO17A_H2F_A,
       SPI1_SS5_MGPIO18A_H2F_A,
       SPI1_SS6_MGPIO23A_H2F_A,
       SPI1_SS7_MGPIO24A_H2F_A,
       TCGF,
       TRACECLK,
       TRACEDATA,
       TX_CLK,
       TX_ENF,
       TX_ERRF,
       TXCTL_EN_RIF,
       TXD_RIF,
       TXDF,
       TXEV,
       WDOGTIMEOUT,
       F_ARREADY_HREADYOUT1,
       F_AWREADY_HREADYOUT0,
       F_BID,
       F_BRESP_HRESP0,
       F_BVALID,
       F_RDATA_HRDATA01,
       F_RID,
       F_RLAST,
       F_RRESP_HRESP1,
       F_RVALID,
       F_WREADY,
       MDDR_FABRIC_PRDATA,
       MDDR_FABRIC_PREADY,
       MDDR_FABRIC_PSLVERR,
       CAN_RXBUS_F2H_SCP,
       CAN_TX_EBL_F2H_SCP,
       CAN_TXBUS_F2H_SCP,
       COLF,
       CRSF,
       F2_DMAREADY,
       F2H_INTERRUPT,
       F2HCALIB,
       F_DMAREADY,
       F_FM0_ADDR,
       F_FM0_ENABLE,
       F_FM0_MASTLOCK,
       F_FM0_READY,
       F_FM0_SEL,
       F_FM0_SIZE,
       F_FM0_TRANS1,
       F_FM0_WDATA,
       F_FM0_WRITE,
       F_HM0_RDATA,
       F_HM0_READY,
       F_HM0_RESP,
       FAB_AVALID,
       FAB_HOSTDISCON,
       FAB_IDDIG,
       FAB_LINESTATE,
       FAB_M3_RESET_N,
       FAB_PLL_LOCK,
       FAB_RXACTIVE,
       FAB_RXERROR,
       FAB_RXVALID,
       FAB_RXVALIDH,
       FAB_SESSEND,
       FAB_TXREADY,
       FAB_VBUSVALID,
       FAB_VSTATUS,
       FAB_XDATAIN,
       GTX_CLKPF,
       I2C0_BCLK,
       I2C0_SCL_F2H_SCP,
       I2C0_SDA_F2H_SCP,
       I2C1_BCLK,
       I2C1_SCL_F2H_SCP,
       I2C1_SDA_F2H_SCP,
       MDIF,
       MGPIO0A_F2H_GPIN,
       MGPIO10A_F2H_GPIN,
       MGPIO11A_F2H_GPIN,
       MGPIO11B_F2H_GPIN,
       MGPIO12A_F2H_GPIN,
       MGPIO13A_F2H_GPIN,
       MGPIO14A_F2H_GPIN,
       MGPIO15A_F2H_GPIN,
       MGPIO16A_F2H_GPIN,
       MGPIO17B_F2H_GPIN,
       MGPIO18B_F2H_GPIN,
       MGPIO19B_F2H_GPIN,
       MGPIO1A_F2H_GPIN,
       MGPIO20B_F2H_GPIN,
       MGPIO21B_F2H_GPIN,
       MGPIO22B_F2H_GPIN,
       MGPIO24B_F2H_GPIN,
       MGPIO25B_F2H_GPIN,
       MGPIO26B_F2H_GPIN,
       MGPIO27B_F2H_GPIN,
       MGPIO28B_F2H_GPIN,
       MGPIO29B_F2H_GPIN,
       MGPIO2A_F2H_GPIN,
       MGPIO30B_F2H_GPIN,
       MGPIO31B_F2H_GPIN,
       MGPIO3A_F2H_GPIN,
       MGPIO4A_F2H_GPIN,
       MGPIO5A_F2H_GPIN,
       MGPIO6A_F2H_GPIN,
       MGPIO7A_F2H_GPIN,
       MGPIO8A_F2H_GPIN,
       MGPIO9A_F2H_GPIN,
       MMUART0_CTS_F2H_SCP,
       MMUART0_DCD_F2H_SCP,
       MMUART0_DSR_F2H_SCP,
       MMUART0_DTR_F2H_SCP,
       MMUART0_RI_F2H_SCP,
       MMUART0_RTS_F2H_SCP,
       MMUART0_RXD_F2H_SCP,
       MMUART0_SCK_F2H_SCP,
       MMUART0_TXD_F2H_SCP,
       MMUART1_CTS_F2H_SCP,
       MMUART1_DCD_F2H_SCP,
       MMUART1_DSR_F2H_SCP,
       MMUART1_RI_F2H_SCP,
       MMUART1_RTS_F2H_SCP,
       MMUART1_RXD_F2H_SCP,
       MMUART1_SCK_F2H_SCP,
       MMUART1_TXD_F2H_SCP,
       PER2_FABRIC_PRDATA,
       PER2_FABRIC_PREADY,
       PER2_FABRIC_PSLVERR,
       RCGF,
       RX_CLKPF,
       RX_DVF,
       RX_ERRF,
       RX_EV,
       RXDF,
       SLEEPHOLDREQ,
       SMBALERT_NI0,
       SMBALERT_NI1,
       SMBSUS_NI0,
       SMBSUS_NI1,
       SPI0_CLK_IN,
       SPI0_SDI_F2H_SCP,
       SPI0_SDO_F2H_SCP,
       SPI0_SS0_F2H_SCP,
       SPI0_SS1_F2H_SCP,
       SPI0_SS2_F2H_SCP,
       SPI0_SS3_F2H_SCP,
       SPI1_CLK_IN,
       SPI1_SDI_F2H_SCP,
       SPI1_SDO_F2H_SCP,
       SPI1_SS0_F2H_SCP,
       SPI1_SS1_F2H_SCP,
       SPI1_SS2_F2H_SCP,
       SPI1_SS3_F2H_SCP,
       TX_CLKPF,
       USER_MSS_GPIO_RESET_N,
       USER_MSS_RESET_N,
       XCLK_FAB,
       CLK_BASE,
       CLK_MDDR_APB,
       F_ARADDR_HADDR1,
       F_ARBURST_HTRANS1,
       F_ARID_HSEL1,
       F_ARLEN_HBURST1,
       F_ARLOCK_HMASTLOCK1,
       F_ARSIZE_HSIZE1,
       F_ARVALID_HWRITE1,
       F_AWADDR_HADDR0,
       F_AWBURST_HTRANS0,
       F_AWID_HSEL0,
       F_AWLEN_HBURST0,
       F_AWLOCK_HMASTLOCK0,
       F_AWSIZE_HSIZE0,
       F_AWVALID_HWRITE0,
       F_BREADY,
       F_RMW_AXI,
       F_RREADY,
       F_WDATA_HWDATA01,
       F_WID_HREADY01,
       F_WLAST,
       F_WSTRB,
       F_WVALID,
       FPGA_MDDR_ARESET_N,
       MDDR_FABRIC_PADDR,
       MDDR_FABRIC_PENABLE,
       MDDR_FABRIC_PSEL,
       MDDR_FABRIC_PWDATA,
       MDDR_FABRIC_PWRITE,
       PRESET_N,
       CAN_RXBUS_USBA_DATA1_MGPIO3A_IN,
       CAN_TX_EBL_USBA_DATA2_MGPIO4A_IN,
       CAN_TXBUS_USBA_DATA0_MGPIO2A_IN,
       DM_IN,
       DRAM_DQ_IN,
       DRAM_DQS_IN,
       DRAM_FIFO_WE_IN,
       I2C0_SCL_USBC_DATA1_MGPIO31B_IN,
       I2C0_SDA_USBC_DATA0_MGPIO30B_IN,
       I2C1_SCL_USBA_DATA4_MGPIO1A_IN,
       I2C1_SDA_USBA_DATA3_MGPIO0A_IN,
       MMUART0_CTS_USBC_DATA7_MGPIO19B_IN,
       MMUART0_DCD_MGPIO22B_IN,
       MMUART0_DSR_MGPIO20B_IN,
       MMUART0_DTR_USBC_DATA6_MGPIO18B_IN,
       MMUART0_RI_MGPIO21B_IN,
       MMUART0_RTS_USBC_DATA5_MGPIO17B_IN,
       MMUART0_RXD_USBC_STP_MGPIO28B_IN,
       MMUART0_SCK_USBC_NXT_MGPIO29B_IN,
       MMUART0_TXD_USBC_DIR_MGPIO27B_IN,
       MMUART1_RXD_USBC_DATA3_MGPIO26B_IN,
       MMUART1_SCK_USBC_DATA4_MGPIO25B_IN,
       MMUART1_TXD_USBC_DATA2_MGPIO24B_IN,
       RGMII_GTX_CLK_RMII_CLK_USBB_XCLK_IN,
       RGMII_MDC_RMII_MDC_IN,
       RGMII_MDIO_RMII_MDIO_USBB_DATA7_IN,
       RGMII_RX_CLK_IN,
       RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_IN,
       RGMII_RXD0_RMII_RXD0_USBB_DATA0_IN,
       RGMII_RXD1_RMII_RXD1_USBB_DATA1_IN,
       RGMII_RXD2_RMII_RX_ER_USBB_DATA3_IN,
       RGMII_RXD3_USBB_DATA4_IN,
       RGMII_TX_CLK_IN,
       RGMII_TX_CTL_RMII_TX_EN_USBB_NXT_IN,
       RGMII_TXD0_RMII_TXD0_USBB_DIR_IN,
       RGMII_TXD1_RMII_TXD1_USBB_STP_IN,
       RGMII_TXD2_USBB_DATA5_IN,
       RGMII_TXD3_USBB_DATA6_IN,
       SPI0_SCK_USBA_XCLK_IN,
       SPI0_SDI_USBA_DIR_MGPIO5A_IN,
       SPI0_SDO_USBA_STP_MGPIO6A_IN,
       SPI0_SS0_USBA_NXT_MGPIO7A_IN,
       SPI0_SS1_USBA_DATA5_MGPIO8A_IN,
       SPI0_SS2_USBA_DATA6_MGPIO9A_IN,
       SPI0_SS3_USBA_DATA7_MGPIO10A_IN,
       SPI1_SCK_IN,
       SPI1_SDI_MGPIO11A_IN,
       SPI1_SDO_MGPIO12A_IN,
       SPI1_SS0_MGPIO13A_IN,
       SPI1_SS1_MGPIO14A_IN,
       SPI1_SS2_MGPIO15A_IN,
       SPI1_SS3_MGPIO16A_IN,
       SPI1_SS4_MGPIO17A_IN,
       SPI1_SS5_MGPIO18A_IN,
       SPI1_SS6_MGPIO23A_IN,
       SPI1_SS7_MGPIO24A_IN,
       USBC_XCLK_IN,
       CAN_RXBUS_USBA_DATA1_MGPIO3A_OUT,
       CAN_TX_EBL_USBA_DATA2_MGPIO4A_OUT,
       CAN_TXBUS_USBA_DATA0_MGPIO2A_OUT,
       DRAM_ADDR,
       DRAM_BA,
       DRAM_CASN,
       DRAM_CKE,
       DRAM_CLK,
       DRAM_CSN,
       DRAM_DM_RDQS_OUT,
       DRAM_DQ_OUT,
       DRAM_DQS_OUT,
       DRAM_FIFO_WE_OUT,
       DRAM_ODT,
       DRAM_RASN,
       DRAM_RSTN,
       DRAM_WEN,
       I2C0_SCL_USBC_DATA1_MGPIO31B_OUT,
       I2C0_SDA_USBC_DATA0_MGPIO30B_OUT,
       I2C1_SCL_USBA_DATA4_MGPIO1A_OUT,
       I2C1_SDA_USBA_DATA3_MGPIO0A_OUT,
       MMUART0_CTS_USBC_DATA7_MGPIO19B_OUT,
       MMUART0_DCD_MGPIO22B_OUT,
       MMUART0_DSR_MGPIO20B_OUT,
       MMUART0_DTR_USBC_DATA6_MGPIO18B_OUT,
       MMUART0_RI_MGPIO21B_OUT,
       MMUART0_RTS_USBC_DATA5_MGPIO17B_OUT,
       MMUART0_RXD_USBC_STP_MGPIO28B_OUT,
       MMUART0_SCK_USBC_NXT_MGPIO29B_OUT,
       MMUART0_TXD_USBC_DIR_MGPIO27B_OUT,
       MMUART1_RXD_USBC_DATA3_MGPIO26B_OUT,
       MMUART1_SCK_USBC_DATA4_MGPIO25B_OUT,
       MMUART1_TXD_USBC_DATA2_MGPIO24B_OUT,
       RGMII_GTX_CLK_RMII_CLK_USBB_XCLK_OUT,
       RGMII_MDC_RMII_MDC_OUT,
       RGMII_MDIO_RMII_MDIO_USBB_DATA7_OUT,
       RGMII_RX_CLK_OUT,
       RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_OUT,
       RGMII_RXD0_RMII_RXD0_USBB_DATA0_OUT,
       RGMII_RXD1_RMII_RXD1_USBB_DATA1_OUT,
       RGMII_RXD2_RMII_RX_ER_USBB_DATA3_OUT,
       RGMII_RXD3_USBB_DATA4_OUT,
       RGMII_TX_CLK_OUT,
       RGMII_TX_CTL_RMII_TX_EN_USBB_NXT_OUT,
       RGMII_TXD0_RMII_TXD0_USBB_DIR_OUT,
       RGMII_TXD1_RMII_TXD1_USBB_STP_OUT,
       RGMII_TXD2_USBB_DATA5_OUT,
       RGMII_TXD3_USBB_DATA6_OUT,
       SPI0_SCK_USBA_XCLK_OUT,
       SPI0_SDI_USBA_DIR_MGPIO5A_OUT,
       SPI0_SDO_USBA_STP_MGPIO6A_OUT,
       SPI0_SS0_USBA_NXT_MGPIO7A_OUT,
       SPI0_SS1_USBA_DATA5_MGPIO8A_OUT,
       SPI0_SS2_USBA_DATA6_MGPIO9A_OUT,
       SPI0_SS3_USBA_DATA7_MGPIO10A_OUT,
       SPI1_SCK_OUT,
       SPI1_SDI_MGPIO11A_OUT,
       SPI1_SDO_MGPIO12A_OUT,
       SPI1_SS0_MGPIO13A_OUT,
       SPI1_SS1_MGPIO14A_OUT,
       SPI1_SS2_MGPIO15A_OUT,
       SPI1_SS3_MGPIO16A_OUT,
       SPI1_SS4_MGPIO17A_OUT,
       SPI1_SS5_MGPIO18A_OUT,
       SPI1_SS6_MGPIO23A_OUT,
       SPI1_SS7_MGPIO24A_OUT,
       USBC_XCLK_OUT,
       CAN_RXBUS_USBA_DATA1_MGPIO3A_OE,
       CAN_TX_EBL_USBA_DATA2_MGPIO4A_OE,
       CAN_TXBUS_USBA_DATA0_MGPIO2A_OE,
       DM_OE,
       DRAM_DQ_OE,
       DRAM_DQS_OE,
       I2C0_SCL_USBC_DATA1_MGPIO31B_OE,
       I2C0_SDA_USBC_DATA0_MGPIO30B_OE,
       I2C1_SCL_USBA_DATA4_MGPIO1A_OE,
       I2C1_SDA_USBA_DATA3_MGPIO0A_OE,
       MMUART0_CTS_USBC_DATA7_MGPIO19B_OE,
       MMUART0_DCD_MGPIO22B_OE,
       MMUART0_DSR_MGPIO20B_OE,
       MMUART0_DTR_USBC_DATA6_MGPIO18B_OE,
       MMUART0_RI_MGPIO21B_OE,
       MMUART0_RTS_USBC_DATA5_MGPIO17B_OE,
       MMUART0_RXD_USBC_STP_MGPIO28B_OE,
       MMUART0_SCK_USBC_NXT_MGPIO29B_OE,
       MMUART0_TXD_USBC_DIR_MGPIO27B_OE,
       MMUART1_RXD_USBC_DATA3_MGPIO26B_OE,
       MMUART1_SCK_USBC_DATA4_MGPIO25B_OE,
       MMUART1_TXD_USBC_DATA2_MGPIO24B_OE,
       RGMII_GTX_CLK_RMII_CLK_USBB_XCLK_OE,
       RGMII_MDC_RMII_MDC_OE,
       RGMII_MDIO_RMII_MDIO_USBB_DATA7_OE,
       RGMII_RX_CLK_OE,
       RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_OE,
       RGMII_RXD0_RMII_RXD0_USBB_DATA0_OE,
       RGMII_RXD1_RMII_RXD1_USBB_DATA1_OE,
       RGMII_RXD2_RMII_RX_ER_USBB_DATA3_OE,
       RGMII_RXD3_USBB_DATA4_OE,
       RGMII_TX_CLK_OE,
       RGMII_TX_CTL_RMII_TX_EN_USBB_NXT_OE,
       RGMII_TXD0_RMII_TXD0_USBB_DIR_OE,
       RGMII_TXD1_RMII_TXD1_USBB_STP_OE,
       RGMII_TXD2_USBB_DATA5_OE,
       RGMII_TXD3_USBB_DATA6_OE,
       SPI0_SCK_USBA_XCLK_OE,
       SPI0_SDI_USBA_DIR_MGPIO5A_OE,
       SPI0_SDO_USBA_STP_MGPIO6A_OE,
       SPI0_SS0_USBA_NXT_MGPIO7A_OE,
       SPI0_SS1_USBA_DATA5_MGPIO8A_OE,
       SPI0_SS2_USBA_DATA6_MGPIO9A_OE,
       SPI0_SS3_USBA_DATA7_MGPIO10A_OE,
       SPI1_SCK_OE,
       SPI1_SDI_MGPIO11A_OE,
       SPI1_SDO_MGPIO12A_OE,
       SPI1_SS0_MGPIO13A_OE,
       SPI1_SS1_MGPIO14A_OE,
       SPI1_SS2_MGPIO15A_OE,
       SPI1_SS3_MGPIO16A_OE,
       SPI1_SS4_MGPIO17A_OE,
       SPI1_SS5_MGPIO18A_OE,
       SPI1_SS6_MGPIO23A_OE,
       SPI1_SS7_MGPIO24A_OE,
       USBC_XCLK_OE
    );
output CAN_RXBUS_MGPIO3A_H2F_A;
output CAN_RXBUS_MGPIO3A_H2F_B;
output CAN_TX_EBL_MGPIO4A_H2F_A;
output CAN_TX_EBL_MGPIO4A_H2F_B;
output CAN_TXBUS_MGPIO2A_H2F_A;
output CAN_TXBUS_MGPIO2A_H2F_B;
output CLK_CONFIG_APB;
output COMMS_INT;
output CONFIG_PRESET_N;
output [7:0] EDAC_ERROR;
output [31:0] F_FM0_RDATA;
output F_FM0_READYOUT;
output F_FM0_RESP;
output [31:0] F_HM0_ADDR;
output F_HM0_ENABLE;
output F_HM0_SEL;
output [1:0] F_HM0_SIZE;
output F_HM0_TRANS1;
output [31:0] F_HM0_WDATA;
output F_HM0_WRITE;
output FAB_CHRGVBUS;
output FAB_DISCHRGVBUS;
output FAB_DMPULLDOWN;
output FAB_DPPULLDOWN;
output FAB_DRVVBUS;
output FAB_IDPULLUP;
output [1:0] FAB_OPMODE;
output FAB_SUSPENDM;
output FAB_TERMSEL;
output FAB_TXVALID;
output [3:0] FAB_VCONTROL;
output FAB_VCONTROLLOADM;
output [1:0] FAB_XCVRSEL;
output [7:0] FAB_XDATAOUT;
output FACC_GLMUX_SEL;
output [1:0] FIC32_0_MASTER;
output [1:0] FIC32_1_MASTER;
output FPGA_RESET_N;
output GTX_CLK;
output [15:0] H2F_INTERRUPT;
output H2F_NMI;
output H2FCALIB;
output I2C0_SCL_MGPIO31B_H2F_A;
output I2C0_SCL_MGPIO31B_H2F_B;
output I2C0_SDA_MGPIO30B_H2F_A;
output I2C0_SDA_MGPIO30B_H2F_B;
output I2C1_SCL_MGPIO1A_H2F_A;
output I2C1_SCL_MGPIO1A_H2F_B;
output I2C1_SDA_MGPIO0A_H2F_A;
output I2C1_SDA_MGPIO0A_H2F_B;
output MDCF;
output MDOENF;
output MDOF;
output MMUART0_CTS_MGPIO19B_H2F_A;
output MMUART0_CTS_MGPIO19B_H2F_B;
output MMUART0_DCD_MGPIO22B_H2F_A;
output MMUART0_DCD_MGPIO22B_H2F_B;
output MMUART0_DSR_MGPIO20B_H2F_A;
output MMUART0_DSR_MGPIO20B_H2F_B;
output MMUART0_DTR_MGPIO18B_H2F_A;
output MMUART0_DTR_MGPIO18B_H2F_B;
output MMUART0_RI_MGPIO21B_H2F_A;
output MMUART0_RI_MGPIO21B_H2F_B;
output MMUART0_RTS_MGPIO17B_H2F_A;
output MMUART0_RTS_MGPIO17B_H2F_B;
output MMUART0_RXD_MGPIO28B_H2F_A;
output MMUART0_RXD_MGPIO28B_H2F_B;
output MMUART0_SCK_MGPIO29B_H2F_A;
output MMUART0_SCK_MGPIO29B_H2F_B;
output MMUART0_TXD_MGPIO27B_H2F_A;
output MMUART0_TXD_MGPIO27B_H2F_B;
output MMUART1_DTR_MGPIO12B_H2F_A;
output MMUART1_RTS_MGPIO11B_H2F_A;
output MMUART1_RTS_MGPIO11B_H2F_B;
output MMUART1_RXD_MGPIO26B_H2F_A;
output MMUART1_RXD_MGPIO26B_H2F_B;
output MMUART1_SCK_MGPIO25B_H2F_A;
output MMUART1_SCK_MGPIO25B_H2F_B;
output MMUART1_TXD_MGPIO24B_H2F_A;
output MMUART1_TXD_MGPIO24B_H2F_B;
output MPLL_LOCK;
output [15:2] PER2_FABRIC_PADDR;
output PER2_FABRIC_PENABLE;
output PER2_FABRIC_PSEL;
output [31:0] PER2_FABRIC_PWDATA;
output PER2_FABRIC_PWRITE;
output RTC_MATCH;
output SLEEPDEEP;
output SLEEPHOLDACK;
output SLEEPING;
output SMBALERT_NO0;
output SMBALERT_NO1;
output SMBSUS_NO0;
output SMBSUS_NO1;
output SPI0_CLK_OUT;
output SPI0_SDI_MGPIO5A_H2F_A;
output SPI0_SDI_MGPIO5A_H2F_B;
output SPI0_SDO_MGPIO6A_H2F_A;
output SPI0_SDO_MGPIO6A_H2F_B;
output SPI0_SS0_MGPIO7A_H2F_A;
output SPI0_SS0_MGPIO7A_H2F_B;
output SPI0_SS1_MGPIO8A_H2F_A;
output SPI0_SS1_MGPIO8A_H2F_B;
output SPI0_SS2_MGPIO9A_H2F_A;
output SPI0_SS2_MGPIO9A_H2F_B;
output SPI0_SS3_MGPIO10A_H2F_A;
output SPI0_SS3_MGPIO10A_H2F_B;
output SPI0_SS4_MGPIO19A_H2F_A;
output SPI0_SS5_MGPIO20A_H2F_A;
output SPI0_SS6_MGPIO21A_H2F_A;
output SPI0_SS7_MGPIO22A_H2F_A;
output SPI1_CLK_OUT;
output SPI1_SDI_MGPIO11A_H2F_A;
output SPI1_SDI_MGPIO11A_H2F_B;
output SPI1_SDO_MGPIO12A_H2F_A;
output SPI1_SDO_MGPIO12A_H2F_B;
output SPI1_SS0_MGPIO13A_H2F_A;
output SPI1_SS0_MGPIO13A_H2F_B;
output SPI1_SS1_MGPIO14A_H2F_A;
output SPI1_SS1_MGPIO14A_H2F_B;
output SPI1_SS2_MGPIO15A_H2F_A;
output SPI1_SS2_MGPIO15A_H2F_B;
output SPI1_SS3_MGPIO16A_H2F_A;
output SPI1_SS3_MGPIO16A_H2F_B;
output SPI1_SS4_MGPIO17A_H2F_A;
output SPI1_SS5_MGPIO18A_H2F_A;
output SPI1_SS6_MGPIO23A_H2F_A;
output SPI1_SS7_MGPIO24A_H2F_A;
output [9:0] TCGF;
output TRACECLK;
output [3:0] TRACEDATA;
output TX_CLK;
output TX_ENF;
output TX_ERRF;
output TXCTL_EN_RIF;
output [3:0] TXD_RIF;
output [7:0] TXDF;
output TXEV;
output WDOGTIMEOUT;
output F_ARREADY_HREADYOUT1;
output F_AWREADY_HREADYOUT0;
output [3:0] F_BID;
output [1:0] F_BRESP_HRESP0;
output F_BVALID;
output [63:0] F_RDATA_HRDATA01;
output [3:0] F_RID;
output F_RLAST;
output [1:0] F_RRESP_HRESP1;
output F_RVALID;
output F_WREADY;
output [15:0] MDDR_FABRIC_PRDATA;
output MDDR_FABRIC_PREADY;
output MDDR_FABRIC_PSLVERR;
input  CAN_RXBUS_F2H_SCP;
input  CAN_TX_EBL_F2H_SCP;
input  CAN_TXBUS_F2H_SCP;
input  COLF;
input  CRSF;
input  [1:0] F2_DMAREADY;
input  [15:0] F2H_INTERRUPT;
input  F2HCALIB;
input  [1:0] F_DMAREADY;
input  [31:0] F_FM0_ADDR;
input  F_FM0_ENABLE;
input  F_FM0_MASTLOCK;
input  F_FM0_READY;
input  F_FM0_SEL;
input  [1:0] F_FM0_SIZE;
input  F_FM0_TRANS1;
input  [31:0] F_FM0_WDATA;
input  F_FM0_WRITE;
input  [31:0] F_HM0_RDATA;
input  F_HM0_READY;
input  F_HM0_RESP;
input  FAB_AVALID;
input  FAB_HOSTDISCON;
input  FAB_IDDIG;
input  [1:0] FAB_LINESTATE;
input  FAB_M3_RESET_N;
input  FAB_PLL_LOCK;
input  FAB_RXACTIVE;
input  FAB_RXERROR;
input  FAB_RXVALID;
input  FAB_RXVALIDH;
input  FAB_SESSEND;
input  FAB_TXREADY;
input  FAB_VBUSVALID;
input  [7:0] FAB_VSTATUS;
input  [7:0] FAB_XDATAIN;
input  GTX_CLKPF;
input  I2C0_BCLK;
input  I2C0_SCL_F2H_SCP;
input  I2C0_SDA_F2H_SCP;
input  I2C1_BCLK;
input  I2C1_SCL_F2H_SCP;
input  I2C1_SDA_F2H_SCP;
input  MDIF;
input  MGPIO0A_F2H_GPIN;
input  MGPIO10A_F2H_GPIN;
input  MGPIO11A_F2H_GPIN;
input  MGPIO11B_F2H_GPIN;
input  MGPIO12A_F2H_GPIN;
input  MGPIO13A_F2H_GPIN;
input  MGPIO14A_F2H_GPIN;
input  MGPIO15A_F2H_GPIN;
input  MGPIO16A_F2H_GPIN;
input  MGPIO17B_F2H_GPIN;
input  MGPIO18B_F2H_GPIN;
input  MGPIO19B_F2H_GPIN;
input  MGPIO1A_F2H_GPIN;
input  MGPIO20B_F2H_GPIN;
input  MGPIO21B_F2H_GPIN;
input  MGPIO22B_F2H_GPIN;
input  MGPIO24B_F2H_GPIN;
input  MGPIO25B_F2H_GPIN;
input  MGPIO26B_F2H_GPIN;
input  MGPIO27B_F2H_GPIN;
input  MGPIO28B_F2H_GPIN;
input  MGPIO29B_F2H_GPIN;
input  MGPIO2A_F2H_GPIN;
input  MGPIO30B_F2H_GPIN;
input  MGPIO31B_F2H_GPIN;
input  MGPIO3A_F2H_GPIN;
input  MGPIO4A_F2H_GPIN;
input  MGPIO5A_F2H_GPIN;
input  MGPIO6A_F2H_GPIN;
input  MGPIO7A_F2H_GPIN;
input  MGPIO8A_F2H_GPIN;
input  MGPIO9A_F2H_GPIN;
input  MMUART0_CTS_F2H_SCP;
input  MMUART0_DCD_F2H_SCP;
input  MMUART0_DSR_F2H_SCP;
input  MMUART0_DTR_F2H_SCP;
input  MMUART0_RI_F2H_SCP;
input  MMUART0_RTS_F2H_SCP;
input  MMUART0_RXD_F2H_SCP;
input  MMUART0_SCK_F2H_SCP;
input  MMUART0_TXD_F2H_SCP;
input  MMUART1_CTS_F2H_SCP;
input  MMUART1_DCD_F2H_SCP;
input  MMUART1_DSR_F2H_SCP;
input  MMUART1_RI_F2H_SCP;
input  MMUART1_RTS_F2H_SCP;
input  MMUART1_RXD_F2H_SCP;
input  MMUART1_SCK_F2H_SCP;
input  MMUART1_TXD_F2H_SCP;
input  [31:0] PER2_FABRIC_PRDATA;
input  PER2_FABRIC_PREADY;
input  PER2_FABRIC_PSLVERR;
input  [9:0] RCGF;
input  RX_CLKPF;
input  RX_DVF;
input  RX_ERRF;
input  RX_EV;
input  [7:0] RXDF;
input  SLEEPHOLDREQ;
input  SMBALERT_NI0;
input  SMBALERT_NI1;
input  SMBSUS_NI0;
input  SMBSUS_NI1;
input  SPI0_CLK_IN;
input  SPI0_SDI_F2H_SCP;
input  SPI0_SDO_F2H_SCP;
input  SPI0_SS0_F2H_SCP;
input  SPI0_SS1_F2H_SCP;
input  SPI0_SS2_F2H_SCP;
input  SPI0_SS3_F2H_SCP;
input  SPI1_CLK_IN;
input  SPI1_SDI_F2H_SCP;
input  SPI1_SDO_F2H_SCP;
input  SPI1_SS0_F2H_SCP;
input  SPI1_SS1_F2H_SCP;
input  SPI1_SS2_F2H_SCP;
input  SPI1_SS3_F2H_SCP;
input  TX_CLKPF;
input  USER_MSS_GPIO_RESET_N;
input  USER_MSS_RESET_N;
input  XCLK_FAB;
input  CLK_BASE;
input  CLK_MDDR_APB;
input  [31:0] F_ARADDR_HADDR1;
input  [1:0] F_ARBURST_HTRANS1;
input  [3:0] F_ARID_HSEL1;
input  [3:0] F_ARLEN_HBURST1;
input  [1:0] F_ARLOCK_HMASTLOCK1;
input  [1:0] F_ARSIZE_HSIZE1;
input  F_ARVALID_HWRITE1;
input  [31:0] F_AWADDR_HADDR0;
input  [1:0] F_AWBURST_HTRANS0;
input  [3:0] F_AWID_HSEL0;
input  [3:0] F_AWLEN_HBURST0;
input  [1:0] F_AWLOCK_HMASTLOCK0;
input  [1:0] F_AWSIZE_HSIZE0;
input  F_AWVALID_HWRITE0;
input  F_BREADY;
input  F_RMW_AXI;
input  F_RREADY;
input  [63:0] F_WDATA_HWDATA01;
input  [3:0] F_WID_HREADY01;
input  F_WLAST;
input  [7:0] F_WSTRB;
input  F_WVALID;
input  FPGA_MDDR_ARESET_N;
input  [10:2] MDDR_FABRIC_PADDR;
input  MDDR_FABRIC_PENABLE;
input  MDDR_FABRIC_PSEL;
input  [15:0] MDDR_FABRIC_PWDATA;
input  MDDR_FABRIC_PWRITE;
input  PRESET_N;
input  CAN_RXBUS_USBA_DATA1_MGPIO3A_IN;
input  CAN_TX_EBL_USBA_DATA2_MGPIO4A_IN;
input  CAN_TXBUS_USBA_DATA0_MGPIO2A_IN;
input  [2:0] DM_IN;
input  [17:0] DRAM_DQ_IN;
input  [2:0] DRAM_DQS_IN;
input  [1:0] DRAM_FIFO_WE_IN;
input  I2C0_SCL_USBC_DATA1_MGPIO31B_IN;
input  I2C0_SDA_USBC_DATA0_MGPIO30B_IN;
input  I2C1_SCL_USBA_DATA4_MGPIO1A_IN;
input  I2C1_SDA_USBA_DATA3_MGPIO0A_IN;
input  MMUART0_CTS_USBC_DATA7_MGPIO19B_IN;
input  MMUART0_DCD_MGPIO22B_IN;
input  MMUART0_DSR_MGPIO20B_IN;
input  MMUART0_DTR_USBC_DATA6_MGPIO18B_IN;
input  MMUART0_RI_MGPIO21B_IN;
input  MMUART0_RTS_USBC_DATA5_MGPIO17B_IN;
input  MMUART0_RXD_USBC_STP_MGPIO28B_IN;
input  MMUART0_SCK_USBC_NXT_MGPIO29B_IN;
input  MMUART0_TXD_USBC_DIR_MGPIO27B_IN;
input  MMUART1_RXD_USBC_DATA3_MGPIO26B_IN;
input  MMUART1_SCK_USBC_DATA4_MGPIO25B_IN;
input  MMUART1_TXD_USBC_DATA2_MGPIO24B_IN;
input  RGMII_GTX_CLK_RMII_CLK_USBB_XCLK_IN;
input  RGMII_MDC_RMII_MDC_IN;
input  RGMII_MDIO_RMII_MDIO_USBB_DATA7_IN;
input  RGMII_RX_CLK_IN;
input  RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_IN;
input  RGMII_RXD0_RMII_RXD0_USBB_DATA0_IN;
input  RGMII_RXD1_RMII_RXD1_USBB_DATA1_IN;
input  RGMII_RXD2_RMII_RX_ER_USBB_DATA3_IN;
input  RGMII_RXD3_USBB_DATA4_IN;
input  RGMII_TX_CLK_IN;
input  RGMII_TX_CTL_RMII_TX_EN_USBB_NXT_IN;
input  RGMII_TXD0_RMII_TXD0_USBB_DIR_IN;
input  RGMII_TXD1_RMII_TXD1_USBB_STP_IN;
input  RGMII_TXD2_USBB_DATA5_IN;
input  RGMII_TXD3_USBB_DATA6_IN;
input  SPI0_SCK_USBA_XCLK_IN;
input  SPI0_SDI_USBA_DIR_MGPIO5A_IN;
input  SPI0_SDO_USBA_STP_MGPIO6A_IN;
input  SPI0_SS0_USBA_NXT_MGPIO7A_IN;
input  SPI0_SS1_USBA_DATA5_MGPIO8A_IN;
input  SPI0_SS2_USBA_DATA6_MGPIO9A_IN;
input  SPI0_SS3_USBA_DATA7_MGPIO10A_IN;
input  SPI1_SCK_IN;
input  SPI1_SDI_MGPIO11A_IN;
input  SPI1_SDO_MGPIO12A_IN;
input  SPI1_SS0_MGPIO13A_IN;
input  SPI1_SS1_MGPIO14A_IN;
input  SPI1_SS2_MGPIO15A_IN;
input  SPI1_SS3_MGPIO16A_IN;
input  SPI1_SS4_MGPIO17A_IN;
input  SPI1_SS5_MGPIO18A_IN;
input  SPI1_SS6_MGPIO23A_IN;
input  SPI1_SS7_MGPIO24A_IN;
input  USBC_XCLK_IN;
output CAN_RXBUS_USBA_DATA1_MGPIO3A_OUT;
output CAN_TX_EBL_USBA_DATA2_MGPIO4A_OUT;
output CAN_TXBUS_USBA_DATA0_MGPIO2A_OUT;
output [15:0] DRAM_ADDR;
output [2:0] DRAM_BA;
output DRAM_CASN;
output DRAM_CKE;
output DRAM_CLK;
output DRAM_CSN;
output [2:0] DRAM_DM_RDQS_OUT;
output [17:0] DRAM_DQ_OUT;
output [2:0] DRAM_DQS_OUT;
output [1:0] DRAM_FIFO_WE_OUT;
output DRAM_ODT;
output DRAM_RASN;
output DRAM_RSTN;
output DRAM_WEN;
output I2C0_SCL_USBC_DATA1_MGPIO31B_OUT;
output I2C0_SDA_USBC_DATA0_MGPIO30B_OUT;
output I2C1_SCL_USBA_DATA4_MGPIO1A_OUT;
output I2C1_SDA_USBA_DATA3_MGPIO0A_OUT;
output MMUART0_CTS_USBC_DATA7_MGPIO19B_OUT;
output MMUART0_DCD_MGPIO22B_OUT;
output MMUART0_DSR_MGPIO20B_OUT;
output MMUART0_DTR_USBC_DATA6_MGPIO18B_OUT;
output MMUART0_RI_MGPIO21B_OUT;
output MMUART0_RTS_USBC_DATA5_MGPIO17B_OUT;
output MMUART0_RXD_USBC_STP_MGPIO28B_OUT;
output MMUART0_SCK_USBC_NXT_MGPIO29B_OUT;
output MMUART0_TXD_USBC_DIR_MGPIO27B_OUT;
output MMUART1_RXD_USBC_DATA3_MGPIO26B_OUT;
output MMUART1_SCK_USBC_DATA4_MGPIO25B_OUT;
output MMUART1_TXD_USBC_DATA2_MGPIO24B_OUT;
output RGMII_GTX_CLK_RMII_CLK_USBB_XCLK_OUT;
output RGMII_MDC_RMII_MDC_OUT;
output RGMII_MDIO_RMII_MDIO_USBB_DATA7_OUT;
output RGMII_RX_CLK_OUT;
output RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_OUT;
output RGMII_RXD0_RMII_RXD0_USBB_DATA0_OUT;
output RGMII_RXD1_RMII_RXD1_USBB_DATA1_OUT;
output RGMII_RXD2_RMII_RX_ER_USBB_DATA3_OUT;
output RGMII_RXD3_USBB_DATA4_OUT;
output RGMII_TX_CLK_OUT;
output RGMII_TX_CTL_RMII_TX_EN_USBB_NXT_OUT;
output RGMII_TXD0_RMII_TXD0_USBB_DIR_OUT;
output RGMII_TXD1_RMII_TXD1_USBB_STP_OUT;
output RGMII_TXD2_USBB_DATA5_OUT;
output RGMII_TXD3_USBB_DATA6_OUT;
output SPI0_SCK_USBA_XCLK_OUT;
output SPI0_SDI_USBA_DIR_MGPIO5A_OUT;
output SPI0_SDO_USBA_STP_MGPIO6A_OUT;
output SPI0_SS0_USBA_NXT_MGPIO7A_OUT;
output SPI0_SS1_USBA_DATA5_MGPIO8A_OUT;
output SPI0_SS2_USBA_DATA6_MGPIO9A_OUT;
output SPI0_SS3_USBA_DATA7_MGPIO10A_OUT;
output SPI1_SCK_OUT;
output SPI1_SDI_MGPIO11A_OUT;
output SPI1_SDO_MGPIO12A_OUT;
output SPI1_SS0_MGPIO13A_OUT;
output SPI1_SS1_MGPIO14A_OUT;
output SPI1_SS2_MGPIO15A_OUT;
output SPI1_SS3_MGPIO16A_OUT;
output SPI1_SS4_MGPIO17A_OUT;
output SPI1_SS5_MGPIO18A_OUT;
output SPI1_SS6_MGPIO23A_OUT;
output SPI1_SS7_MGPIO24A_OUT;
output USBC_XCLK_OUT;
output CAN_RXBUS_USBA_DATA1_MGPIO3A_OE;
output CAN_TX_EBL_USBA_DATA2_MGPIO4A_OE;
output CAN_TXBUS_USBA_DATA0_MGPIO2A_OE;
output [2:0] DM_OE;
output [17:0] DRAM_DQ_OE;
output [2:0] DRAM_DQS_OE;
output I2C0_SCL_USBC_DATA1_MGPIO31B_OE;
output I2C0_SDA_USBC_DATA0_MGPIO30B_OE;
output I2C1_SCL_USBA_DATA4_MGPIO1A_OE;
output I2C1_SDA_USBA_DATA3_MGPIO0A_OE;
output MMUART0_CTS_USBC_DATA7_MGPIO19B_OE;
output MMUART0_DCD_MGPIO22B_OE;
output MMUART0_DSR_MGPIO20B_OE;
output MMUART0_DTR_USBC_DATA6_MGPIO18B_OE;
output MMUART0_RI_MGPIO21B_OE;
output MMUART0_RTS_USBC_DATA5_MGPIO17B_OE;
output MMUART0_RXD_USBC_STP_MGPIO28B_OE;
output MMUART0_SCK_USBC_NXT_MGPIO29B_OE;
output MMUART0_TXD_USBC_DIR_MGPIO27B_OE;
output MMUART1_RXD_USBC_DATA3_MGPIO26B_OE;
output MMUART1_SCK_USBC_DATA4_MGPIO25B_OE;
output MMUART1_TXD_USBC_DATA2_MGPIO24B_OE;
output RGMII_GTX_CLK_RMII_CLK_USBB_XCLK_OE;
output RGMII_MDC_RMII_MDC_OE;
output RGMII_MDIO_RMII_MDIO_USBB_DATA7_OE;
output RGMII_RX_CLK_OE;
output RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_OE;
output RGMII_RXD0_RMII_RXD0_USBB_DATA0_OE;
output RGMII_RXD1_RMII_RXD1_USBB_DATA1_OE;
output RGMII_RXD2_RMII_RX_ER_USBB_DATA3_OE;
output RGMII_RXD3_USBB_DATA4_OE;
output RGMII_TX_CLK_OE;
output RGMII_TX_CTL_RMII_TX_EN_USBB_NXT_OE;
output RGMII_TXD0_RMII_TXD0_USBB_DIR_OE;
output RGMII_TXD1_RMII_TXD1_USBB_STP_OE;
output RGMII_TXD2_USBB_DATA5_OE;
output RGMII_TXD3_USBB_DATA6_OE;
output SPI0_SCK_USBA_XCLK_OE;
output SPI0_SDI_USBA_DIR_MGPIO5A_OE;
output SPI0_SDO_USBA_STP_MGPIO6A_OE;
output SPI0_SS0_USBA_NXT_MGPIO7A_OE;
output SPI0_SS1_USBA_DATA5_MGPIO8A_OE;
output SPI0_SS2_USBA_DATA6_MGPIO9A_OE;
output SPI0_SS3_USBA_DATA7_MGPIO10A_OE;
output SPI1_SCK_OE;
output SPI1_SDI_MGPIO11A_OE;
output SPI1_SDO_MGPIO12A_OE;
output SPI1_SS0_MGPIO13A_OE;
output SPI1_SS1_MGPIO14A_OE;
output SPI1_SS2_MGPIO15A_OE;
output SPI1_SS3_MGPIO16A_OE;
output SPI1_SS4_MGPIO17A_OE;
output SPI1_SS5_MGPIO18A_OE;
output SPI1_SS6_MGPIO23A_OE;
output SPI1_SS7_MGPIO24A_OE;
output USBC_XCLK_OE;

    parameter INIT = 'h0 ;
    parameter ACT_UBITS = 'hFFFFFFFFFFFFFF ;
    parameter MEMORYFILE = "" ;
    parameter RTC_MAIN_XTL_FREQ = 0.0 ;
    parameter RTC_MAIN_XTL_MODE = "1" ;
    
endmodule


module COREAPB3_MUXPTOB3(
       GPOUT_reg,
       INTR_reg,
       CoreAPB3_0_APBmslave5_PRDATA_m_d_0,
       CoreAPB3_0_APBmslave3_PRDATA_2,
       CoreAPB3_0_APBmslave3_PRDATA_3,
       CoreAPB3_0_APBmslave3_PRDATA_0,
       CoreAPB3_0_APBmslave2_PADDR_1,
       CoreAPB3_0_APBmslave2_PADDR_2,
       CoreAPB3_0_APBmslave2_PADDR_0,
       CoreAPB3_0_APBmslave2_PADDR_3,
       CoreAPB3_0_APBmslave2_PADDR_5,
       PRDATA_reg_4,
       PRDATA_reg_0,
       PRDATA_reg_3,
       PRDATA_reg_1,
       PRDATA_reg_5,
       PRDATA_reg_10,
       PRDATA_reg_19,
       PRDATA_reg_20,
       PRDATA_reg_6,
       PRDATA_reg_17,
       PRDATA_reg_18,
       PRDATA_reg_7,
       PRDATA_reg_15,
       PRDATA_reg_16,
       PRDATA_reg_8,
       PRDATA_reg_13,
       PRDATA_reg_14,
       PRDATA_reg_9,
       PRDATA_reg_11,
       PRDATA_reg_12,
       PRDATA_reg_21,
       PRDATA_reg_22,
       PRDATA_reg_23,
       PRDATA_reg_24,
       PRDATA_reg_25,
       PRDATA_reg_26,
       PRDATA_reg_27,
       PRDATA_reg_28,
       lsram_width32_PRDATA_4,
       lsram_width32_PRDATA_0,
       lsram_width32_PRDATA_3,
       lsram_width32_PRDATA_1,
       lsram_width32_PRDATA_5,
       lsram_width32_PRDATA_10,
       lsram_width32_PRDATA_19,
       lsram_width32_PRDATA_20,
       lsram_width32_PRDATA_6,
       lsram_width32_PRDATA_17,
       lsram_width32_PRDATA_18,
       lsram_width32_PRDATA_7,
       lsram_width32_PRDATA_15,
       lsram_width32_PRDATA_16,
       lsram_width32_PRDATA_8,
       lsram_width32_PRDATA_13,
       lsram_width32_PRDATA_14,
       lsram_width32_PRDATA_9,
       lsram_width32_PRDATA_11,
       lsram_width32_PRDATA_12,
       lsram_width32_PRDATA_21,
       lsram_width32_PRDATA_22,
       lsram_width32_PRDATA_23,
       lsram_width32_PRDATA_24,
       lsram_width32_PRDATA_25,
       lsram_width32_PRDATA_26,
       lsram_width32_PRDATA_27,
       lsram_width32_PRDATA_28,
       FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_4,
       FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_9,
       FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_18,
       FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_19,
       FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_5,
       FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_16,
       FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_17,
       FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_6,
       FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_14,
       FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_15,
       FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_7,
       FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_12,
       FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_13,
       FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_8,
       FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_10,
       FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_11,
       FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_20,
       FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_21,
       FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_22,
       FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_23,
       FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_24,
       FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_25,
       FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_26,
       FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_27,
       FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_0,
       FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_3,
       CoreAPB3_0_APBmslave2_PENABLE,
       CoreAPB3_0_APBmslave2_PWRITE,
       PRDATA4_out,
       iPRDATA29,
       PRDATA_N_8_mux_0,
       CoreAPB3_m8_0,
       CoreAPB3_N_8_0_i_1,
       CoreAPB3_N_3_i_0_li_0,
       CoreAPB3_N_8_0_i_0,
       N_4762,
       N_4738,
       N_4706,
       N_4682,
       N_4882,
       N_4858,
       N_4826,
       N_4802,
       CoreAPB3_0_APBmslave3_PSELx,
       CoreAPB3_0_APBmslave5_PSELx,
       N_245,
       PRDATA_m1_e_1,
       CoreAPB3_m2_0_a2_1_1,
       N_247,
       CoreAPB3_0_APBmslave3_PREADY,
       CoreAPB3_0_APBmslave2_PREADY,
       PREADY_0_iv_i_0,
       \CONFIG_reg[4]2_0_a4_0_a2_0_RNIBB9M2 ,
       CoreAPB3_m6_0_ns,
       N_452
    );
input  [31:8] GPOUT_reg;
input  [31:7] INTR_reg;
input  [4:4] CoreAPB3_0_APBmslave5_PRDATA_m_d_0;
input  CoreAPB3_0_APBmslave3_PRDATA_2;
input  CoreAPB3_0_APBmslave3_PRDATA_3;
input  CoreAPB3_0_APBmslave3_PRDATA_0;
input  CoreAPB3_0_APBmslave2_PADDR_1;
input  CoreAPB3_0_APBmslave2_PADDR_2;
input  CoreAPB3_0_APBmslave2_PADDR_0;
input  CoreAPB3_0_APBmslave2_PADDR_3;
input  CoreAPB3_0_APBmslave2_PADDR_5;
input  PRDATA_reg_4;
input  PRDATA_reg_0;
input  PRDATA_reg_3;
input  PRDATA_reg_1;
input  PRDATA_reg_5;
input  PRDATA_reg_10;
input  PRDATA_reg_19;
input  PRDATA_reg_20;
input  PRDATA_reg_6;
input  PRDATA_reg_17;
input  PRDATA_reg_18;
input  PRDATA_reg_7;
input  PRDATA_reg_15;
input  PRDATA_reg_16;
input  PRDATA_reg_8;
input  PRDATA_reg_13;
input  PRDATA_reg_14;
input  PRDATA_reg_9;
input  PRDATA_reg_11;
input  PRDATA_reg_12;
input  PRDATA_reg_21;
input  PRDATA_reg_22;
input  PRDATA_reg_23;
input  PRDATA_reg_24;
input  PRDATA_reg_25;
input  PRDATA_reg_26;
input  PRDATA_reg_27;
input  PRDATA_reg_28;
input  lsram_width32_PRDATA_4;
input  lsram_width32_PRDATA_0;
input  lsram_width32_PRDATA_3;
input  lsram_width32_PRDATA_1;
input  lsram_width32_PRDATA_5;
input  lsram_width32_PRDATA_10;
input  lsram_width32_PRDATA_19;
input  lsram_width32_PRDATA_20;
input  lsram_width32_PRDATA_6;
input  lsram_width32_PRDATA_17;
input  lsram_width32_PRDATA_18;
input  lsram_width32_PRDATA_7;
input  lsram_width32_PRDATA_15;
input  lsram_width32_PRDATA_16;
input  lsram_width32_PRDATA_8;
input  lsram_width32_PRDATA_13;
input  lsram_width32_PRDATA_14;
input  lsram_width32_PRDATA_9;
input  lsram_width32_PRDATA_11;
input  lsram_width32_PRDATA_12;
input  lsram_width32_PRDATA_21;
input  lsram_width32_PRDATA_22;
input  lsram_width32_PRDATA_23;
input  lsram_width32_PRDATA_24;
input  lsram_width32_PRDATA_25;
input  lsram_width32_PRDATA_26;
input  lsram_width32_PRDATA_27;
input  lsram_width32_PRDATA_28;
output FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_4;
output FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_9;
output FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_18;
output FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_19;
output FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_5;
output FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_16;
output FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_17;
output FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_6;
output FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_14;
output FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_15;
output FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_7;
output FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_12;
output FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_13;
output FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_8;
output FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_10;
output FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_11;
output FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_20;
output FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_21;
output FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_22;
output FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_23;
output FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_24;
output FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_25;
output FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_26;
output FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_27;
output FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_0;
output FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_3;
input  CoreAPB3_0_APBmslave2_PENABLE;
input  CoreAPB3_0_APBmslave2_PWRITE;
input  PRDATA4_out;
input  iPRDATA29;
output PRDATA_N_8_mux_0;
input  CoreAPB3_m8_0;
input  CoreAPB3_N_8_0_i_1;
input  CoreAPB3_N_3_i_0_li_0;
output CoreAPB3_N_8_0_i_0;
input  N_4762;
input  N_4738;
input  N_4706;
input  N_4682;
input  N_4882;
input  N_4858;
input  N_4826;
input  N_4802;
input  CoreAPB3_0_APBmslave3_PSELx;
input  CoreAPB3_0_APBmslave5_PSELx;
input  N_245;
input  PRDATA_m1_e_1;
input  CoreAPB3_m2_0_a2_1_1;
input  N_247;
input  CoreAPB3_0_APBmslave3_PREADY;
input  CoreAPB3_0_APBmslave2_PREADY;
output PREADY_0_iv_i_0;
input  \CONFIG_reg[4]2_0_a4_0_a2_0_RNIBB9M2 ;
input  CoreAPB3_m6_0_ns;
input  N_452;

    wire \PRDATA_0_iv_1_0_RNO[7]_net_1 , CoreAPB3_m7_0_1, 
        PRDATA_m4_am_1_1_net_1, PRDATA_m4_am_net_1, 
        PRDATA_m4_bm_1_1_net_1, PRDATA_m4_bm_net_1, PRDATA_m4_ns_net_1, 
        CoreAPB3_m4_2_0, CoreAPB3_m4_10_0, CoreAPB3_m4_5_0, 
        CoreAPB3_m4_1_0, CoreAPB3_m4_9_0, CoreAPB3_m4_13_0, 
        CoreAPB3_m4_4_0, CoreAPB3_m4_0_0, CoreAPB3_m4_12_0, 
        CoreAPB3_m4_11_0, CoreAPB3_m4_3_0, CoreAPB3_m4_0, 
        CoreAPB3_m4_6_0, CoreAPB3_m4_0_1, CoreAPB3_m4_5_0_0, 
        CoreAPB3_m4_8_0, CoreAPB3_m4_3_0_0, CoreAPB3_m4_14_0, 
        CoreAPB3_m4_1_0_0, CoreAPB3_m4_0_0_0, CoreAPB3_m4_2_0_0, 
        CoreAPB3_m4_6_0_0, CoreAPB3_m4_7_0, CoreAPB3_m4_4_0_0, 
        PRDATA_m2_1_net_1, PRDATA_m2_net_1, CoreAPB3_m7_0_0, 
        \PRDATA_0_iv_1_0[7]_net_1 , 
        \CoreAPB3_0_APBmslave5_PRDATA_m_0[4] , PRDATA_m6_i_0_1_net_1, 
        \PRDATA_0_iv_1_1[7]_net_1 , 
        \CoreAPB3_0_APBmslave5_PRDATA_m_1[4] , 
        \CoreAPB3_0_APBmslave2_PRDATA_m[8] , 
        \CoreAPB3_0_APBmslave2_PRDATA_m[13] , 
        \CoreAPB3_0_APBmslave2_PRDATA_m[22] , 
        \CoreAPB3_0_APBmslave2_PRDATA_m[23] , 
        \CoreAPB3_0_APBmslave2_PRDATA_m[9] , 
        \CoreAPB3_0_APBmslave2_PRDATA_m[20] , 
        \CoreAPB3_0_APBmslave2_PRDATA_m[21] , 
        \CoreAPB3_0_APBmslave2_PRDATA_m[10] , 
        \CoreAPB3_0_APBmslave2_PRDATA_m[18] , 
        \CoreAPB3_0_APBmslave2_PRDATA_m[19] , 
        \CoreAPB3_0_APBmslave2_PRDATA_m[11] , 
        \CoreAPB3_0_APBmslave2_PRDATA_m[16] , 
        \CoreAPB3_0_APBmslave2_PRDATA_m[17] , 
        \CoreAPB3_0_APBmslave2_PRDATA_m[12] , 
        \CoreAPB3_0_APBmslave2_PRDATA_m[14] , 
        \CoreAPB3_0_APBmslave2_PRDATA_m[15] , 
        \CoreAPB3_0_APBmslave2_PRDATA_m[24] , 
        \CoreAPB3_0_APBmslave2_PRDATA_m[25] , 
        \CoreAPB3_0_APBmslave2_PRDATA_m[26] , 
        \CoreAPB3_0_APBmslave2_PRDATA_m[27] , 
        \CoreAPB3_0_APBmslave2_PRDATA_m[28] , 
        \CoreAPB3_0_APBmslave2_PRDATA_m[29] , 
        \CoreAPB3_0_APBmslave2_PRDATA_m[30] , 
        \CoreAPB3_0_APBmslave2_PRDATA_m[31] , GND_net_1, VCC_net_1;
    
    CFG4 #( .INIT(16'h0A0C) )  \PRDATA_0_iv_RNO[31]  (.A(GPOUT_reg[31])
        , .B(INTR_reg[31]), .C(CoreAPB3_0_APBmslave2_PADDR_2), .D(
        CoreAPB3_0_APBmslave2_PADDR_3), .Y(CoreAPB3_m4_5_0));
    CFG4 #( .INIT(16'h0A0C) )  \PRDATA_0_iv_RNO[13]  (.A(GPOUT_reg[13])
        , .B(INTR_reg[13]), .C(CoreAPB3_0_APBmslave2_PADDR_2), .D(
        CoreAPB3_0_APBmslave2_PADDR_3), .Y(CoreAPB3_m4_1_0_0));
    CFG4 #( .INIT(16'hF0F8) )  \PRDATA_0_iv[12]  (.A(
        CoreAPB3_0_APBmslave5_PSELx), .B(CoreAPB3_m4_12_0), .C(
        \CoreAPB3_0_APBmslave2_PRDATA_m[12] ), .D(N_245), .Y(
        FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_8));
    CFG4 #( .INIT(16'h34F4) )  PRDATA_m4_am (.A(N_4762), .B(
        CoreAPB3_0_APBmslave2_PADDR_1), .C(PRDATA_m4_am_1_1_net_1), .D(
        N_4738), .Y(PRDATA_m4_am_net_1));
    CFG4 #( .INIT(16'h0A0C) )  \PRDATA_0_iv_RNO[14]  (.A(GPOUT_reg[14])
        , .B(INTR_reg[14]), .C(CoreAPB3_0_APBmslave2_PADDR_2), .D(
        CoreAPB3_0_APBmslave2_PADDR_3), .Y(CoreAPB3_m4_9_0));
    CFG4 #( .INIT(16'hF0F8) )  \PRDATA_0_iv[19]  (.A(
        CoreAPB3_0_APBmslave5_PSELx), .B(CoreAPB3_m4_10_0), .C(
        \CoreAPB3_0_APBmslave2_PRDATA_m[19] ), .D(N_245), .Y(
        FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_15));
    CFG4 #( .INIT(16'h0A0C) )  \PRDATA_0_iv_RNO[19]  (.A(GPOUT_reg[19])
        , .B(INTR_reg[19]), .C(CoreAPB3_0_APBmslave2_PADDR_2), .D(
        CoreAPB3_0_APBmslave2_PADDR_3), .Y(CoreAPB3_m4_10_0));
    CFG4 #( .INIT(16'hC840) )  \PRDATA_0_iv_RNO_0[13]  (.A(PRDATA4_out)
        , .B(iPRDATA29), .C(PRDATA_reg_10), .D(lsram_width32_PRDATA_10)
        , .Y(\CoreAPB3_0_APBmslave2_PRDATA_m[13] ));
    CFG4 #( .INIT(16'h0A0C) )  \PRDATA_0_iv_RNO[9]  (.A(GPOUT_reg[9]), 
        .B(INTR_reg[9]), .C(CoreAPB3_0_APBmslave2_PADDR_2), .D(
        CoreAPB3_0_APBmslave2_PADDR_3), .Y(CoreAPB3_m4_0_1));
    CFG4 #( .INIT(16'h0A0C) )  \PRDATA_0_iv_RNO[26]  (.A(GPOUT_reg[26])
        , .B(INTR_reg[26]), .C(CoreAPB3_0_APBmslave2_PADDR_2), .D(
        CoreAPB3_0_APBmslave2_PADDR_3), .Y(CoreAPB3_m4_6_0));
    CFG4 #( .INIT(16'h2A0A) )  PRDATA_m6_i_0_1 (.A(
        CoreAPB3_0_APBmslave5_PSELx), .B(N_245), .C(
        CoreAPB3_0_APBmslave2_PADDR_5), .D(PRDATA_m1_e_1), .Y(
        PRDATA_m6_i_0_1_net_1));
    CFG4 #( .INIT(16'hF070) )  PRDATA_m2_1_RNIJAJR4 (.A(
        CoreAPB3_0_APBmslave5_PSELx), .B(CoreAPB3_m2_0_a2_1_1), .C(
        CoreAPB3_m7_0_0), .D(N_245), .Y(CoreAPB3_m7_0_1));
    CFG4 #( .INIT(16'hC840) )  \PRDATA_0_iv_RNO_0[16]  (.A(PRDATA4_out)
        , .B(iPRDATA29), .C(PRDATA_reg_13), .D(lsram_width32_PRDATA_13)
        , .Y(\CoreAPB3_0_APBmslave2_PRDATA_m[16] ));
    CFG4 #( .INIT(16'hFF8A) )  \PRDATA_0_iv_1[7]  (.A(
        PRDATA_m6_i_0_1_net_1), .B(N_452), .C(PRDATA_m4_ns_net_1), .D(
        \PRDATA_0_iv_1_1[7]_net_1 ), .Y(
        FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_3));
    CFG4 #( .INIT(16'hC840) )  \PRDATA_0_iv_RNO_0[19]  (.A(PRDATA4_out)
        , .B(iPRDATA29), .C(PRDATA_reg_16), .D(lsram_width32_PRDATA_16)
        , .Y(\CoreAPB3_0_APBmslave2_PRDATA_m[19] ));
    CFG4 #( .INIT(16'hC840) )  \PRDATA_0_iv_RNO_0[12]  (.A(PRDATA4_out)
        , .B(iPRDATA29), .C(PRDATA_reg_9), .D(lsram_width32_PRDATA_9), 
        .Y(\CoreAPB3_0_APBmslave2_PRDATA_m[12] ));
    CFG4 #( .INIT(16'hC840) )  \PRDATA_0_iv_RNO_0[23]  (.A(PRDATA4_out)
        , .B(iPRDATA29), .C(PRDATA_reg_20), .D(lsram_width32_PRDATA_20)
        , .Y(\CoreAPB3_0_APBmslave2_PRDATA_m[23] ));
    CFG4 #( .INIT(16'hC840) )  \PRDATA_0_iv_RNO_0[26]  (.A(PRDATA4_out)
        , .B(iPRDATA29), .C(PRDATA_reg_23), .D(lsram_width32_PRDATA_23)
        , .Y(\CoreAPB3_0_APBmslave2_PRDATA_m[26] ));
    CFG4 #( .INIT(16'h0A0C) )  \PRDATA_0_iv_RNO[20]  (.A(GPOUT_reg[20])
        , .B(INTR_reg[20]), .C(CoreAPB3_0_APBmslave2_PADDR_2), .D(
        CoreAPB3_0_APBmslave2_PADDR_3), .Y(CoreAPB3_m4_8_0));
    CFG4 #( .INIT(16'hC840) )  \PRDATA_0_iv_RNO_0[17]  (.A(PRDATA4_out)
        , .B(iPRDATA29), .C(PRDATA_reg_14), .D(lsram_width32_PRDATA_14)
        , .Y(\CoreAPB3_0_APBmslave2_PRDATA_m[17] ));
    CFG4 #( .INIT(16'hC840) )  \PRDATA_0_iv_RNO_0[10]  (.A(PRDATA4_out)
        , .B(iPRDATA29), .C(PRDATA_reg_7), .D(lsram_width32_PRDATA_7), 
        .Y(\CoreAPB3_0_APBmslave2_PRDATA_m[10] ));
    CFG4 #( .INIT(16'hC840) )  \PRDATA_0_iv_RNO_0[29]  (.A(PRDATA4_out)
        , .B(iPRDATA29), .C(PRDATA_reg_26), .D(lsram_width32_PRDATA_26)
        , .Y(\CoreAPB3_0_APBmslave2_PRDATA_m[29] ));
    CFG4 #( .INIT(16'hC840) )  \PRDATA_0_iv_RNO_0[22]  (.A(PRDATA4_out)
        , .B(iPRDATA29), .C(PRDATA_reg_19), .D(lsram_width32_PRDATA_19)
        , .Y(\CoreAPB3_0_APBmslave2_PRDATA_m[22] ));
    CFG4 #( .INIT(16'hF0F8) )  \PRDATA_0_iv[18]  (.A(
        CoreAPB3_0_APBmslave5_PSELx), .B(CoreAPB3_m4_14_0), .C(
        \CoreAPB3_0_APBmslave2_PRDATA_m[18] ), .D(N_245), .Y(
        FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_14));
    CFG4 #( .INIT(16'hF0F8) )  \PRDATA_0_iv[16]  (.A(
        CoreAPB3_0_APBmslave5_PSELx), .B(CoreAPB3_m4_2_0_0), .C(
        \CoreAPB3_0_APBmslave2_PRDATA_m[16] ), .D(N_245), .Y(
        FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_12));
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'hF0F8) )  \PRDATA_0_iv[11]  (.A(
        CoreAPB3_0_APBmslave5_PSELx), .B(CoreAPB3_m4_3_0_0), .C(
        \CoreAPB3_0_APBmslave2_PRDATA_m[11] ), .D(N_245), .Y(
        FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_7));
    CFG4 #( .INIT(16'hF0F8) )  \PRDATA_0_iv[10]  (.A(
        CoreAPB3_0_APBmslave5_PSELx), .B(CoreAPB3_m4_13_0), .C(
        \CoreAPB3_0_APBmslave2_PRDATA_m[10] ), .D(N_245), .Y(
        FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_6));
    CFG4 #( .INIT(16'hC840) )  \PRDATA_0_iv_RNO_0[27]  (.A(PRDATA4_out)
        , .B(iPRDATA29), .C(PRDATA_reg_24), .D(lsram_width32_PRDATA_24)
        , .Y(\CoreAPB3_0_APBmslave2_PRDATA_m[27] ));
    CFG4 #( .INIT(16'hC840) )  \PRDATA_0_iv_RNO_0[20]  (.A(PRDATA4_out)
        , .B(iPRDATA29), .C(PRDATA_reg_17), .D(lsram_width32_PRDATA_17)
        , .Y(\CoreAPB3_0_APBmslave2_PRDATA_m[20] ));
    CFG4 #( .INIT(16'hF351) )  PREADY_0_iv_i (.A(iPRDATA29), .B(
        CoreAPB3_0_APBmslave3_PSELx), .C(CoreAPB3_0_APBmslave3_PREADY), 
        .D(CoreAPB3_0_APBmslave2_PREADY), .Y(PREADY_0_iv_i_0));
    CFG4 #( .INIT(16'hDCCC) )  PRDATA_m2_RNI74LF4 (.A(N_245), .B(
        \CoreAPB3_0_APBmslave5_PRDATA_m_0[4] ), .C(
        CoreAPB3_0_APBmslave5_PRDATA_m_d_0[4]), .D(
        CoreAPB3_0_APBmslave5_PSELx), .Y(
        \CoreAPB3_0_APBmslave5_PRDATA_m_1[4] ));
    CFG4 #( .INIT(16'h0A0C) )  \PRDATA_0_iv_RNO[16]  (.A(GPOUT_reg[16])
        , .B(INTR_reg[16]), .C(CoreAPB3_0_APBmslave2_PADDR_2), .D(
        CoreAPB3_0_APBmslave2_PADDR_3), .Y(CoreAPB3_m4_2_0_0));
    CFG4 #( .INIT(16'hFCFE) )  PRDATA_m2_RNI6H2OT (.A(CoreAPB3_m8_0), 
        .B(\CONFIG_reg[4]2_0_a4_0_a2_0_RNIBB9M2 ), .C(
        \CoreAPB3_0_APBmslave5_PRDATA_m_1[4] ), .D(CoreAPB3_m6_0_ns), 
        .Y(FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_0));
    CFG4 #( .INIT(16'hF0F8) )  \PRDATA_0_iv[14]  (.A(
        CoreAPB3_0_APBmslave5_PSELx), .B(CoreAPB3_m4_9_0), .C(
        \CoreAPB3_0_APBmslave2_PRDATA_m[14] ), .D(N_245), .Y(
        FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_10));
    CFG4 #( .INIT(16'h4657) )  PRDATA_m4_bm_1_1 (.A(
        CoreAPB3_0_APBmslave2_PADDR_2), .B(
        CoreAPB3_0_APBmslave2_PADDR_1), .C(N_4826), .D(N_4802), .Y(
        PRDATA_m4_bm_1_1_net_1));
    CFG4 #( .INIT(16'hC840) )  \PRDATA_0_iv_RNO_0[31]  (.A(PRDATA4_out)
        , .B(iPRDATA29), .C(PRDATA_reg_28), .D(lsram_width32_PRDATA_28)
        , .Y(\CoreAPB3_0_APBmslave2_PRDATA_m[31] ));
    CFG4 #( .INIT(16'h0A0C) )  \PRDATA_0_iv_RNO[10]  (.A(GPOUT_reg[10])
        , .B(INTR_reg[10]), .C(CoreAPB3_0_APBmslave2_PADDR_2), .D(
        CoreAPB3_0_APBmslave2_PADDR_3), .Y(CoreAPB3_m4_13_0));
    CFG4 #( .INIT(16'h0A0C) )  \PRDATA_0_iv_RNO[8]  (.A(GPOUT_reg[8]), 
        .B(INTR_reg[8]), .C(CoreAPB3_0_APBmslave2_PADDR_2), .D(
        CoreAPB3_0_APBmslave2_PADDR_3), .Y(CoreAPB3_m4_6_0_0));
    CFG4 #( .INIT(16'h0A0C) )  \PRDATA_0_iv_RNO[30]  (.A(GPOUT_reg[30])
        , .B(INTR_reg[30]), .C(CoreAPB3_0_APBmslave2_PADDR_2), .D(
        CoreAPB3_0_APBmslave2_PADDR_3), .Y(CoreAPB3_m4_0_0_0));
    CFG4 #( .INIT(16'hF0F8) )  \PRDATA_0_iv[9]  (.A(
        CoreAPB3_0_APBmslave5_PSELx), .B(CoreAPB3_m4_0_1), .C(
        \CoreAPB3_0_APBmslave2_PRDATA_m[9] ), .D(N_245), .Y(
        FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_5));
    CFG4 #( .INIT(16'h0A0C) )  \PRDATA_0_iv_RNO[28]  (.A(GPOUT_reg[28])
        , .B(INTR_reg[28]), .C(CoreAPB3_0_APBmslave2_PADDR_2), .D(
        CoreAPB3_0_APBmslave2_PADDR_3), .Y(CoreAPB3_m4_2_0));
    CFG4 #( .INIT(16'h0A0C) )  \PRDATA_0_iv_RNO[22]  (.A(GPOUT_reg[22])
        , .B(INTR_reg[22]), .C(CoreAPB3_0_APBmslave2_PADDR_2), .D(
        CoreAPB3_0_APBmslave2_PADDR_3), .Y(CoreAPB3_m4_4_0));
    CFG4 #( .INIT(16'hF0F8) )  \PRDATA_0_iv[22]  (.A(
        CoreAPB3_0_APBmslave5_PSELx), .B(CoreAPB3_m4_4_0), .C(
        \CoreAPB3_0_APBmslave2_PRDATA_m[22] ), .D(N_245), .Y(
        FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_18));
    CFG4 #( .INIT(16'hC840) )  \PRDATA_0_iv_RNO_0[18]  (.A(PRDATA4_out)
        , .B(iPRDATA29), .C(PRDATA_reg_15), .D(lsram_width32_PRDATA_15)
        , .Y(\CoreAPB3_0_APBmslave2_PRDATA_m[18] ));
    CFG4 #( .INIT(16'hF0F8) )  \PRDATA_0_iv[13]  (.A(
        CoreAPB3_0_APBmslave5_PSELx), .B(CoreAPB3_m4_1_0_0), .C(
        \CoreAPB3_0_APBmslave2_PRDATA_m[13] ), .D(N_245), .Y(
        FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_9));
    CFG4 #( .INIT(16'hF0F8) )  \PRDATA_0_iv[29]  (.A(
        CoreAPB3_0_APBmslave5_PSELx), .B(CoreAPB3_m4_0), .C(
        \CoreAPB3_0_APBmslave2_PRDATA_m[29] ), .D(N_245), .Y(
        FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_25));
    CFG4 #( .INIT(16'h2A3F) )  PRDATA_m2_1_RNIQL321 (.A(
        PRDATA_m2_1_net_1), .B(CoreAPB3_0_APBmslave3_PRDATA_2), .C(
        CoreAPB3_0_APBmslave3_PSELx), .D(iPRDATA29), .Y(
        CoreAPB3_m7_0_0));
    CFG4 #( .INIT(16'hC840) )  \PRDATA_0_iv_RNO_0[14]  (.A(PRDATA4_out)
        , .B(iPRDATA29), .C(PRDATA_reg_11), .D(lsram_width32_PRDATA_11)
        , .Y(\CoreAPB3_0_APBmslave2_PRDATA_m[14] ));
    CFG4 #( .INIT(16'hF0F8) )  \PRDATA_0_iv[15]  (.A(
        CoreAPB3_0_APBmslave5_PSELx), .B(CoreAPB3_m4_11_0), .C(
        \CoreAPB3_0_APBmslave2_PRDATA_m[15] ), .D(N_245), .Y(
        FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_11));
    CFG4 #( .INIT(16'h0A0C) )  \PRDATA_0_iv_RNO[27]  (.A(GPOUT_reg[27])
        , .B(INTR_reg[27]), .C(CoreAPB3_0_APBmslave2_PADDR_2), .D(
        CoreAPB3_0_APBmslave2_PADDR_3), .Y(CoreAPB3_m4_3_0));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'hD5C0) )  PRDATA_m2_RNI82L11 (.A(PRDATA_m2_net_1), 
        .B(CoreAPB3_0_APBmslave3_PRDATA_0), .C(
        CoreAPB3_0_APBmslave3_PSELx), .D(iPRDATA29), .Y(
        \CoreAPB3_0_APBmslave5_PRDATA_m_0[4] ));
    CFG4 #( .INIT(16'hFF08) )  \PRDATA_0_iv_1_1[7]  (.A(INTR_reg[7]), 
        .B(CoreAPB3_0_APBmslave5_PSELx), .C(N_247), .D(
        \PRDATA_0_iv_1_0[7]_net_1 ), .Y(\PRDATA_0_iv_1_1[7]_net_1 ));
    CFG4 #( .INIT(16'hF0F8) )  \PRDATA_0_iv[17]  (.A(
        CoreAPB3_0_APBmslave5_PSELx), .B(CoreAPB3_m4_7_0), .C(
        \CoreAPB3_0_APBmslave2_PRDATA_m[17] ), .D(N_245), .Y(
        FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_13));
    CFG4 #( .INIT(16'hBF3F) )  PRDATA_m2_1_RNIF0DK01 (.A(CoreAPB3_m8_0)
        , .B(CoreAPB3_m7_0_1), .C(CoreAPB3_N_8_0_i_1), .D(
        CoreAPB3_N_3_i_0_li_0), .Y(CoreAPB3_N_8_0_i_0));
    CFG4 #( .INIT(16'hC840) )  \PRDATA_0_iv_RNO_0[28]  (.A(PRDATA4_out)
        , .B(iPRDATA29), .C(PRDATA_reg_25), .D(lsram_width32_PRDATA_25)
        , .Y(\CoreAPB3_0_APBmslave2_PRDATA_m[28] ));
    CFG4 #( .INIT(16'hC840) )  g0 (.A(PRDATA4_out), .B(iPRDATA29), .C(
        PRDATA_reg_0), .D(lsram_width32_PRDATA_0), .Y(PRDATA_N_8_mux_0)
        );
    CFG4 #( .INIT(16'hC840) )  \PRDATA_0_iv_RNO_0[8]  (.A(PRDATA4_out), 
        .B(iPRDATA29), .C(PRDATA_reg_5), .D(lsram_width32_PRDATA_5), 
        .Y(\CoreAPB3_0_APBmslave2_PRDATA_m[8] ));
    CFG4 #( .INIT(16'hC840) )  \PRDATA_0_iv_RNO_0[24]  (.A(PRDATA4_out)
        , .B(iPRDATA29), .C(PRDATA_reg_21), .D(lsram_width32_PRDATA_21)
        , .Y(\CoreAPB3_0_APBmslave2_PRDATA_m[24] ));
    CFG3 #( .INIT(8'hE2) )  PRDATA_m4_ns (.A(PRDATA_m4_am_net_1), .B(
        CoreAPB3_0_APBmslave2_PADDR_0), .C(PRDATA_m4_bm_net_1), .Y(
        PRDATA_m4_ns_net_1));
    CFG4 #( .INIT(16'h4657) )  PRDATA_m4_am_1_1 (.A(
        CoreAPB3_0_APBmslave2_PADDR_2), .B(
        CoreAPB3_0_APBmslave2_PADDR_1), .C(N_4706), .D(N_4682), .Y(
        PRDATA_m4_am_1_1_net_1));
    CFG4 #( .INIT(16'hC840) )  \PRDATA_0_iv_RNO_0[9]  (.A(PRDATA4_out), 
        .B(iPRDATA29), .C(PRDATA_reg_6), .D(lsram_width32_PRDATA_6), 
        .Y(\CoreAPB3_0_APBmslave2_PRDATA_m[9] ));
    CFG4 #( .INIT(16'hC840) )  \PRDATA_0_iv_RNO_0[15]  (.A(PRDATA4_out)
        , .B(iPRDATA29), .C(PRDATA_reg_12), .D(lsram_width32_PRDATA_12)
        , .Y(\CoreAPB3_0_APBmslave2_PRDATA_m[15] ));
    CFG4 #( .INIT(16'hF0F8) )  \PRDATA_0_iv[28]  (.A(
        CoreAPB3_0_APBmslave5_PSELx), .B(CoreAPB3_m4_2_0), .C(
        \CoreAPB3_0_APBmslave2_PRDATA_m[28] ), .D(N_245), .Y(
        FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_24));
    CFG4 #( .INIT(16'h34F4) )  PRDATA_m4_bm (.A(N_4882), .B(
        CoreAPB3_0_APBmslave2_PADDR_1), .C(PRDATA_m4_bm_1_1_net_1), .D(
        N_4858), .Y(PRDATA_m4_bm_net_1));
    CFG4 #( .INIT(16'hC840) )  \PRDATA_0_iv_RNO_0[25]  (.A(PRDATA4_out)
        , .B(iPRDATA29), .C(PRDATA_reg_22), .D(lsram_width32_PRDATA_22)
        , .Y(\CoreAPB3_0_APBmslave2_PRDATA_m[25] ));
    CFG4 #( .INIT(16'h0A0C) )  \PRDATA_0_iv_RNO[18]  (.A(GPOUT_reg[18])
        , .B(INTR_reg[18]), .C(CoreAPB3_0_APBmslave2_PADDR_2), .D(
        CoreAPB3_0_APBmslave2_PADDR_3), .Y(CoreAPB3_m4_14_0));
    CFG4 #( .INIT(16'h0A0C) )  \PRDATA_0_iv_RNO[12]  (.A(GPOUT_reg[12])
        , .B(INTR_reg[12]), .C(CoreAPB3_0_APBmslave2_PADDR_2), .D(
        CoreAPB3_0_APBmslave2_PADDR_3), .Y(CoreAPB3_m4_12_0));
    CFG4 #( .INIT(16'hF0F8) )  \PRDATA_0_iv[26]  (.A(
        CoreAPB3_0_APBmslave5_PSELx), .B(CoreAPB3_m4_6_0), .C(
        \CoreAPB3_0_APBmslave2_PRDATA_m[26] ), .D(N_245), .Y(
        FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_22));
    CFG4 #( .INIT(16'hF0F8) )  \PRDATA_0_iv[21]  (.A(
        CoreAPB3_0_APBmslave5_PSELx), .B(CoreAPB3_m4_5_0_0), .C(
        \CoreAPB3_0_APBmslave2_PRDATA_m[21] ), .D(N_245), .Y(
        FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_17));
    CFG4 #( .INIT(16'hF0F8) )  \PRDATA_0_iv[20]  (.A(
        CoreAPB3_0_APBmslave5_PSELx), .B(CoreAPB3_m4_8_0), .C(
        \CoreAPB3_0_APBmslave2_PRDATA_m[20] ), .D(N_245), .Y(
        FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_16));
    CFG4 #( .INIT(16'hF0F8) )  \PRDATA_0_iv[8]  (.A(
        CoreAPB3_0_APBmslave5_PSELx), .B(CoreAPB3_m4_6_0_0), .C(
        \CoreAPB3_0_APBmslave2_PRDATA_m[8] ), .D(N_245), .Y(
        FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_4));
    CFG4 #( .INIT(16'h0A0C) )  \PRDATA_0_iv_RNO[17]  (.A(GPOUT_reg[17])
        , .B(INTR_reg[17]), .C(CoreAPB3_0_APBmslave2_PADDR_2), .D(
        CoreAPB3_0_APBmslave2_PADDR_3), .Y(CoreAPB3_m4_7_0));
    CFG4 #( .INIT(16'hF0F8) )  \PRDATA_0_iv[24]  (.A(
        CoreAPB3_0_APBmslave5_PSELx), .B(CoreAPB3_m4_1_0), .C(
        \CoreAPB3_0_APBmslave2_PRDATA_m[24] ), .D(N_245), .Y(
        FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_20));
    CFG4 #( .INIT(16'h3353) )  PRDATA_m2 (.A(lsram_width32_PRDATA_1), 
        .B(PRDATA_reg_1), .C(CoreAPB3_0_APBmslave2_PENABLE), .D(
        CoreAPB3_0_APBmslave2_PWRITE), .Y(PRDATA_m2_net_1));
    CFG4 #( .INIT(16'hC840) )  \PRDATA_0_iv_RNO_0[30]  (.A(PRDATA4_out)
        , .B(iPRDATA29), .C(PRDATA_reg_27), .D(lsram_width32_PRDATA_27)
        , .Y(\CoreAPB3_0_APBmslave2_PRDATA_m[30] ));
    CFG4 #( .INIT(16'h0A0C) )  \PRDATA_0_iv_RNO[25]  (.A(GPOUT_reg[25])
        , .B(INTR_reg[25]), .C(CoreAPB3_0_APBmslave2_PADDR_2), .D(
        CoreAPB3_0_APBmslave2_PADDR_3), .Y(CoreAPB3_m4_4_0_0));
    CFG4 #( .INIT(16'hC840) )  \PRDATA_0_iv_RNO_0[11]  (.A(PRDATA4_out)
        , .B(iPRDATA29), .C(PRDATA_reg_8), .D(lsram_width32_PRDATA_8), 
        .Y(\CoreAPB3_0_APBmslave2_PRDATA_m[11] ));
    CFG4 #( .INIT(16'hF0F8) )  \PRDATA_0_iv[31]  (.A(
        CoreAPB3_0_APBmslave5_PSELx), .B(CoreAPB3_m4_5_0), .C(
        \CoreAPB3_0_APBmslave2_PRDATA_m[31] ), .D(N_245), .Y(
        FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_27));
    CFG4 #( .INIT(16'hF0F8) )  \PRDATA_0_iv[30]  (.A(
        CoreAPB3_0_APBmslave5_PSELx), .B(CoreAPB3_m4_0_0_0), .C(
        \CoreAPB3_0_APBmslave2_PRDATA_m[30] ), .D(N_245), .Y(
        FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_26));
    CFG4 #( .INIT(16'hF0F8) )  \PRDATA_0_iv[23]  (.A(
        CoreAPB3_0_APBmslave5_PSELx), .B(CoreAPB3_m4_0_0), .C(
        \CoreAPB3_0_APBmslave2_PRDATA_m[23] ), .D(N_245), .Y(
        FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_19));
    CFG4 #( .INIT(16'h0A0C) )  \PRDATA_0_iv_RNO[21]  (.A(GPOUT_reg[21])
        , .B(INTR_reg[21]), .C(CoreAPB3_0_APBmslave2_PADDR_2), .D(
        CoreAPB3_0_APBmslave2_PADDR_3), .Y(CoreAPB3_m4_5_0_0));
    CFG4 #( .INIT(16'hD5C0) )  \PRDATA_0_iv_1_0[7]  (.A(
        \PRDATA_0_iv_1_0_RNO[7]_net_1 ), .B(
        CoreAPB3_0_APBmslave3_PRDATA_3), .C(
        CoreAPB3_0_APBmslave3_PSELx), .D(iPRDATA29), .Y(
        \PRDATA_0_iv_1_0[7]_net_1 ));
    CFG4 #( .INIT(16'hF0F8) )  \PRDATA_0_iv[25]  (.A(
        CoreAPB3_0_APBmslave5_PSELx), .B(CoreAPB3_m4_4_0_0), .C(
        \CoreAPB3_0_APBmslave2_PRDATA_m[25] ), .D(N_245), .Y(
        FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_21));
    CFG4 #( .INIT(16'hC840) )  \PRDATA_0_iv_RNO_0[21]  (.A(PRDATA4_out)
        , .B(iPRDATA29), .C(PRDATA_reg_18), .D(lsram_width32_PRDATA_18)
        , .Y(\CoreAPB3_0_APBmslave2_PRDATA_m[21] ));
    CFG4 #( .INIT(16'hF0F8) )  \PRDATA_0_iv[27]  (.A(
        CoreAPB3_0_APBmslave5_PSELx), .B(CoreAPB3_m4_3_0), .C(
        \CoreAPB3_0_APBmslave2_PRDATA_m[27] ), .D(N_245), .Y(
        FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_23));
    CFG4 #( .INIT(16'h0A0C) )  \PRDATA_0_iv_RNO[23]  (.A(GPOUT_reg[23])
        , .B(INTR_reg[23]), .C(CoreAPB3_0_APBmslave2_PADDR_2), .D(
        CoreAPB3_0_APBmslave2_PADDR_3), .Y(CoreAPB3_m4_0_0));
    CFG4 #( .INIT(16'h0A0C) )  \PRDATA_0_iv_RNO[24]  (.A(GPOUT_reg[24])
        , .B(INTR_reg[24]), .C(CoreAPB3_0_APBmslave2_PADDR_2), .D(
        CoreAPB3_0_APBmslave2_PADDR_3), .Y(CoreAPB3_m4_1_0));
    CFG4 #( .INIT(16'h0A0C) )  \PRDATA_0_iv_RNO[29]  (.A(GPOUT_reg[29])
        , .B(INTR_reg[29]), .C(CoreAPB3_0_APBmslave2_PADDR_2), .D(
        CoreAPB3_0_APBmslave2_PADDR_3), .Y(CoreAPB3_m4_0));
    CFG4 #( .INIT(16'h0A0C) )  \PRDATA_0_iv_RNO[15]  (.A(GPOUT_reg[15])
        , .B(INTR_reg[15]), .C(CoreAPB3_0_APBmslave2_PADDR_2), .D(
        CoreAPB3_0_APBmslave2_PADDR_3), .Y(CoreAPB3_m4_11_0));
    CFG4 #( .INIT(16'h3353) )  \PRDATA_0_iv_1_0_RNO[7]  (.A(
        lsram_width32_PRDATA_4), .B(PRDATA_reg_4), .C(
        CoreAPB3_0_APBmslave2_PENABLE), .D(
        CoreAPB3_0_APBmslave2_PWRITE), .Y(
        \PRDATA_0_iv_1_0_RNO[7]_net_1 ));
    CFG4 #( .INIT(16'h3353) )  PRDATA_m2_1 (.A(lsram_width32_PRDATA_3), 
        .B(PRDATA_reg_3), .C(CoreAPB3_0_APBmslave2_PENABLE), .D(
        CoreAPB3_0_APBmslave2_PWRITE), .Y(PRDATA_m2_1_net_1));
    CFG4 #( .INIT(16'h0A0C) )  \PRDATA_0_iv_RNO[11]  (.A(GPOUT_reg[11])
        , .B(INTR_reg[11]), .C(CoreAPB3_0_APBmslave2_PADDR_2), .D(
        CoreAPB3_0_APBmslave2_PADDR_3), .Y(CoreAPB3_m4_3_0_0));
    
endmodule


module CoreAPB3_Z1(
       FIC_MSS_0_FIC_0_APB_MASTER_PADDR,
       iPSELS_2,
       \CONFIG_reg[3] ,
       \CONFIG_reg[5] ,
       \CONFIG_reg[6] ,
       \CONFIG_reg[2] ,
       \CONFIG_reg[1] ,
       \CONFIG_reg[0] ,
       CoreAPB3_0_APBmslave3_PRDATA,
       PRDATA_reg,
       lsram_width32_PRDATA,
       CoreAPB3_0_APBmslave2_PADDR_5,
       CoreAPB3_0_APBmslave2_PADDR_2,
       CoreAPB3_0_APBmslave2_PADDR_1,
       CoreAPB3_0_APBmslave2_PADDR_0,
       CoreAPB3_0_APBmslave2_PADDR_3,
       gpin3_3,
       gpin3_5,
       gpin3_6,
       gpin3_2,
       gpin3_1,
       gpin3_0,
       GPOUT_reg_4,
       GPOUT_reg_0,
       GPOUT_reg_6,
       GPOUT_reg_5,
       GPOUT_reg_1,
       GPOUT_reg_2,
       GPOUT_reg_8,
       GPOUT_reg_9,
       GPOUT_reg_10,
       GPOUT_reg_11,
       GPOUT_reg_12,
       GPOUT_reg_13,
       GPOUT_reg_14,
       GPOUT_reg_15,
       GPOUT_reg_16,
       GPOUT_reg_17,
       GPOUT_reg_18,
       GPOUT_reg_19,
       GPOUT_reg_20,
       GPOUT_reg_21,
       GPOUT_reg_22,
       GPOUT_reg_23,
       GPOUT_reg_24,
       GPOUT_reg_25,
       GPOUT_reg_26,
       GPOUT_reg_27,
       GPOUT_reg_28,
       GPOUT_reg_29,
       GPOUT_reg_30,
       GPOUT_reg_31,
       INTR_reg_2,
       INTR_reg_1,
       INTR_reg_5,
       INTR_reg_6,
       INTR_reg_0,
       INTR_reg_4,
       INTR_reg_7,
       INTR_reg_8,
       INTR_reg_9,
       INTR_reg_10,
       INTR_reg_11,
       INTR_reg_12,
       INTR_reg_13,
       INTR_reg_14,
       INTR_reg_15,
       INTR_reg_16,
       INTR_reg_17,
       INTR_reg_18,
       INTR_reg_19,
       INTR_reg_20,
       INTR_reg_21,
       INTR_reg_22,
       INTR_reg_23,
       INTR_reg_24,
       INTR_reg_25,
       INTR_reg_26,
       INTR_reg_27,
       INTR_reg_28,
       INTR_reg_29,
       INTR_reg_30,
       INTR_reg_31,
       FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_0,
       FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_5,
       FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_10,
       FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_19,
       FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_20,
       FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_6,
       FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_17,
       FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_18,
       FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_7,
       FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_15,
       FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_16,
       FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_8,
       FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_13,
       FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_14,
       FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_9,
       FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_11,
       FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_12,
       FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_21,
       FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_22,
       FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_23,
       FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_24,
       FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_25,
       FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_26,
       FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_27,
       FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_28,
       FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_1,
       FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_4,
       iPRDATA29,
       FIC_MSS_0_FIC_0_APB_MASTER_PSELx,
       CoreAPB3_0_APBmslave5_PSELx,
       N_245,
       N_603,
       PRDATA_N_3_0,
       CoreAPB3_0_APBmslave3_PSELx,
       CoreAPB3_N_8_3_i_0,
       N_247,
       CoreAPB3_N_8_2_i_0,
       CoreAPB3_N_8_1_i_0,
       CoreAPB3_N_8_i_0,
       N_4755,
       N_4731,
       N_4699,
       N_4675,
       N_4875,
       N_4851,
       N_4819,
       N_4795,
       N_4761,
       N_4737,
       N_4705,
       N_4681,
       N_4881,
       N_4857,
       N_4825,
       N_4801,
       N_4760,
       N_4736,
       N_4704,
       N_4680,
       N_4880,
       N_4856,
       N_4824,
       N_4800,
       N_4756,
       N_4732,
       N_4700,
       N_4676,
       N_4876,
       N_4852,
       N_4820,
       N_4796,
       N_4757,
       N_4733,
       N_4701,
       N_4677,
       N_4877,
       N_4853,
       N_4821,
       N_4797,
       N_4759,
       N_4735,
       N_4703,
       N_4679,
       N_4879,
       N_4855,
       N_4823,
       N_4799,
       N_4758,
       N_4734,
       N_4702,
       N_4678,
       N_4878,
       N_4854,
       N_4822,
       N_4798,
       CoreAPB3_0_APBmslave2_PENABLE,
       CoreAPB3_0_APBmslave2_PWRITE,
       N_610,
       PRDATA4_out,
       CoreAPB3_N_8_0_i_0,
       N_4762,
       N_4738,
       N_4706,
       N_4682,
       N_4882,
       N_4858,
       N_4826,
       N_4802,
       PRDATA_m1_e_1,
       CoreAPB3_0_APBmslave3_PREADY,
       CoreAPB3_0_APBmslave2_PREADY,
       PREADY_0_iv_i_0,
       \CONFIG_reg[4]2_0_a4_0_a2_0_RNIBB9M2 ,
       N_452
    );
input  [31:28] FIC_MSS_0_FIC_0_APB_MASTER_PADDR;
output [5:5] iPSELS_2;
input  [1:1] \CONFIG_reg[3] ;
input  [1:1] \CONFIG_reg[5] ;
input  [1:1] \CONFIG_reg[6] ;
input  [1:1] \CONFIG_reg[2] ;
input  [1:1] \CONFIG_reg[1] ;
input  [1:1] \CONFIG_reg[0] ;
input  [7:0] CoreAPB3_0_APBmslave3_PRDATA;
input  [31:0] PRDATA_reg;
input  [31:0] lsram_width32_PRDATA;
input  CoreAPB3_0_APBmslave2_PADDR_5;
input  CoreAPB3_0_APBmslave2_PADDR_2;
input  CoreAPB3_0_APBmslave2_PADDR_1;
input  CoreAPB3_0_APBmslave2_PADDR_0;
input  CoreAPB3_0_APBmslave2_PADDR_3;
input  gpin3_3;
input  gpin3_5;
input  gpin3_6;
input  gpin3_2;
input  gpin3_1;
input  gpin3_0;
input  GPOUT_reg_4;
input  GPOUT_reg_0;
input  GPOUT_reg_6;
input  GPOUT_reg_5;
input  GPOUT_reg_1;
input  GPOUT_reg_2;
input  GPOUT_reg_8;
input  GPOUT_reg_9;
input  GPOUT_reg_10;
input  GPOUT_reg_11;
input  GPOUT_reg_12;
input  GPOUT_reg_13;
input  GPOUT_reg_14;
input  GPOUT_reg_15;
input  GPOUT_reg_16;
input  GPOUT_reg_17;
input  GPOUT_reg_18;
input  GPOUT_reg_19;
input  GPOUT_reg_20;
input  GPOUT_reg_21;
input  GPOUT_reg_22;
input  GPOUT_reg_23;
input  GPOUT_reg_24;
input  GPOUT_reg_25;
input  GPOUT_reg_26;
input  GPOUT_reg_27;
input  GPOUT_reg_28;
input  GPOUT_reg_29;
input  GPOUT_reg_30;
input  GPOUT_reg_31;
input  INTR_reg_2;
input  INTR_reg_1;
input  INTR_reg_5;
input  INTR_reg_6;
input  INTR_reg_0;
input  INTR_reg_4;
input  INTR_reg_7;
input  INTR_reg_8;
input  INTR_reg_9;
input  INTR_reg_10;
input  INTR_reg_11;
input  INTR_reg_12;
input  INTR_reg_13;
input  INTR_reg_14;
input  INTR_reg_15;
input  INTR_reg_16;
input  INTR_reg_17;
input  INTR_reg_18;
input  INTR_reg_19;
input  INTR_reg_20;
input  INTR_reg_21;
input  INTR_reg_22;
input  INTR_reg_23;
input  INTR_reg_24;
input  INTR_reg_25;
input  INTR_reg_26;
input  INTR_reg_27;
input  INTR_reg_28;
input  INTR_reg_29;
input  INTR_reg_30;
input  INTR_reg_31;
output FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_0;
output FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_5;
output FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_10;
output FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_19;
output FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_20;
output FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_6;
output FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_17;
output FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_18;
output FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_7;
output FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_15;
output FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_16;
output FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_8;
output FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_13;
output FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_14;
output FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_9;
output FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_11;
output FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_12;
output FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_21;
output FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_22;
output FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_23;
output FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_24;
output FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_25;
output FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_26;
output FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_27;
output FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_28;
output FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_1;
output FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_4;
output iPRDATA29;
input  FIC_MSS_0_FIC_0_APB_MASTER_PSELx;
output CoreAPB3_0_APBmslave5_PSELx;
input  N_245;
input  N_603;
input  PRDATA_N_3_0;
output CoreAPB3_0_APBmslave3_PSELx;
output CoreAPB3_N_8_3_i_0;
input  N_247;
output CoreAPB3_N_8_2_i_0;
output CoreAPB3_N_8_1_i_0;
output CoreAPB3_N_8_i_0;
input  N_4755;
input  N_4731;
input  N_4699;
input  N_4675;
input  N_4875;
input  N_4851;
input  N_4819;
input  N_4795;
input  N_4761;
input  N_4737;
input  N_4705;
input  N_4681;
input  N_4881;
input  N_4857;
input  N_4825;
input  N_4801;
input  N_4760;
input  N_4736;
input  N_4704;
input  N_4680;
input  N_4880;
input  N_4856;
input  N_4824;
input  N_4800;
input  N_4756;
input  N_4732;
input  N_4700;
input  N_4676;
input  N_4876;
input  N_4852;
input  N_4820;
input  N_4796;
input  N_4757;
input  N_4733;
input  N_4701;
input  N_4677;
input  N_4877;
input  N_4853;
input  N_4821;
input  N_4797;
input  N_4759;
input  N_4735;
input  N_4703;
input  N_4679;
input  N_4879;
input  N_4855;
input  N_4823;
input  N_4799;
input  N_4758;
input  N_4734;
input  N_4702;
input  N_4678;
input  N_4878;
input  N_4854;
input  N_4822;
input  N_4798;
input  CoreAPB3_0_APBmslave2_PENABLE;
input  CoreAPB3_0_APBmslave2_PWRITE;
input  N_610;
input  PRDATA4_out;
output CoreAPB3_N_8_0_i_0;
input  N_4762;
input  N_4738;
input  N_4706;
input  N_4682;
input  N_4882;
input  N_4858;
input  N_4826;
input  N_4802;
input  PRDATA_m1_e_1;
input  CoreAPB3_0_APBmslave3_PREADY;
input  CoreAPB3_0_APBmslave2_PREADY;
output PREADY_0_iv_i_0;
input  \CONFIG_reg[4]2_0_a4_0_a2_0_RNIBB9M2 ;
input  N_452;

    wire \iPSELS_sx[2]_net_1 , g0_0_0, g0_0_net_1, g2_3_net_1, 
        g0_2_3_net_1, g2_4_net_1, CoreAPB3_m8_0, r_N_4_0_0, 
        \CoreAPB3_0_APBmslave5_PRDATA_m_c_0[3] , PRDATA_N_8_mux_0, 
        g0_4_1, CoreAPB3_m6_ns_net_1, CoreAPB3_m7_3_1, 
        CoreAPB3_N_8_3_i_1_net_1, CoreAPB3_N_3_i_0_li_3, 
        \CoreAPB3_0_APBmslave5_PRDATA_m_d_a0[2]_net_1 , 
        CoreAPB3_m7_2_1, CoreAPB3_N_8_2_i_1_net_1, 
        CoreAPB3_N_3_i_0_li_2, 
        \CoreAPB3_0_APBmslave5_PRDATA_m_d_a0[1]_net_1 , 
        CoreAPB3_m7_1_1, CoreAPB3_N_8_1_i_1_net_1, 
        CoreAPB3_N_3_i_0_li_1, 
        \CoreAPB3_0_APBmslave5_PRDATA_m_d_a0[5]_net_1 , 
        \CoreAPB3_0_APBmslave5_PRDATA_m_d_a0[6]_net_1 , 
        CoreAPB3_N_8_0_i_1_net_1, CoreAPB3_m7_1, 
        CoreAPB3_N_8_i_1_net_1, CoreAPB3_N_3_i_0_li, 
        \CoreAPB3_0_APBmslave5_PRDATA_m_d_a0[0]_net_1 , 
        CoreAPB3_m2_0_am_1, CoreAPB3_m2_0_am_net_1, CoreAPB3_m2_0_bm_1, 
        CoreAPB3_m2_0_bm_net_1, CoreAPB3_m2_2_am_1_1_net_1, 
        CoreAPB3_m2_2_am_net_1, CoreAPB3_m2_2_bm_1_1_net_1, 
        CoreAPB3_m2_2_bm_net_1, CoreAPB3_m2_4_am_1_1_net_1, 
        CoreAPB3_m2_4_am_net_1, CoreAPB3_m2_4_bm_1_1_net_1, 
        CoreAPB3_m2_4_bm_net_1, CoreAPB3_m2_6_am_1_1_net_1, 
        CoreAPB3_m2_6_am_net_1, CoreAPB3_m2_6_bm_1_1_net_1, 
        CoreAPB3_m2_6_bm_net_1, CoreAPB3_m2_8_am_1_1_net_1, 
        CoreAPB3_m2_8_am_net_1, CoreAPB3_m2_8_bm_1_1_net_1, 
        CoreAPB3_m2_8_bm_net_1, CoreAPB3_m6_0_am_1, 
        CoreAPB3_m6_0_am_net_1, CoreAPB3_m6_0_bm_1, 
        CoreAPB3_m6_0_bm_net_1, CoreAPB3_m2_14_1, CoreAPB3_N_3_9, 
        CoreAPB3_m5_1, CoreAPB3_N_6_4, CoreAPB3_N_3_i_0_li_0, 
        CoreAPB3_m6_0_ns_net_1, \iPSELS_1[3] , 
        CoreAPB3_m2_0_a2_3_1_net_1, CoreAPB3_m2_0_a2_1_1_net_1, 
        CoreAPB3_m2_0_a2_7_1_net_1, CoreAPB3_m2_0_a2_5_1_net_1, 
        CoreAPB3_m2_0_a2_1, 
        \CoreAPB3_0_APBmslave5_PRDATA_m_d_0[4]_net_1 , 
        CoreAPB3_m2_12_net_1, CoreAPB3_m2_11_net_1, 
        CoreAPB3_m2_10_net_1, CoreAPB3_m2_9_net_1, CoreAPB3_m7_2_0, 
        CoreAPB3_m7_0, CoreAPB3_m7_1_0, CoreAPB3_m7_3_0, GND_net_1, 
        VCC_net_1;
    
    CFG4 #( .INIT(16'h4657) )  CoreAPB3_m2_0_bm_1_1 (.A(
        CoreAPB3_0_APBmslave2_PADDR_2), .B(
        CoreAPB3_0_APBmslave2_PADDR_1), .C(N_4819), .D(N_4795), .Y(
        CoreAPB3_m2_0_bm_1));
    CFG4 #( .INIT(16'h3353) )  CoreAPB3_m2_10 (.A(
        lsram_width32_PRDATA[2]), .B(PRDATA_reg[2]), .C(
        CoreAPB3_0_APBmslave2_PENABLE), .D(
        CoreAPB3_0_APBmslave2_PWRITE), .Y(CoreAPB3_m2_10_net_1));
    CFG4 #( .INIT(16'h0080) )  CoreAPB3_m2_0_a2_5_1 (.A(
        \CONFIG_reg[1] [1]), .B(gpin3_1), .C(
        CoreAPB3_0_APBmslave2_PADDR_2), .D(
        CoreAPB3_0_APBmslave2_PADDR_3), .Y(CoreAPB3_m2_0_a2_5_1_net_1));
    CFG4 #( .INIT(16'h0800) )  
        \CoreAPB3_0_APBmslave5_PRDATA_m_d_a0[1]  (.A(N_610), .B(
        GPOUT_reg_1), .C(N_245), .D(CoreAPB3_0_APBmslave5_PSELx), .Y(
        \CoreAPB3_0_APBmslave5_PRDATA_m_d_a0[1]_net_1 ));
    CFG3 #( .INIT(8'hE2) )  CoreAPB3_m2_4_ns (.A(
        CoreAPB3_m2_4_am_net_1), .B(CoreAPB3_0_APBmslave2_PADDR_0), .C(
        CoreAPB3_m2_4_bm_net_1), .Y(CoreAPB3_N_3_i_0_li_1));
    CFG4 #( .INIT(16'h4657) )  CoreAPB3_m2_4_am_1_1 (.A(
        CoreAPB3_0_APBmslave2_PADDR_2), .B(
        CoreAPB3_0_APBmslave2_PADDR_1), .C(N_4704), .D(N_4680), .Y(
        CoreAPB3_m2_4_am_1_1_net_1));
    CFG4 #( .INIT(16'h0080) )  CoreAPB3_m2_0_a2_3_1 (.A(
        \CONFIG_reg[5] [1]), .B(gpin3_5), .C(
        CoreAPB3_0_APBmslave2_PADDR_2), .D(
        CoreAPB3_0_APBmslave2_PADDR_3), .Y(CoreAPB3_m2_0_a2_3_1_net_1));
    CFG4 #( .INIT(16'h00AC) )  \CoreAPB3_0_APBmslave5_PRDATA_m_d_0[4]  
        (.A(GPOUT_reg_4), .B(INTR_reg_4), .C(
        CoreAPB3_0_APBmslave2_PADDR_3), .D(
        CoreAPB3_0_APBmslave2_PADDR_2), .Y(
        \CoreAPB3_0_APBmslave5_PRDATA_m_d_0[4]_net_1 ));
    CFG2 #( .INIT(4'h8) )  g0_0 (.A(gpin3_3), .B(\CONFIG_reg[3] [1]), 
        .Y(g0_0_net_1));
    CFG4 #( .INIT(16'h0800) )  
        \CoreAPB3_0_APBmslave5_PRDATA_m_d_a0[5]  (.A(N_610), .B(
        GPOUT_reg_5), .C(N_245), .D(CoreAPB3_0_APBmslave5_PSELx), .Y(
        \CoreAPB3_0_APBmslave5_PRDATA_m_d_a0[5]_net_1 ));
    CFG4 #( .INIT(16'h0002) )  g0_1 (.A(CoreAPB3_0_APBmslave5_PSELx), 
        .B(N_245), .C(CoreAPB3_0_APBmslave2_PADDR_2), .D(PRDATA_N_3_0), 
        .Y(\CoreAPB3_0_APBmslave5_PRDATA_m_c_0[3] ));
    CFG4 #( .INIT(16'h34F4) )  CoreAPB3_m6_0_bm (.A(N_4879), .B(
        CoreAPB3_0_APBmslave2_PADDR_1), .C(CoreAPB3_m6_0_bm_1), .D(
        N_4855), .Y(CoreAPB3_m6_0_bm_net_1));
    CFG4 #( .INIT(16'h34F4) )  CoreAPB3_m2_14 (.A(N_4758), .B(
        CoreAPB3_0_APBmslave2_PADDR_1), .C(CoreAPB3_m2_14_1), .D(
        N_4734), .Y(CoreAPB3_N_3_9));
    CFG4 #( .INIT(16'h0F07) )  CoreAPB3_N_8_1_i_1 (.A(INTR_reg_5), .B(
        CoreAPB3_0_APBmslave5_PSELx), .C(
        \CoreAPB3_0_APBmslave5_PRDATA_m_d_a0[5]_net_1 ), .D(N_247), .Y(
        CoreAPB3_N_8_1_i_1_net_1));
    CFG3 #( .INIT(8'hE2) )  CoreAPB3_m2_6_ns (.A(
        CoreAPB3_m2_6_am_net_1), .B(CoreAPB3_0_APBmslave2_PADDR_0), .C(
        CoreAPB3_m2_6_bm_net_1), .Y(CoreAPB3_N_3_i_0_li_2));
    CFG4 #( .INIT(16'h4657) )  CoreAPB3_m2_6_am_1_1 (.A(
        CoreAPB3_0_APBmslave2_PADDR_2), .B(
        CoreAPB3_0_APBmslave2_PADDR_1), .C(N_4700), .D(N_4676), .Y(
        CoreAPB3_m2_6_am_1_1_net_1));
    COREAPB3_MUXPTOB3 u_mux_p_to_b3 (.GPOUT_reg({GPOUT_reg_31, 
        GPOUT_reg_30, GPOUT_reg_29, GPOUT_reg_28, GPOUT_reg_27, 
        GPOUT_reg_26, GPOUT_reg_25, GPOUT_reg_24, GPOUT_reg_23, 
        GPOUT_reg_22, GPOUT_reg_21, GPOUT_reg_20, GPOUT_reg_19, 
        GPOUT_reg_18, GPOUT_reg_17, GPOUT_reg_16, GPOUT_reg_15, 
        GPOUT_reg_14, GPOUT_reg_13, GPOUT_reg_12, GPOUT_reg_11, 
        GPOUT_reg_10, GPOUT_reg_9, GPOUT_reg_8}), .INTR_reg({
        INTR_reg_31, INTR_reg_30, INTR_reg_29, INTR_reg_28, 
        INTR_reg_27, INTR_reg_26, INTR_reg_25, INTR_reg_24, 
        INTR_reg_23, INTR_reg_22, INTR_reg_21, INTR_reg_20, 
        INTR_reg_19, INTR_reg_18, INTR_reg_17, INTR_reg_16, 
        INTR_reg_15, INTR_reg_14, INTR_reg_13, INTR_reg_12, 
        INTR_reg_11, INTR_reg_10, INTR_reg_9, INTR_reg_8, INTR_reg_7}), 
        .CoreAPB3_0_APBmslave5_PRDATA_m_d_0({
        \CoreAPB3_0_APBmslave5_PRDATA_m_d_0[4]_net_1 }), 
        .CoreAPB3_0_APBmslave3_PRDATA_2(
        CoreAPB3_0_APBmslave3_PRDATA[6]), 
        .CoreAPB3_0_APBmslave3_PRDATA_3(
        CoreAPB3_0_APBmslave3_PRDATA[7]), 
        .CoreAPB3_0_APBmslave3_PRDATA_0(
        CoreAPB3_0_APBmslave3_PRDATA[4]), 
        .CoreAPB3_0_APBmslave2_PADDR_1(CoreAPB3_0_APBmslave2_PADDR_1), 
        .CoreAPB3_0_APBmslave2_PADDR_2(CoreAPB3_0_APBmslave2_PADDR_2), 
        .CoreAPB3_0_APBmslave2_PADDR_0(CoreAPB3_0_APBmslave2_PADDR_0), 
        .CoreAPB3_0_APBmslave2_PADDR_3(CoreAPB3_0_APBmslave2_PADDR_3), 
        .CoreAPB3_0_APBmslave2_PADDR_5(CoreAPB3_0_APBmslave2_PADDR_5), 
        .PRDATA_reg_4(PRDATA_reg[7]), .PRDATA_reg_0(PRDATA_reg[3]), 
        .PRDATA_reg_3(PRDATA_reg[6]), .PRDATA_reg_1(PRDATA_reg[4]), 
        .PRDATA_reg_5(PRDATA_reg[8]), .PRDATA_reg_10(PRDATA_reg[13]), 
        .PRDATA_reg_19(PRDATA_reg[22]), .PRDATA_reg_20(PRDATA_reg[23]), 
        .PRDATA_reg_6(PRDATA_reg[9]), .PRDATA_reg_17(PRDATA_reg[20]), 
        .PRDATA_reg_18(PRDATA_reg[21]), .PRDATA_reg_7(PRDATA_reg[10]), 
        .PRDATA_reg_15(PRDATA_reg[18]), .PRDATA_reg_16(PRDATA_reg[19]), 
        .PRDATA_reg_8(PRDATA_reg[11]), .PRDATA_reg_13(PRDATA_reg[16]), 
        .PRDATA_reg_14(PRDATA_reg[17]), .PRDATA_reg_9(PRDATA_reg[12]), 
        .PRDATA_reg_11(PRDATA_reg[14]), .PRDATA_reg_12(PRDATA_reg[15]), 
        .PRDATA_reg_21(PRDATA_reg[24]), .PRDATA_reg_22(PRDATA_reg[25]), 
        .PRDATA_reg_23(PRDATA_reg[26]), .PRDATA_reg_24(PRDATA_reg[27]), 
        .PRDATA_reg_25(PRDATA_reg[28]), .PRDATA_reg_26(PRDATA_reg[29]), 
        .PRDATA_reg_27(PRDATA_reg[30]), .PRDATA_reg_28(PRDATA_reg[31]), 
        .lsram_width32_PRDATA_4(lsram_width32_PRDATA[7]), 
        .lsram_width32_PRDATA_0(lsram_width32_PRDATA[3]), 
        .lsram_width32_PRDATA_3(lsram_width32_PRDATA[6]), 
        .lsram_width32_PRDATA_1(lsram_width32_PRDATA[4]), 
        .lsram_width32_PRDATA_5(lsram_width32_PRDATA[8]), 
        .lsram_width32_PRDATA_10(lsram_width32_PRDATA[13]), 
        .lsram_width32_PRDATA_19(lsram_width32_PRDATA[22]), 
        .lsram_width32_PRDATA_20(lsram_width32_PRDATA[23]), 
        .lsram_width32_PRDATA_6(lsram_width32_PRDATA[9]), 
        .lsram_width32_PRDATA_17(lsram_width32_PRDATA[20]), 
        .lsram_width32_PRDATA_18(lsram_width32_PRDATA[21]), 
        .lsram_width32_PRDATA_7(lsram_width32_PRDATA[10]), 
        .lsram_width32_PRDATA_15(lsram_width32_PRDATA[18]), 
        .lsram_width32_PRDATA_16(lsram_width32_PRDATA[19]), 
        .lsram_width32_PRDATA_8(lsram_width32_PRDATA[11]), 
        .lsram_width32_PRDATA_13(lsram_width32_PRDATA[16]), 
        .lsram_width32_PRDATA_14(lsram_width32_PRDATA[17]), 
        .lsram_width32_PRDATA_9(lsram_width32_PRDATA[12]), 
        .lsram_width32_PRDATA_11(lsram_width32_PRDATA[14]), 
        .lsram_width32_PRDATA_12(lsram_width32_PRDATA[15]), 
        .lsram_width32_PRDATA_21(lsram_width32_PRDATA[24]), 
        .lsram_width32_PRDATA_22(lsram_width32_PRDATA[25]), 
        .lsram_width32_PRDATA_23(lsram_width32_PRDATA[26]), 
        .lsram_width32_PRDATA_24(lsram_width32_PRDATA[27]), 
        .lsram_width32_PRDATA_25(lsram_width32_PRDATA[28]), 
        .lsram_width32_PRDATA_26(lsram_width32_PRDATA[29]), 
        .lsram_width32_PRDATA_27(lsram_width32_PRDATA[30]), 
        .lsram_width32_PRDATA_28(lsram_width32_PRDATA[31]), 
        .FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_4(
        FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_5), 
        .FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_9(
        FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_10), 
        .FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_18(
        FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_19), 
        .FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_19(
        FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_20), 
        .FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_5(
        FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_6), 
        .FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_16(
        FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_17), 
        .FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_17(
        FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_18), 
        .FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_6(
        FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_7), 
        .FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_14(
        FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_15), 
        .FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_15(
        FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_16), 
        .FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_7(
        FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_8), 
        .FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_12(
        FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_13), 
        .FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_13(
        FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_14), 
        .FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_8(
        FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_9), 
        .FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_10(
        FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_11), 
        .FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_11(
        FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_12), 
        .FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_20(
        FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_21), 
        .FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_21(
        FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_22), 
        .FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_22(
        FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_23), 
        .FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_23(
        FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_24), 
        .FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_24(
        FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_25), 
        .FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_25(
        FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_26), 
        .FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_26(
        FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_27), 
        .FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_27(
        FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_28), 
        .FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_0(
        FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_1), 
        .FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_3(
        FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_4), 
        .CoreAPB3_0_APBmslave2_PENABLE(CoreAPB3_0_APBmslave2_PENABLE), 
        .CoreAPB3_0_APBmslave2_PWRITE(CoreAPB3_0_APBmslave2_PWRITE), 
        .PRDATA4_out(PRDATA4_out), .iPRDATA29(iPRDATA29), 
        .PRDATA_N_8_mux_0(PRDATA_N_8_mux_0), .CoreAPB3_m8_0(
        CoreAPB3_m8_0), .CoreAPB3_N_8_0_i_1(CoreAPB3_N_8_0_i_1_net_1), 
        .CoreAPB3_N_3_i_0_li_0(CoreAPB3_N_3_i_0_li_0), 
        .CoreAPB3_N_8_0_i_0(CoreAPB3_N_8_0_i_0), .N_4762(N_4762), 
        .N_4738(N_4738), .N_4706(N_4706), .N_4682(N_4682), .N_4882(
        N_4882), .N_4858(N_4858), .N_4826(N_4826), .N_4802(N_4802), 
        .CoreAPB3_0_APBmslave3_PSELx(CoreAPB3_0_APBmslave3_PSELx), 
        .CoreAPB3_0_APBmslave5_PSELx(CoreAPB3_0_APBmslave5_PSELx), 
        .N_245(N_245), .PRDATA_m1_e_1(PRDATA_m1_e_1), 
        .CoreAPB3_m2_0_a2_1_1(CoreAPB3_m2_0_a2_1_1_net_1), .N_247(
        N_247), .CoreAPB3_0_APBmslave3_PREADY(
        CoreAPB3_0_APBmslave3_PREADY), .CoreAPB3_0_APBmslave2_PREADY(
        CoreAPB3_0_APBmslave2_PREADY), .PREADY_0_iv_i_0(
        PREADY_0_iv_i_0), .\CONFIG_reg[4]2_0_a4_0_a2_0_RNIBB9M2 (
        \CONFIG_reg[4]2_0_a4_0_a2_0_RNIBB9M2 ), .CoreAPB3_m6_0_ns(
        CoreAPB3_m6_0_ns_net_1), .N_452(N_452));
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hE2) )  CoreAPB3_m2_2_ns (.A(
        CoreAPB3_m2_2_am_net_1), .B(CoreAPB3_0_APBmslave2_PADDR_0), .C(
        CoreAPB3_m2_2_bm_net_1), .Y(CoreAPB3_N_3_i_0_li_0));
    CFG4 #( .INIT(16'h4657) )  CoreAPB3_m2_6_bm_1_1 (.A(
        CoreAPB3_0_APBmslave2_PADDR_2), .B(
        CoreAPB3_0_APBmslave2_PADDR_1), .C(N_4820), .D(N_4796), .Y(
        CoreAPB3_m2_6_bm_1_1_net_1));
    CFG4 #( .INIT(16'hFBFF) )  \iPSELS_sx[2]  (.A(
        FIC_MSS_0_FIC_0_APB_MASTER_PADDR[30]), .B(
        FIC_MSS_0_FIC_0_APB_MASTER_PSELx), .C(
        FIC_MSS_0_FIC_0_APB_MASTER_PADDR[31]), .D(
        FIC_MSS_0_FIC_0_APB_MASTER_PADDR[29]), .Y(\iPSELS_sx[2]_net_1 )
        );
    CFG4 #( .INIT(16'h2A3F) )  \iPSELS_RNIC0HC2[3]  (.A(
        CoreAPB3_m2_10_net_1), .B(CoreAPB3_0_APBmslave3_PRDATA[2]), .C(
        CoreAPB3_0_APBmslave3_PSELx), .D(iPRDATA29), .Y(
        CoreAPB3_m7_3_0));
    CFG4 #( .INIT(16'h0800) )  
        \CoreAPB3_0_APBmslave5_PRDATA_m_d_a0[6]  (.A(N_610), .B(
        GPOUT_reg_6), .C(N_245), .D(CoreAPB3_0_APBmslave5_PSELx), .Y(
        \CoreAPB3_0_APBmslave5_PRDATA_m_d_a0[6]_net_1 ));
    CFG4 #( .INIT(16'hBF3F) )  \iPSELS_RNIVREC11[3]  (.A(CoreAPB3_m8_0)
        , .B(CoreAPB3_m7_1_1), .C(CoreAPB3_N_8_1_i_1_net_1), .D(
        CoreAPB3_N_3_i_0_li_1), .Y(CoreAPB3_N_8_1_i_0));
    CFG4 #( .INIT(16'h4657) )  CoreAPB3_m5_1_2 (.A(
        CoreAPB3_0_APBmslave2_PADDR_2), .B(
        CoreAPB3_0_APBmslave2_PADDR_1), .C(N_4822), .D(N_4798), .Y(
        CoreAPB3_m5_1));
    CFG4 #( .INIT(16'hCB0B) )  CoreAPB3_m2_4_bm (.A(N_4880), .B(
        CoreAPB3_0_APBmslave2_PADDR_1), .C(CoreAPB3_m2_4_bm_1_1_net_1), 
        .D(N_4856), .Y(CoreAPB3_m2_4_bm_net_1));
    CFG4 #( .INIT(16'hBF3F) )  \iPSELS_RNI1MB511[3]  (.A(CoreAPB3_m8_0)
        , .B(CoreAPB3_m7_3_1), .C(CoreAPB3_N_8_3_i_1_net_1), .D(
        CoreAPB3_N_3_i_0_li_3), .Y(CoreAPB3_N_8_3_i_0));
    CFG4 #( .INIT(16'h0F07) )  CoreAPB3_N_8_i_1 (.A(INTR_reg_0), .B(
        CoreAPB3_0_APBmslave5_PSELx), .C(
        \CoreAPB3_0_APBmslave5_PRDATA_m_d_a0[0]_net_1 ), .D(N_247), .Y(
        CoreAPB3_N_8_i_1_net_1));
    CFG3 #( .INIT(8'hE2) )  CoreAPB3_m2_8_ns (.A(
        CoreAPB3_m2_8_am_net_1), .B(CoreAPB3_0_APBmslave2_PADDR_0), .C(
        CoreAPB3_m2_8_bm_net_1), .Y(CoreAPB3_N_3_i_0_li_3));
    CFG4 #( .INIT(16'hFFBA) )  \iPSELS_RNI61LRU[3]  (.A(g0_4_1), .B(
        CoreAPB3_m6_ns_net_1), .C(g2_4_net_1), .D(
        \CoreAPB3_0_APBmslave5_PRDATA_m_c_0[3] ), .Y(
        FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_0));
    CFG3 #( .INIT(8'hE2) )  CoreAPB3_m2_0_ns (.A(
        CoreAPB3_m2_0_am_net_1), .B(CoreAPB3_0_APBmslave2_PADDR_0), .C(
        CoreAPB3_m2_0_bm_net_1), .Y(CoreAPB3_N_3_i_0_li));
    CFG4 #( .INIT(16'h4657) )  CoreAPB3_m2_0_am_1_1 (.A(
        CoreAPB3_0_APBmslave2_PADDR_2), .B(
        CoreAPB3_0_APBmslave2_PADDR_1), .C(N_4699), .D(N_4675), .Y(
        CoreAPB3_m2_0_am_1));
    CFG4 #( .INIT(16'h0F07) )  CoreAPB3_N_8_3_i_1 (.A(INTR_reg_2), .B(
        CoreAPB3_0_APBmslave5_PSELx), .C(
        \CoreAPB3_0_APBmslave5_PRDATA_m_d_a0[2]_net_1 ), .D(N_247), .Y(
        CoreAPB3_N_8_3_i_1_net_1));
    CFG4 #( .INIT(16'h0800) )  
        \CoreAPB3_0_APBmslave5_PRDATA_m_d_a0[0]  (.A(N_610), .B(
        GPOUT_reg_0), .C(N_245), .D(CoreAPB3_0_APBmslave5_PSELx), .Y(
        \CoreAPB3_0_APBmslave5_PRDATA_m_d_a0[0]_net_1 ));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h4657) )  CoreAPB3_m6_0_am_1_1 (.A(
        CoreAPB3_0_APBmslave2_PADDR_2), .B(
        CoreAPB3_0_APBmslave2_PADDR_1), .C(N_4703), .D(N_4679), .Y(
        CoreAPB3_m6_0_am_1));
    CFG4 #( .INIT(16'hF070) )  \iPSELS_RNI9Q8N5[3]  (.A(
        CoreAPB3_0_APBmslave5_PSELx), .B(CoreAPB3_m2_0_a2_1), .C(
        CoreAPB3_m7_0), .D(N_245), .Y(CoreAPB3_m7_1));
    CFG4 #( .INIT(16'h0800) )  g2_3 (.A(
        FIC_MSS_0_FIC_0_APB_MASTER_PSELx), .B(
        FIC_MSS_0_FIC_0_APB_MASTER_PADDR[30]), .C(
        FIC_MSS_0_FIC_0_APB_MASTER_PADDR[29]), .D(
        FIC_MSS_0_FIC_0_APB_MASTER_PADDR[28]), .Y(g2_3_net_1));
    CFG3 #( .INIT(8'h04) )  g2_4 (.A(
        FIC_MSS_0_FIC_0_APB_MASTER_PADDR[31]), .B(g2_3_net_1), .C(
        CoreAPB3_0_APBmslave2_PADDR_5), .Y(g2_4_net_1));
    CFG3 #( .INIT(8'h80) )  g0_6 (.A(FIC_MSS_0_FIC_0_APB_MASTER_PSELx), 
        .B(FIC_MSS_0_FIC_0_APB_MASTER_PADDR[30]), .C(
        FIC_MSS_0_FIC_0_APB_MASTER_PADDR[28]), .Y(iPSELS_2[5]));
    CFG4 #( .INIT(16'h34F4) )  CoreAPB3_m5 (.A(N_4878), .B(
        CoreAPB3_0_APBmslave2_PADDR_1), .C(CoreAPB3_m5_1), .D(N_4854), 
        .Y(CoreAPB3_N_6_4));
    CFG4 #( .INIT(16'h2000) )  \iPSELS[3]  (.A(
        FIC_MSS_0_FIC_0_APB_MASTER_PSELx), .B(
        FIC_MSS_0_FIC_0_APB_MASTER_PADDR[30]), .C(
        FIC_MSS_0_FIC_0_APB_MASTER_PADDR[28]), .D(\iPSELS_1[3] ), .Y(
        CoreAPB3_0_APBmslave3_PSELx));
    CFG4 #( .INIT(16'h2000) )  g0 (.A(CoreAPB3_0_APBmslave5_PSELx), .B(
        N_245), .C(g0_0_net_1), .D(N_603), .Y(r_N_4_0_0));
    CFG4 #( .INIT(16'h2A3F) )  \iPSELS_RNI8SGC2[3]  (.A(
        CoreAPB3_m2_9_net_1), .B(CoreAPB3_0_APBmslave3_PRDATA[0]), .C(
        CoreAPB3_0_APBmslave3_PSELx), .D(iPRDATA29), .Y(CoreAPB3_m7_0));
    CFG3 #( .INIT(8'hD8) )  CoreAPB3_m6_ns (.A(
        CoreAPB3_0_APBmslave2_PADDR_0), .B(CoreAPB3_N_6_4), .C(
        CoreAPB3_N_3_9), .Y(CoreAPB3_m6_ns_net_1));
    CFG2 #( .INIT(4'h4) )  \iPSELS_0[2]  (.A(
        FIC_MSS_0_FIC_0_APB_MASTER_PADDR[31]), .B(
        FIC_MSS_0_FIC_0_APB_MASTER_PADDR[29]), .Y(\iPSELS_1[3] ));
    CFG4 #( .INIT(16'h2A3F) )  \iPSELS_RNII6HC2[3]  (.A(
        CoreAPB3_m2_11_net_1), .B(CoreAPB3_0_APBmslave3_PRDATA[5]), .C(
        CoreAPB3_0_APBmslave3_PSELx), .D(iPRDATA29), .Y(
        CoreAPB3_m7_1_0));
    CFG4 #( .INIT(16'hCB0B) )  CoreAPB3_m2_6_bm (.A(N_4876), .B(
        CoreAPB3_0_APBmslave2_PADDR_1), .C(CoreAPB3_m2_6_bm_1_1_net_1), 
        .D(N_4852), .Y(CoreAPB3_m2_6_bm_net_1));
    CFG4 #( .INIT(16'h4657) )  CoreAPB3_m2_4_bm_1_1 (.A(
        CoreAPB3_0_APBmslave2_PADDR_2), .B(
        CoreAPB3_0_APBmslave2_PADDR_1), .C(N_4824), .D(N_4800), .Y(
        CoreAPB3_m2_4_bm_1_1_net_1));
    CFG4 #( .INIT(16'hBF3F) )  \iPSELS_RNID7K011[3]  (.A(CoreAPB3_m8_0)
        , .B(CoreAPB3_m7_1), .C(CoreAPB3_N_8_i_1_net_1), .D(
        CoreAPB3_N_3_i_0_li), .Y(CoreAPB3_N_8_i_0));
    CFG4 #( .INIT(16'hCB0B) )  CoreAPB3_m2_8_am (.A(N_4757), .B(
        CoreAPB3_0_APBmslave2_PADDR_1), .C(CoreAPB3_m2_8_am_1_1_net_1), 
        .D(N_4733), .Y(CoreAPB3_m2_8_am_net_1));
    CFG4 #( .INIT(16'hF070) )  \iPSELS_RNI7I7M5[3]  (.A(
        CoreAPB3_0_APBmslave5_PSELx), .B(CoreAPB3_m2_0_a2_3_1_net_1), 
        .C(CoreAPB3_m7_1_0), .D(N_245), .Y(CoreAPB3_m7_1_1));
    CFG4 #( .INIT(16'hCB0B) )  CoreAPB3_m2_4_am (.A(N_4760), .B(
        CoreAPB3_0_APBmslave2_PADDR_1), .C(CoreAPB3_m2_4_am_1_1_net_1), 
        .D(N_4736), .Y(CoreAPB3_m2_4_am_net_1));
    CFG4 #( .INIT(16'hFEEE) )  \iPSELS_RNIN93E4[3]  (.A(
        PRDATA_N_8_mux_0), .B(r_N_4_0_0), .C(
        CoreAPB3_0_APBmslave3_PRDATA[3]), .D(
        CoreAPB3_0_APBmslave3_PSELx), .Y(g0_4_1));
    CFG4 #( .INIT(16'h0800) )  g0_2_3 (.A(
        FIC_MSS_0_FIC_0_APB_MASTER_PSELx), .B(
        FIC_MSS_0_FIC_0_APB_MASTER_PADDR[30]), .C(
        FIC_MSS_0_FIC_0_APB_MASTER_PADDR[29]), .D(
        FIC_MSS_0_FIC_0_APB_MASTER_PADDR[28]), .Y(g0_2_3_net_1));
    CFG2 #( .INIT(4'h1) )  \iPSELS[2]  (.A(\iPSELS_sx[2]_net_1 ), .B(
        FIC_MSS_0_FIC_0_APB_MASTER_PADDR[28]), .Y(iPRDATA29));
    CFG4 #( .INIT(16'h0080) )  CoreAPB3_m2_0_a2_7_1 (.A(
        \CONFIG_reg[2] [1]), .B(gpin3_2), .C(
        CoreAPB3_0_APBmslave2_PADDR_2), .D(
        CoreAPB3_0_APBmslave2_PADDR_3), .Y(CoreAPB3_m2_0_a2_7_1_net_1));
    CFG4 #( .INIT(16'hBF3F) )  \iPSELS_RNINUV221[3]  (.A(CoreAPB3_m8_0)
        , .B(CoreAPB3_m7_2_1), .C(CoreAPB3_N_8_2_i_1_net_1), .D(
        CoreAPB3_N_3_i_0_li_2), .Y(CoreAPB3_N_8_2_i_0));
    CFG4 #( .INIT(16'hCB0B) )  CoreAPB3_m2_0_bm (.A(N_4875), .B(
        CoreAPB3_0_APBmslave2_PADDR_1), .C(CoreAPB3_m2_0_bm_1), .D(
        N_4851), .Y(CoreAPB3_m2_0_bm_net_1));
    CFG4 #( .INIT(16'h4657) )  CoreAPB3_m2_8_bm_1_1 (.A(
        CoreAPB3_0_APBmslave2_PADDR_2), .B(
        CoreAPB3_0_APBmslave2_PADDR_1), .C(N_4821), .D(N_4797), .Y(
        CoreAPB3_m2_8_bm_1_1_net_1));
    CFG4 #( .INIT(16'hF070) )  \iPSELS_RNIF5276[3]  (.A(
        CoreAPB3_0_APBmslave5_PSELx), .B(CoreAPB3_m2_0_a2_5_1_net_1), 
        .C(CoreAPB3_m7_2_0), .D(N_245), .Y(CoreAPB3_m7_2_1));
    CFG4 #( .INIT(16'hCB0B) )  CoreAPB3_m2_8_bm (.A(N_4877), .B(
        CoreAPB3_0_APBmslave2_PADDR_1), .C(CoreAPB3_m2_8_bm_1_1_net_1), 
        .D(N_4853), .Y(CoreAPB3_m2_8_bm_net_1));
    CFG4 #( .INIT(16'h4657) )  CoreAPB3_m2_8_am_1_1 (.A(
        CoreAPB3_0_APBmslave2_PADDR_2), .B(
        CoreAPB3_0_APBmslave2_PADDR_1), .C(N_4701), .D(N_4677), .Y(
        CoreAPB3_m2_8_am_1_1_net_1));
    CFG4 #( .INIT(16'hCB0B) )  CoreAPB3_m2_0_am (.A(N_4755), .B(
        CoreAPB3_0_APBmslave2_PADDR_1), .C(CoreAPB3_m2_0_am_1), .D(
        N_4731), .Y(CoreAPB3_m2_0_am_net_1));
    CFG4 #( .INIT(16'h3353) )  CoreAPB3_m2_11 (.A(
        lsram_width32_PRDATA[5]), .B(PRDATA_reg[5]), .C(
        CoreAPB3_0_APBmslave2_PENABLE), .D(
        CoreAPB3_0_APBmslave2_PWRITE), .Y(CoreAPB3_m2_11_net_1));
    CFG4 #( .INIT(16'h0080) )  CoreAPB3_m2_0_a2_1_1 (.A(
        \CONFIG_reg[6] [1]), .B(gpin3_6), .C(
        CoreAPB3_0_APBmslave2_PADDR_2), .D(
        CoreAPB3_0_APBmslave2_PADDR_3), .Y(CoreAPB3_m2_0_a2_1_1_net_1));
    CFG4 #( .INIT(16'h4657) )  CoreAPB3_m2_2_bm_1_1 (.A(
        CoreAPB3_0_APBmslave2_PADDR_2), .B(
        CoreAPB3_0_APBmslave2_PADDR_1), .C(N_4825), .D(N_4801), .Y(
        CoreAPB3_m2_2_bm_1_1_net_1));
    CFG4 #( .INIT(16'hCB0B) )  CoreAPB3_m2_2_am (.A(N_4761), .B(
        CoreAPB3_0_APBmslave2_PADDR_1), .C(CoreAPB3_m2_2_am_1_1_net_1), 
        .D(N_4737), .Y(CoreAPB3_m2_2_am_net_1));
    CFG4 #( .INIT(16'h4657) )  CoreAPB3_m6_0_bm_1_1 (.A(
        CoreAPB3_0_APBmslave2_PADDR_2), .B(
        CoreAPB3_0_APBmslave2_PADDR_1), .C(N_4823), .D(N_4799), .Y(
        CoreAPB3_m6_0_bm_1));
    CFG4 #( .INIT(16'h3353) )  CoreAPB3_m2_9 (.A(
        lsram_width32_PRDATA[0]), .B(PRDATA_reg[0]), .C(
        CoreAPB3_0_APBmslave2_PENABLE), .D(
        CoreAPB3_0_APBmslave2_PWRITE), .Y(CoreAPB3_m2_9_net_1));
    CFG4 #( .INIT(16'h0F07) )  CoreAPB3_N_8_0_i_1 (.A(INTR_reg_6), .B(
        CoreAPB3_0_APBmslave5_PSELx), .C(
        \CoreAPB3_0_APBmslave5_PRDATA_m_d_a0[6]_net_1 ), .D(N_247), .Y(
        CoreAPB3_N_8_0_i_1_net_1));
    CFG4 #( .INIT(16'h3353) )  CoreAPB3_m2_12 (.A(
        lsram_width32_PRDATA[1]), .B(PRDATA_reg[1]), .C(
        CoreAPB3_0_APBmslave2_PENABLE), .D(
        CoreAPB3_0_APBmslave2_PWRITE), .Y(CoreAPB3_m2_12_net_1));
    CFG4 #( .INIT(16'h0F07) )  CoreAPB3_N_8_2_i_1 (.A(INTR_reg_1), .B(
        CoreAPB3_0_APBmslave5_PSELx), .C(
        \CoreAPB3_0_APBmslave5_PRDATA_m_d_a0[1]_net_1 ), .D(N_247), .Y(
        CoreAPB3_N_8_2_i_1_net_1));
    CFG4 #( .INIT(16'h0080) )  CoreAPB3_m2_0_a2_1_0 (.A(
        \CONFIG_reg[0] [1]), .B(gpin3_0), .C(
        CoreAPB3_0_APBmslave2_PADDR_2), .D(
        CoreAPB3_0_APBmslave2_PADDR_3), .Y(CoreAPB3_m2_0_a2_1));
    CFG4 #( .INIT(16'h4657) )  CoreAPB3_m2_2_am_1_1 (.A(
        CoreAPB3_0_APBmslave2_PADDR_2), .B(
        CoreAPB3_0_APBmslave2_PADDR_1), .C(N_4705), .D(N_4681), .Y(
        CoreAPB3_m2_2_am_1_1_net_1));
    CFG3 #( .INIT(8'h04) )  g0_2 (.A(
        FIC_MSS_0_FIC_0_APB_MASTER_PADDR[31]), .B(g0_2_3_net_1), .C(
        CoreAPB3_0_APBmslave2_PADDR_5), .Y(CoreAPB3_m8_0));
    CFG4 #( .INIT(16'hCB0B) )  CoreAPB3_m2_6_am (.A(N_4756), .B(
        CoreAPB3_0_APBmslave2_PADDR_1), .C(CoreAPB3_m2_6_am_1_1_net_1), 
        .D(N_4732), .Y(CoreAPB3_m2_6_am_net_1));
    CFG4 #( .INIT(16'h4657) )  CoreAPB3_m2_14_1_2 (.A(
        CoreAPB3_0_APBmslave2_PADDR_2), .B(
        CoreAPB3_0_APBmslave2_PADDR_1), .C(N_4702), .D(N_4678), .Y(
        CoreAPB3_m2_14_1));
    CFG4 #( .INIT(16'h34F4) )  CoreAPB3_m6_0_am (.A(N_4759), .B(
        CoreAPB3_0_APBmslave2_PADDR_1), .C(CoreAPB3_m6_0_am_1), .D(
        N_4735), .Y(CoreAPB3_m6_0_am_net_1));
    CFG4 #( .INIT(16'h2A3F) )  \iPSELS_RNIAUGC2[3]  (.A(
        CoreAPB3_m2_12_net_1), .B(CoreAPB3_0_APBmslave3_PRDATA[1]), .C(
        CoreAPB3_0_APBmslave3_PSELx), .D(iPRDATA29), .Y(
        CoreAPB3_m7_2_0));
    CFG2 #( .INIT(4'h8) )  g0_0_1 (.A(
        FIC_MSS_0_FIC_0_APB_MASTER_PADDR[30]), .B(
        FIC_MSS_0_FIC_0_APB_MASTER_PSELx), .Y(g0_0_0));
    CFG4 #( .INIT(16'hCB0B) )  CoreAPB3_m2_2_bm (.A(N_4881), .B(
        CoreAPB3_0_APBmslave2_PADDR_1), .C(CoreAPB3_m2_2_bm_1_1_net_1), 
        .D(N_4857), .Y(CoreAPB3_m2_2_bm_net_1));
    CFG3 #( .INIT(8'hE2) )  CoreAPB3_m6_0_ns (.A(
        CoreAPB3_m6_0_am_net_1), .B(CoreAPB3_0_APBmslave2_PADDR_0), .C(
        CoreAPB3_m6_0_bm_net_1), .Y(CoreAPB3_m6_0_ns_net_1));
    CFG4 #( .INIT(16'h0800) )  
        \CoreAPB3_0_APBmslave5_PRDATA_m_d_a0[2]  (.A(N_610), .B(
        GPOUT_reg_2), .C(N_245), .D(CoreAPB3_0_APBmslave5_PSELx), .Y(
        \CoreAPB3_0_APBmslave5_PRDATA_m_d_a0[2]_net_1 ));
    CFG4 #( .INIT(16'hF070) )  \iPSELS_RNILGRM5[3]  (.A(
        CoreAPB3_0_APBmslave5_PSELx), .B(CoreAPB3_m2_0_a2_7_1_net_1), 
        .C(CoreAPB3_m7_3_0), .D(N_245), .Y(CoreAPB3_m7_3_1));
    CFG4 #( .INIT(16'h1000) )  g0_5 (.A(
        FIC_MSS_0_FIC_0_APB_MASTER_PADDR[31]), .B(
        FIC_MSS_0_FIC_0_APB_MASTER_PADDR[29]), .C(g0_0_0), .D(
        FIC_MSS_0_FIC_0_APB_MASTER_PADDR[28]), .Y(
        CoreAPB3_0_APBmslave5_PSELx));
    
endmodule


module FIC_OSC_0_OSC(
       OSC_0_RCOSC_25_50MHZ_CCC_OUT_RCOSC_25_50MHZ_CCC
    );
output OSC_0_RCOSC_25_50MHZ_CCC_OUT_RCOSC_25_50MHZ_CCC;

    wire GND_net_1, VCC_net_1;
    
    RCOSC_25_50MHZ #( .FREQUENCY(50.0) )  I_RCOSC_25_50MHZ (.CLKOUT(
        OSC_0_RCOSC_25_50MHZ_CCC_OUT_RCOSC_25_50MHZ_CCC));
    VCC VCC (.Y(VCC_net_1));
    GND GND (.Y(GND_net_1));
    
endmodule


module FIC_FCCC_0_FCCC(
       FCCC_0_GL1,
       FCCC_0_LOCK,
       OSC_0_RCOSC_25_50MHZ_CCC_OUT_RCOSC_25_50MHZ_CCC
    );
output FCCC_0_GL1;
output FCCC_0_LOCK;
input  OSC_0_RCOSC_25_50MHZ_CCC_OUT_RCOSC_25_50MHZ_CCC;

    wire GL1_net, VCC_net_1, GND_net_1;
    
    CLKINT GL1_INST (.A(GL1_net), .Y(FCCC_0_GL1));
    VCC VCC (.Y(VCC_net_1));
    GND GND (.Y(GND_net_1));
    CCC #( .INIT(210'h0000007FB8000044D64000318C6307C6318C61EC0404040400301)
        , .VCOFREQUENCY(800.0) )  CCC_INST (.Y0(), .Y1(), .Y2(), .Y3(), 
        .PRDATA({nc0, nc1, nc2, nc3, nc4, nc5, nc6, nc7}), .LOCK(
        FCCC_0_LOCK), .BUSY(), .CLK0(VCC_net_1), .CLK1(VCC_net_1), 
        .CLK2(VCC_net_1), .CLK3(VCC_net_1), .NGMUX0_SEL(GND_net_1), 
        .NGMUX1_SEL(GND_net_1), .NGMUX2_SEL(GND_net_1), .NGMUX3_SEL(
        GND_net_1), .NGMUX0_HOLD_N(VCC_net_1), .NGMUX1_HOLD_N(
        VCC_net_1), .NGMUX2_HOLD_N(VCC_net_1), .NGMUX3_HOLD_N(
        VCC_net_1), .NGMUX0_ARST_N(VCC_net_1), .NGMUX1_ARST_N(
        VCC_net_1), .NGMUX2_ARST_N(VCC_net_1), .NGMUX3_ARST_N(
        VCC_net_1), .PLL_BYPASS_N(VCC_net_1), .PLL_ARST_N(VCC_net_1), 
        .PLL_POWERDOWN_N(VCC_net_1), .GPD0_ARST_N(VCC_net_1), 
        .GPD1_ARST_N(VCC_net_1), .GPD2_ARST_N(VCC_net_1), .GPD3_ARST_N(
        VCC_net_1), .PRESET_N(GND_net_1), .PCLK(VCC_net_1), .PSEL(
        VCC_net_1), .PENABLE(VCC_net_1), .PWRITE(VCC_net_1), .PADDR({
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1}), .PWDATA({VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1}), 
        .CLK0_PAD(GND_net_1), .CLK1_PAD(GND_net_1), .CLK2_PAD(
        GND_net_1), .CLK3_PAD(GND_net_1), .GL0(), .GL1(GL1_net), .GL2()
        , .GL3(), .RCOSC_25_50MHZ(
        OSC_0_RCOSC_25_50MHZ_CCC_OUT_RCOSC_25_50MHZ_CCC), .RCOSC_1MHZ(
        GND_net_1), .XTLOSC(GND_net_1));
    
endmodule


module reg16x8(
       CoreAPB3_0_APBmslave3_PRDATA,
       CoreAPB3_0_APBmslave2_PWDATA,
       CoreAPB3_0_APBmslave2_PADDR,
       MSS_RESET_N_F2M_c,
       FCCC_0_GL1,
       rd_enable,
       wr_enable
    );
output [7:0] CoreAPB3_0_APBmslave3_PRDATA;
input  [7:0] CoreAPB3_0_APBmslave2_PWDATA;
input  [3:0] CoreAPB3_0_APBmslave2_PADDR;
input  MSS_RESET_N_F2M_c;
input  FCCC_0_GL1;
input  rd_enable;
input  wr_enable;

    wire un1_mem_0_5_122_net_1, un1_mem_0_5_122_i, 
        un1_mem_0_5_26_net_1, un1_mem_0_5_26_i, un1_mem_0_5_10_net_1, 
        un1_mem_0_5_10_i, un1_mem_0_5_80_net_1, un1_mem_0_5_80_i, 
        un1_mem_0_5_28_net_1, un1_mem_0_5_28_i, un1_mem_0_5_12_net_1, 
        un1_mem_0_5_12_i, un1_mem_0_5_81_net_1, un1_mem_0_5_81_i, 
        un1_mem_0_5_57_net_1, un1_mem_0_5_57_i, un1_mem_0_5_112_net_1, 
        un1_mem_0_5_112_i, un1_mem_0_5_104_net_1, un1_mem_0_5_104_i, 
        un1_mem_0_5_16_net_1, un1_mem_0_5_16_i, un1_mem_0_5_88_net_1, 
        un1_mem_0_5_88_i, un1_mem_0_5_97_net_1, un1_mem_0_5_97_i, 
        un1_mem_0_5_72_net_1, un1_mem_0_5_72_i, un1_mem_0_5_7_net_1, 
        un1_mem_0_5_7_i, un1_mem_0_5_125_net_1, un1_mem_0_5_125_i, 
        un1_mem_0_5_29_net_1, un1_mem_0_5_29_i, un1_mem_0_5_13_net_1, 
        un1_mem_0_5_13_i, un1_mem_0_5_net_1, un1_mem_0_5_i, 
        un1_mem_0_5_14_net_1, un1_mem_0_5_14_i, un1_mem_0_5_82_net_1, 
        un1_mem_0_5_82_i, un1_mem_0_5_59_net_1, un1_mem_0_5_59_i, 
        un1_mem_0_5_113_net_1, un1_mem_0_5_113_i, 
        un1_mem_0_5_105_net_1, un1_mem_0_5_105_i, un1_mem_0_5_17_net_1, 
        un1_mem_0_5_17_i, un1_mem_0_5_89_net_1, un1_mem_0_5_89_i, 
        un1_mem_0_5_98_net_1, un1_mem_0_5_98_i, un1_mem_0_5_73_net_1, 
        un1_mem_0_5_73_i, un1_mem_0_5_5_net_1, un1_mem_0_5_5_i, 
        un1_mem_0_5_127_net_1, un1_mem_0_5_127_i, un1_mem_0_5_31_net_1, 
        un1_mem_0_5_31_i, un1_mem_0_5_15_net_1, un1_mem_0_5_15_i, 
        un1_mem_0_5_2_net_1, un1_mem_0_5_2_i, un1_mem_0_5_124_net_1, 
        un1_mem_0_5_124_i, un1_mem_0_5_84_net_1, un1_mem_0_5_84_i, 
        un1_mem_0_5_56_net_1, un1_mem_0_5_56_i, un1_mem_0_5_114_net_1, 
        un1_mem_0_5_114_i, un1_mem_0_5_106_net_1, un1_mem_0_5_106_i, 
        un1_mem_0_5_18_net_1, un1_mem_0_5_18_i, un1_mem_0_5_90_net_1, 
        un1_mem_0_5_90_i, un1_mem_0_5_99_net_1, un1_mem_0_5_99_i, 
        un1_mem_0_5_74_net_1, un1_mem_0_5_74_i, un1_mem_0_5_64_net_1, 
        un1_mem_0_5_64_i, un1_mem_0_5_49_net_1, un1_mem_0_5_49_i, 
        un1_mem_0_5_33_net_1, un1_mem_0_5_33_i, un1_mem_0_5_40_net_1, 
        un1_mem_0_5_40_i, un1_mem_0_5_4_net_1, un1_mem_0_5_4_i, 
        un1_mem_0_5_126_net_1, un1_mem_0_5_126_i, un1_mem_0_5_30_net_1, 
        un1_mem_0_5_30_i, un1_mem_0_5_61_net_1, un1_mem_0_5_61_i, 
        un1_mem_0_5_115_net_1, un1_mem_0_5_115_i, 
        un1_mem_0_5_107_net_1, un1_mem_0_5_107_i, un1_mem_0_5_19_net_1, 
        un1_mem_0_5_19_i, un1_mem_0_5_91_net_1, un1_mem_0_5_91_i, 
        un1_mem_0_5_96_net_1, un1_mem_0_5_96_i, un1_mem_0_5_75_net_1, 
        un1_mem_0_5_75_i, un1_mem_0_5_66_net_1, un1_mem_0_5_66_i, 
        un1_mem_0_5_51_net_1, un1_mem_0_5_51_i, un1_mem_0_5_35_net_1, 
        un1_mem_0_5_35_i, un1_mem_0_5_42_net_1, un1_mem_0_5_42_i, 
        un1_mem_0_5_6_net_1, un1_mem_0_5_6_i, un1_mem_0_5_48_net_1, 
        un1_mem_0_5_48_i, un1_mem_0_5_32_net_1, un1_mem_0_5_32_i, 
        un1_mem_0_5_43_net_1, un1_mem_0_5_43_i, un1_mem_0_5_116_net_1, 
        un1_mem_0_5_116_i, un1_mem_0_5_108_net_1, un1_mem_0_5_108_i, 
        un1_mem_0_5_20_net_1, un1_mem_0_5_20_i, un1_mem_0_5_92_net_1, 
        un1_mem_0_5_92_i, un1_mem_0_5_101_net_1, un1_mem_0_5_101_i, 
        un1_mem_0_5_76_net_1, un1_mem_0_5_76_i, un1_mem_0_5_68_net_1, 
        un1_mem_0_5_68_i, un1_mem_0_5_53_net_1, un1_mem_0_5_53_i, 
        un1_mem_0_5_37_net_1, un1_mem_0_5_37_i, un1_mem_0_5_44_net_1, 
        un1_mem_0_5_44_i, un1_mem_0_5_65_net_1, un1_mem_0_5_65_i, 
        un1_mem_0_5_50_net_1, un1_mem_0_5_50_i, un1_mem_0_5_34_net_1, 
        un1_mem_0_5_34_i, un1_mem_0_5_41_net_1, un1_mem_0_5_41_i, 
        un1_mem_0_5_85_net_1, un1_mem_0_5_85_i, un1_mem_0_5_109_net_1, 
        un1_mem_0_5_109_i, un1_mem_0_5_21_net_1, un1_mem_0_5_21_i, 
        un1_mem_0_5_93_net_1, un1_mem_0_5_93_i, un1_mem_0_5_102_net_1, 
        un1_mem_0_5_102_i, un1_mem_0_5_77_net_1, un1_mem_0_5_77_i, 
        un1_mem_0_5_69_net_1, un1_mem_0_5_69_i, un1_mem_0_5_54_net_1, 
        un1_mem_0_5_54_i, un1_mem_0_5_39_net_1, un1_mem_0_5_39_i, 
        un1_mem_0_5_46_net_1, un1_mem_0_5_46_i, un1_mem_0_5_67_net_1, 
        un1_mem_0_5_67_i, un1_mem_0_5_52_net_1, un1_mem_0_5_52_i, 
        un1_mem_0_5_36_net_1, un1_mem_0_5_36_i, un1_mem_0_5_47_net_1, 
        un1_mem_0_5_47_i, un1_mem_0_5_86_net_1, un1_mem_0_5_86_i, 
        un1_mem_0_5_58_net_1, un1_mem_0_5_58_i, un1_mem_0_5_22_net_1, 
        un1_mem_0_5_22_i, un1_mem_0_5_94_net_1, un1_mem_0_5_94_i, 
        un1_mem_0_5_103_net_1, un1_mem_0_5_103_i, un1_mem_0_5_78_net_1, 
        un1_mem_0_5_78_i, un1_mem_0_5_70_net_1, un1_mem_0_5_70_i, 
        un1_mem_0_5_3_net_1, un1_mem_0_5_3_i, un1_mem_0_5_121_net_1, 
        un1_mem_0_5_121_i, un1_mem_0_5_25_net_1, un1_mem_0_5_25_i, 
        un1_mem_0_5_9_net_1, un1_mem_0_5_9_i, un1_mem_0_5_83_net_1, 
        un1_mem_0_5_83_i, un1_mem_0_5_38_net_1, un1_mem_0_5_38_i, 
        un1_mem_0_5_45_net_1, un1_mem_0_5_45_i, un1_mem_0_5_87_net_1, 
        un1_mem_0_5_87_i, un1_mem_0_5_62_net_1, un1_mem_0_5_62_i, 
        un1_mem_0_5_117_net_1, un1_mem_0_5_117_i, un1_mem_0_5_95_net_1, 
        un1_mem_0_5_95_i, un1_mem_0_5_100_net_1, un1_mem_0_5_100_i, 
        un1_mem_0_5_79_net_1, un1_mem_0_5_79_i, un1_mem_0_5_71_net_1, 
        un1_mem_0_5_71_i, un1_mem_0_5_1_net_1, un1_mem_0_5_1_i, 
        un1_mem_0_5_123_net_1, un1_mem_0_5_123_i, un1_mem_0_5_27_net_1, 
        un1_mem_0_5_27_i, un1_mem_0_5_11_net_1, un1_mem_0_5_11_i, 
        un1_mem_0_5_55_net_1, un1_mem_0_5_55_i, un1_mem_0_5_120_net_1, 
        un1_mem_0_5_120_i, un1_mem_0_5_24_net_1, un1_mem_0_5_24_i, 
        un1_mem_0_5_8_net_1, un1_mem_0_5_8_i, un1_mem_0_5_63_net_1, 
        un1_mem_0_5_63_i, un1_mem_0_5_118_net_1, un1_mem_0_5_118_i, 
        un1_mem_0_5_110_net_1, un1_mem_0_5_110_i, un1_mem_0_5_60_net_1, 
        un1_mem_0_5_60_i, un1_mem_0_5_119_net_1, un1_mem_0_5_119_i, 
        un1_mem_0_5_111_net_1, un1_mem_0_5_111_i, un1_mem_0_5_23_net_1, 
        un1_mem_0_5_23_i, \temp_data[0]_net_1 , VCC_net_1, N_4_i_0, 
        GND_net_1, \temp_data[1]_net_1 , N_8_i_0, \temp_data[2]_net_1 , 
        N_10_i_0, \temp_data[3]_net_1 , N_12_i_0, \temp_data[4]_net_1 , 
        N_16_i_0, \temp_data[5]_net_1 , N_39_i_0, \temp_data[6]_net_1 , 
        N_47_i_0, \temp_data[7]_net_1 , N_64_i_0, 
        un1_mem_0_5_23_set_net_1, un1_mem_0_5_231_rs_net_1, 
        \mem_12_rs[7] , \mem_12_[7]_net_1 , un1_mem_0_5_231_i, 
        mem_12__1_sqmuxa, un1_mem_0_5_111_set_net_1, 
        un1_mem_0_5_239_rs_net_1, \mem_13_rs[7] , \mem_13_[7]_net_1 , 
        un1_mem_0_5_239_i, mem_13__1_sqmuxa, un1_mem_0_5_119_set_net_1, 
        un1_mem_0_5_247_rs_net_1, \mem_14_rs[7] , \mem_14_[7]_net_1 , 
        un1_mem_0_5_247_i, mem_14__1_sqmuxa, un1_mem_0_5_60_set_net_1, 
        un1_mem_0_5_252_rs_net_1, \mem_15_rs[7] , \mem_15_[7]_net_1 , 
        un1_mem_0_5_252_i, mem_15__1_sqmuxa, un1_mem_0_5_110_set_net_1, 
        un1_mem_0_5_238_rs_net_1, \mem_13_rs[6] , \mem_13_[6]_net_1 , 
        un1_mem_0_5_238_i, un1_mem_0_5_118_set_net_1, 
        un1_mem_0_5_246_rs_net_1, \mem_14_rs[6] , \mem_14_[6]_net_1 , 
        un1_mem_0_5_246_i, un1_mem_0_5_63_set_net_1, 
        un1_mem_0_5_255_rs_net_1, \mem_15_rs[6] , \mem_15_[6]_net_1 , 
        un1_mem_0_5_255_i, un1_mem_0_5_8_set_net_1, 
        un1_mem_0_5_135_rs_net_1, \mem_0_rs[7] , \mem_0_[7]_net_1 , 
        un1_mem_0_5_135_i, mem_0__1_sqmuxa, un1_mem_0_5_24_set_net_1, 
        un1_mem_0_5_143_rs_net_1, \mem_1_rs[7] , \mem_1_[7]_net_1 , 
        un1_mem_0_5_143_i, mem_1__1_sqmuxa, un1_mem_0_5_120_set_net_1, 
        un1_mem_0_5_151_rs_net_1, \mem_2_rs[7] , \mem_2_[7]_net_1 , 
        un1_mem_0_5_151_i, mem_2__1_sqmuxa, un1_mem_0_5_55_set_net_1, 
        un1_mem_0_5_160_rs_net_1, \mem_3_rs[7] , \mem_3_[7]_net_1 , 
        un1_mem_0_5_160_i, mem_3__1_sqmuxa, un1_mem_0_5_11_set_net_1, 
        un1_mem_0_5_170_rs_net_1, \mem_4_rs[7] , \mem_4_[7]_net_1 , 
        un1_mem_0_5_170_i, mem_4__1_sqmuxa, un1_mem_0_5_27_set_net_1, 
        un1_mem_0_5_186_rs_net_1, \mem_5_rs[7] , \mem_5_[7]_net_1 , 
        un1_mem_0_5_186_i, mem_5__1_sqmuxa, un1_mem_0_5_123_set_net_1, 
        un1_mem_0_5_202_rs_net_1, \mem_6_rs[7] , \mem_6_[7]_net_1 , 
        un1_mem_0_5_202_i, mem_6__1_sqmuxa, un1_mem_0_5_1_set_net_1, 
        un1_mem_0_5_217_rs_net_1, \mem_7_rs[7] , \mem_7_[7]_net_1 , 
        un1_mem_0_5_217_i, mem_7__1_sqmuxa, un1_mem_0_5_71_set_net_1, 
        un1_mem_0_5_173_rs_net_1, \mem_8_rs[7] , \mem_8_[7]_net_1 , 
        un1_mem_0_5_173_i, mem_8__1_sqmuxa, un1_mem_0_5_79_set_net_1, 
        un1_mem_0_5_189_rs_net_1, \mem_9_rs[7] , \mem_9_[7]_net_1 , 
        un1_mem_0_5_189_i, mem_9__1_sqmuxa, un1_mem_0_5_100_set_net_1, 
        un1_mem_0_5_205_rs_net_1, \mem_10_rs[7] , \mem_10_[7]_net_1 , 
        un1_mem_0_5_205_i, mem_10__1_sqmuxa, un1_mem_0_5_95_set_net_1, 
        un1_mem_0_5_220_rs_net_1, \mem_11_rs[7] , \mem_11_[7]_net_1 , 
        un1_mem_0_5_220_i, mem_11__1_sqmuxa, un1_mem_0_5_117_set_net_1, 
        un1_mem_0_5_245_rs_net_1, \mem_14_rs[5] , \mem_14_[5]_net_1 , 
        un1_mem_0_5_245_i, un1_mem_0_5_62_set_net_1, 
        un1_mem_0_5_254_rs_net_1, \mem_15_rs[5] , \mem_15_[5]_net_1 , 
        un1_mem_0_5_254_i, un1_mem_0_5_87_set_net_1, 
        un1_mem_0_5_134_rs_net_1, \mem_0_rs[6] , \mem_0_[6]_net_1 , 
        un1_mem_0_5_134_i, un1_mem_0_5_45_set_net_1, 
        un1_mem_0_5_142_rs_net_1, \mem_1_rs[6] , \mem_1_[6]_net_1 , 
        un1_mem_0_5_142_i, un1_mem_0_5_38_set_net_1, 
        un1_mem_0_5_150_rs_net_1, \mem_2_rs[6] , \mem_2_[6]_net_1 , 
        un1_mem_0_5_150_i, un1_mem_0_5_83_set_net_1, 
        un1_mem_0_5_159_rs_net_1, \mem_3_rs[6] , \mem_3_[6]_net_1 , 
        un1_mem_0_5_159_i, un1_mem_0_5_9_set_net_1, 
        un1_mem_0_5_168_rs_net_1, \mem_4_rs[6] , \mem_4_[6]_net_1 , 
        un1_mem_0_5_168_i, un1_mem_0_5_25_set_net_1, 
        un1_mem_0_5_184_rs_net_1, \mem_5_rs[6] , \mem_5_[6]_net_1 , 
        un1_mem_0_5_184_i, un1_mem_0_5_121_set_net_1, 
        un1_mem_0_5_200_rs_net_1, \mem_6_rs[6] , \mem_6_[6]_net_1 , 
        un1_mem_0_5_200_i, un1_mem_0_5_3_set_net_1, 
        un1_mem_0_5_215_rs_net_1, \mem_7_rs[6] , \mem_7_[6]_net_1 , 
        un1_mem_0_5_215_i, un1_mem_0_5_70_set_net_1, 
        un1_mem_0_5_171_rs_net_1, \mem_8_rs[6] , \mem_8_[6]_net_1 , 
        un1_mem_0_5_171_i, un1_mem_0_5_78_set_net_1, 
        un1_mem_0_5_187_rs_net_1, \mem_9_rs[6] , \mem_9_[6]_net_1 , 
        un1_mem_0_5_187_i, un1_mem_0_5_103_set_net_1, 
        un1_mem_0_5_203_rs_net_1, \mem_10_rs[6] , \mem_10_[6]_net_1 , 
        un1_mem_0_5_203_i, un1_mem_0_5_94_set_net_1, 
        un1_mem_0_5_218_rs_net_1, \mem_11_rs[6] , \mem_11_[6]_net_1 , 
        un1_mem_0_5_218_i, un1_mem_0_5_22_set_net_1, 
        un1_mem_0_5_230_rs_net_1, \mem_12_rs[6] , \mem_12_[6]_net_1 , 
        un1_mem_0_5_230_i, un1_mem_0_5_58_set_net_1, 
        un1_mem_0_5_253_rs_net_1, \mem_15_rs[4] , \mem_15_[4]_net_1 , 
        un1_mem_0_5_253_i, un1_mem_0_5_86_set_net_1, 
        un1_mem_0_5_133_rs_net_1, \mem_0_rs[5] , \mem_0_[5]_net_1 , 
        un1_mem_0_5_133_i, un1_mem_0_5_47_set_net_1, 
        un1_mem_0_5_141_rs_net_1, \mem_1_rs[5] , \mem_1_[5]_net_1 , 
        un1_mem_0_5_141_i, un1_mem_0_5_36_set_net_1, 
        un1_mem_0_5_149_rs_net_1, \mem_2_rs[5] , \mem_2_[5]_net_1 , 
        un1_mem_0_5_149_i, un1_mem_0_5_52_set_net_1, 
        un1_mem_0_5_157_rs_net_1, \mem_3_rs[5] , \mem_3_[5]_net_1 , 
        un1_mem_0_5_157_i, un1_mem_0_5_67_set_net_1, 
        un1_mem_0_5_166_rs_net_1, \mem_4_rs[5] , \mem_4_[5]_net_1 , 
        un1_mem_0_5_166_i, un1_mem_0_5_46_set_net_1, 
        un1_mem_0_5_182_rs_net_1, \mem_5_rs[5] , \mem_5_[5]_net_1 , 
        un1_mem_0_5_182_i, un1_mem_0_5_39_set_net_1, 
        un1_mem_0_5_198_rs_net_1, \mem_6_rs[5] , \mem_6_[5]_net_1 , 
        un1_mem_0_5_198_i, un1_mem_0_5_54_set_net_1, 
        un1_mem_0_5_213_rs_net_1, \mem_7_rs[5] , \mem_7_[5]_net_1 , 
        un1_mem_0_5_213_i, un1_mem_0_5_69_set_net_1, 
        un1_mem_0_5_169_rs_net_1, \mem_8_rs[5] , \mem_8_[5]_net_1 , 
        un1_mem_0_5_169_i, un1_mem_0_5_77_set_net_1, 
        un1_mem_0_5_185_rs_net_1, \mem_9_rs[5] , \mem_9_[5]_net_1 , 
        un1_mem_0_5_185_i, un1_mem_0_5_102_set_net_1, 
        un1_mem_0_5_201_rs_net_1, \mem_10_rs[5] , \mem_10_[5]_net_1 , 
        un1_mem_0_5_201_i, un1_mem_0_5_93_set_net_1, 
        un1_mem_0_5_216_rs_net_1, \mem_11_rs[5] , \mem_11_[5]_net_1 , 
        un1_mem_0_5_216_i, un1_mem_0_5_21_set_net_1, 
        un1_mem_0_5_229_rs_net_1, \mem_12_rs[5] , \mem_12_[5]_net_1 , 
        un1_mem_0_5_229_i, un1_mem_0_5_109_set_net_1, 
        un1_mem_0_5_237_rs_net_1, \mem_13_rs[5] , \mem_13_[5]_net_1 , 
        un1_mem_0_5_237_i, un1_mem_0_5_85_set_net_1, 
        un1_mem_0_5_132_rs_net_1, \mem_0_rs[4] , \mem_0_[4]_net_1 , 
        un1_mem_0_5_132_i, un1_mem_0_5_41_set_net_1, 
        un1_mem_0_5_140_rs_net_1, \mem_1_rs[4] , \mem_1_[4]_net_1 , 
        un1_mem_0_5_140_i, un1_mem_0_5_34_set_net_1, 
        un1_mem_0_5_148_rs_net_1, \mem_2_rs[4] , \mem_2_[4]_net_1 , 
        un1_mem_0_5_148_i, un1_mem_0_5_50_set_net_1, 
        un1_mem_0_5_156_rs_net_1, \mem_3_rs[4] , \mem_3_[4]_net_1 , 
        un1_mem_0_5_156_i, un1_mem_0_5_65_set_net_1, 
        un1_mem_0_5_165_rs_net_1, \mem_4_rs[4] , \mem_4_[4]_net_1 , 
        un1_mem_0_5_165_i, un1_mem_0_5_44_set_net_1, 
        un1_mem_0_5_180_rs_net_1, \mem_5_rs[4] , \mem_5_[4]_net_1 , 
        un1_mem_0_5_180_i, un1_mem_0_5_37_set_net_1, 
        un1_mem_0_5_196_rs_net_1, \mem_6_rs[4] , \mem_6_[4]_net_1 , 
        un1_mem_0_5_196_i, un1_mem_0_5_53_set_net_1, 
        un1_mem_0_5_158_rs_net_1, \mem_7_rs[4] , \mem_7_[4]_net_1 , 
        un1_mem_0_5_158_i, un1_mem_0_5_68_set_net_1, 
        un1_mem_0_5_167_rs_net_1, \mem_8_rs[4] , \mem_8_[4]_net_1 , 
        un1_mem_0_5_167_i, un1_mem_0_5_76_set_net_1, 
        un1_mem_0_5_183_rs_net_1, \mem_9_rs[4] , \mem_9_[4]_net_1 , 
        un1_mem_0_5_183_i, un1_mem_0_5_101_set_net_1, 
        un1_mem_0_5_199_rs_net_1, \mem_10_rs[4] , \mem_10_[4]_net_1 , 
        un1_mem_0_5_199_i, un1_mem_0_5_92_set_net_1, 
        un1_mem_0_5_214_rs_net_1, \mem_11_rs[4] , \mem_11_[4]_net_1 , 
        un1_mem_0_5_214_i, un1_mem_0_5_20_set_net_1, 
        un1_mem_0_5_228_rs_net_1, \mem_12_rs[4] , \mem_12_[4]_net_1 , 
        un1_mem_0_5_228_i, un1_mem_0_5_108_set_net_1, 
        un1_mem_0_5_236_rs_net_1, \mem_13_rs[4] , \mem_13_[4]_net_1 , 
        un1_mem_0_5_236_i, un1_mem_0_5_116_set_net_1, 
        un1_mem_0_5_244_rs_net_1, \mem_14_rs[4] , \mem_14_[4]_net_1 , 
        un1_mem_0_5_244_i, un1_mem_0_5_43_set_net_1, 
        un1_mem_0_5_139_rs_net_1, \mem_1_rs[3] , \mem_1_[3]_net_1 , 
        un1_mem_0_5_139_i, un1_mem_0_5_32_set_net_1, 
        un1_mem_0_5_147_rs_net_1, \mem_2_rs[3] , \mem_2_[3]_net_1 , 
        un1_mem_0_5_147_i, un1_mem_0_5_48_set_net_1, 
        un1_mem_0_5_155_rs_net_1, \mem_3_rs[3] , \mem_3_[3]_net_1 , 
        un1_mem_0_5_155_i, un1_mem_0_5_6_set_net_1, 
        un1_mem_0_5_164_rs_net_1, \mem_4_rs[3] , \mem_4_[3]_net_1 , 
        un1_mem_0_5_164_i, un1_mem_0_5_42_set_net_1, 
        un1_mem_0_5_178_rs_net_1, \mem_5_rs[3] , \mem_5_[3]_net_1 , 
        un1_mem_0_5_178_i, un1_mem_0_5_35_set_net_1, 
        un1_mem_0_5_194_rs_net_1, \mem_6_rs[3] , \mem_6_[3]_net_1 , 
        un1_mem_0_5_194_i, un1_mem_0_5_51_set_net_1, 
        un1_mem_0_5_210_rs_net_1, \mem_7_rs[3] , \mem_7_[3]_net_1 , 
        un1_mem_0_5_210_i, un1_mem_0_5_66_set_net_1, 
        un1_mem_0_5_225_rs_net_1, \mem_8_rs[3] , \mem_8_[3]_net_1 , 
        un1_mem_0_5_225_i, un1_mem_0_5_75_set_net_1, 
        un1_mem_0_5_181_rs_net_1, \mem_9_rs[3] , \mem_9_[3]_net_1 , 
        un1_mem_0_5_181_i, un1_mem_0_5_96_set_net_1, 
        un1_mem_0_5_197_rs_net_1, \mem_10_rs[3] , \mem_10_[3]_net_1 , 
        un1_mem_0_5_197_i, un1_mem_0_5_91_set_net_1, 
        un1_mem_0_5_212_rs_net_1, \mem_11_rs[3] , \mem_11_[3]_net_1 , 
        un1_mem_0_5_212_i, un1_mem_0_5_19_set_net_1, 
        un1_mem_0_5_227_rs_net_1, \mem_12_rs[3] , \mem_12_[3]_net_1 , 
        un1_mem_0_5_227_i, un1_mem_0_5_107_set_net_1, 
        un1_mem_0_5_235_rs_net_1, \mem_13_rs[3] , \mem_13_[3]_net_1 , 
        un1_mem_0_5_235_i, un1_mem_0_5_115_set_net_1, 
        un1_mem_0_5_243_rs_net_1, \mem_14_rs[3] , \mem_14_[3]_net_1 , 
        un1_mem_0_5_243_i, un1_mem_0_5_61_set_net_1, 
        un1_mem_0_5_251_rs_net_1, \mem_15_rs[3] , \mem_15_[3]_net_1 , 
        un1_mem_0_5_251_i, un1_mem_0_5_30_set_net_1, 
        un1_mem_0_5_146_rs_net_1, \mem_2_rs[2] , \mem_2_[2]_net_1 , 
        un1_mem_0_5_146_i, un1_mem_0_5_126_set_net_1, 
        un1_mem_0_5_154_rs_net_1, \mem_3_rs[2] , \mem_3_[2]_net_1 , 
        un1_mem_0_5_154_i, un1_mem_0_5_4_set_net_1, 
        un1_mem_0_5_163_rs_net_1, \mem_4_rs[2] , \mem_4_[2]_net_1 , 
        un1_mem_0_5_163_i, un1_mem_0_5_40_set_net_1, 
        un1_mem_0_5_176_rs_net_1, \mem_5_rs[2] , \mem_5_[2]_net_1 , 
        un1_mem_0_5_176_i, un1_mem_0_5_33_set_net_1, 
        un1_mem_0_5_192_rs_net_1, \mem_6_rs[2] , \mem_6_[2]_net_1 , 
        un1_mem_0_5_192_i, un1_mem_0_5_49_set_net_1, 
        un1_mem_0_5_208_rs_net_1, \mem_7_rs[2] , \mem_7_[2]_net_1 , 
        un1_mem_0_5_208_i, un1_mem_0_5_64_set_net_1, 
        un1_mem_0_5_223_rs_net_1, \mem_8_rs[2] , \mem_8_[2]_net_1 , 
        un1_mem_0_5_223_i, un1_mem_0_5_74_set_net_1, 
        un1_mem_0_5_179_rs_net_1, \mem_9_rs[2] , \mem_9_[2]_net_1 , 
        un1_mem_0_5_179_i, un1_mem_0_5_99_set_net_1, 
        un1_mem_0_5_195_rs_net_1, \mem_10_rs[2] , \mem_10_[2]_net_1 , 
        un1_mem_0_5_195_i, un1_mem_0_5_90_set_net_1, 
        un1_mem_0_5_211_rs_net_1, \mem_11_rs[2] , \mem_11_[2]_net_1 , 
        un1_mem_0_5_211_i, un1_mem_0_5_18_set_net_1, 
        un1_mem_0_5_226_rs_net_1, \mem_12_rs[2] , \mem_12_[2]_net_1 , 
        un1_mem_0_5_226_i, un1_mem_0_5_106_set_net_1, 
        un1_mem_0_5_234_rs_net_1, \mem_13_rs[2] , \mem_13_[2]_net_1 , 
        un1_mem_0_5_234_i, un1_mem_0_5_114_set_net_1, 
        un1_mem_0_5_242_rs_net_1, \mem_14_rs[2] , \mem_14_[2]_net_1 , 
        un1_mem_0_5_242_i, un1_mem_0_5_56_set_net_1, 
        un1_mem_0_5_250_rs_net_1, \mem_15_rs[2] , \mem_15_[2]_net_1 , 
        un1_mem_0_5_250_i, un1_mem_0_5_84_set_net_1, 
        un1_mem_0_5_130_rs_net_1, \mem_0_rs[3] , \mem_0_[3]_net_1 , 
        un1_mem_0_5_130_i, un1_mem_0_5_124_set_net_1, 
        un1_mem_0_5_153_rs_net_1, \mem_3_rs[1] , \mem_3_[1]_net_1 , 
        un1_mem_0_5_153_i, un1_mem_0_5_2_set_net_1, 
        un1_mem_0_5_162_rs_net_1, \mem_4_rs[1] , \mem_4_[1]_net_1 , 
        un1_mem_0_5_162_i, un1_mem_0_5_15_set_net_1, 
        un1_mem_0_5_174_rs_net_1, \mem_5_rs[1] , \mem_5_[1]_net_1 , 
        un1_mem_0_5_174_i, un1_mem_0_5_31_set_net_1, 
        un1_mem_0_5_190_rs_net_1, \mem_6_rs[1] , \mem_6_[1]_net_1 , 
        un1_mem_0_5_190_i, un1_mem_0_5_127_set_net_1, 
        un1_mem_0_5_206_rs_net_1, \mem_7_rs[1] , \mem_7_[1]_net_1 , 
        un1_mem_0_5_206_i, un1_mem_0_5_5_set_net_1, 
        un1_mem_0_5_221_rs_net_1, \mem_8_rs[1] , \mem_8_[1]_net_1 , 
        un1_mem_0_5_221_i, un1_mem_0_5_73_set_net_1, 
        un1_mem_0_5_177_rs_net_1, \mem_9_rs[1] , \mem_9_[1]_net_1 , 
        un1_mem_0_5_177_i, un1_mem_0_5_98_set_net_1, 
        un1_mem_0_5_193_rs_net_1, \mem_10_rs[1] , \mem_10_[1]_net_1 , 
        un1_mem_0_5_193_i, un1_mem_0_5_89_set_net_1, 
        un1_mem_0_5_209_rs_net_1, \mem_11_rs[1] , \mem_11_[1]_net_1 , 
        un1_mem_0_5_209_i, un1_mem_0_5_17_set_net_1, 
        un1_mem_0_5_224_rs_net_1, \mem_12_rs[1] , \mem_12_[1]_net_1 , 
        un1_mem_0_5_224_i, un1_mem_0_5_105_set_net_1, 
        un1_mem_0_5_233_rs_net_1, \mem_13_rs[1] , \mem_13_[1]_net_1 , 
        un1_mem_0_5_233_i, un1_mem_0_5_113_set_net_1, 
        un1_mem_0_5_241_rs_net_1, \mem_14_rs[1] , \mem_14_[1]_net_1 , 
        un1_mem_0_5_241_i, un1_mem_0_5_59_set_net_1, 
        un1_mem_0_5_249_rs_net_1, \mem_15_rs[1] , \mem_15_[1]_net_1 , 
        un1_mem_0_5_249_i, un1_mem_0_5_82_set_net_1, 
        un1_mem_0_5_129_rs_net_1, \mem_0_rs[2] , \mem_0_[2]_net_1 , 
        un1_mem_0_5_129_i, un1_mem_0_5_14_set_net_1, 
        un1_mem_0_5_138_rs_net_1, \mem_1_rs[2] , \mem_1_[2]_net_1 , 
        un1_mem_0_5_138_i, un1_mem_0_5_set_net_1, 
        un1_mem_0_5_161_rs_net_1, \mem_4_rs[0] , \mem_4_[0]_net_1 , 
        un1_mem_0_5_161_i, un1_mem_0_5_13_set_net_1, 
        un1_mem_0_5_172_rs_net_1, \mem_5_rs[0] , \mem_5_[0]_net_1 , 
        un1_mem_0_5_172_i, un1_mem_0_5_29_set_net_1, 
        un1_mem_0_5_188_rs_net_1, \mem_6_rs[0] , \mem_6_[0]_net_1 , 
        un1_mem_0_5_188_i, un1_mem_0_5_125_set_net_1, 
        un1_mem_0_5_204_rs_net_1, \mem_7_rs[0] , \mem_7_[0]_net_1 , 
        un1_mem_0_5_204_i, un1_mem_0_5_7_set_net_1, 
        un1_mem_0_5_219_rs_net_1, \mem_8_rs[0] , \mem_8_[0]_net_1 , 
        un1_mem_0_5_219_i, un1_mem_0_5_72_set_net_1, 
        un1_mem_0_5_175_rs_net_1, \mem_9_rs[0] , \mem_9_[0]_net_1 , 
        un1_mem_0_5_175_i, un1_mem_0_5_97_set_net_1, 
        un1_mem_0_5_191_rs_net_1, \mem_10_rs[0] , \mem_10_[0]_net_1 , 
        un1_mem_0_5_191_i, un1_mem_0_5_88_set_net_1, 
        un1_mem_0_5_207_rs_net_1, \mem_11_rs[0] , \mem_11_[0]_net_1 , 
        un1_mem_0_5_207_i, un1_mem_0_5_16_set_net_1, 
        un1_mem_0_5_222_rs_net_1, \mem_12_rs[0] , \mem_12_[0]_net_1 , 
        un1_mem_0_5_222_i, un1_mem_0_5_104_set_net_1, 
        un1_mem_0_5_232_rs_net_1, \mem_13_rs[0] , \mem_13_[0]_net_1 , 
        un1_mem_0_5_232_i, un1_mem_0_5_112_set_net_1, 
        un1_mem_0_5_240_rs_net_1, \mem_14_rs[0] , \mem_14_[0]_net_1 , 
        un1_mem_0_5_240_i, un1_mem_0_5_57_set_net_1, 
        un1_mem_0_5_248_rs_net_1, \mem_15_rs[0] , \mem_15_[0]_net_1 , 
        un1_mem_0_5_248_i, un1_mem_0_5_81_set_net_1, 
        un1_mem_0_5_128_rs_net_1, \mem_0_rs[1] , \mem_0_[1]_net_1 , 
        un1_mem_0_5_128_i, un1_mem_0_5_12_set_net_1, 
        un1_mem_0_5_137_rs_net_1, \mem_1_rs[1] , \mem_1_[1]_net_1 , 
        un1_mem_0_5_137_i, un1_mem_0_5_28_set_net_1, 
        un1_mem_0_5_145_rs_net_1, \mem_2_rs[1] , \mem_2_[1]_net_1 , 
        un1_mem_0_5_145_i, un1_mem_0_5_80_set_net_1, 
        un1_mem_0_5_131_rs_net_1, \mem_0_rs[0] , \mem_0_[0]_net_1 , 
        un1_mem_0_5_131_i, un1_mem_0_5_10_set_net_1, 
        un1_mem_0_5_136_rs_net_1, \mem_1_rs[0] , \mem_1_[0]_net_1 , 
        un1_mem_0_5_136_i, un1_mem_0_5_26_set_net_1, 
        un1_mem_0_5_144_rs_net_1, \mem_2_rs[0] , \mem_2_[0]_net_1 , 
        un1_mem_0_5_144_i, un1_mem_0_5_122_set_net_1, 
        un1_mem_0_5_152_rs_net_1, \mem_3_rs[0] , \mem_3_[0]_net_1 , 
        un1_mem_0_5_152_i, N_467, N_468, N_469, N_470, N_471, N_472, 
        N_473, N_474, N_475, N_476, N_477, N_478, N_479, N_480, N_481, 
        N_482, N_329, N_345, N_361, N_377, N_393, N_416, N_434, N_455, 
        \temp_data_2_15_i_7[3]_net_1 , \temp_data_2_15_i_5[3]_net_1 , 
        \temp_data_2_15_i_4[3]_net_1 , \temp_data_2_15_i_3[3]_net_1 , 
        \temp_data_2_15_i_2[3]_net_1 , \temp_data_2_15_i_1[3]_net_1 , 
        \temp_data_2_15_i_0[3]_net_1 , \temp_data_2_15_i_7[4]_net_1 , 
        \temp_data_2_15_i_5[4]_net_1 , \temp_data_2_15_i_4[4]_net_1 , 
        \temp_data_2_15_i_3[4]_net_1 , \temp_data_2_15_i_2[4]_net_1 , 
        \temp_data_2_15_i_1[4]_net_1 , \temp_data_2_15_i_0[4]_net_1 , 
        \temp_data_2_15_i_7[0]_net_1 , \temp_data_2_15_i_5[0]_net_1 , 
        \temp_data_2_15_i_4[0]_net_1 , \temp_data_2_15_i_3[0]_net_1 , 
        \temp_data_2_15_i_2[0]_net_1 , \temp_data_2_15_i_1[0]_net_1 , 
        \temp_data_2_15_i_0[0]_net_1 , \temp_data_2_15_i_7[5]_net_1 , 
        \temp_data_2_15_i_5[5]_net_1 , \temp_data_2_15_i_4[5]_net_1 , 
        \temp_data_2_15_i_3[5]_net_1 , \temp_data_2_15_i_2[5]_net_1 , 
        \temp_data_2_15_i_1[5]_net_1 , \temp_data_2_15_i_0[5]_net_1 , 
        \temp_data_2_15_i_7[1]_net_1 , \temp_data_2_15_i_5[1]_net_1 , 
        \temp_data_2_15_i_4[1]_net_1 , \temp_data_2_15_i_3[1]_net_1 , 
        \temp_data_2_15_i_2[1]_net_1 , \temp_data_2_15_i_1[1]_net_1 , 
        \temp_data_2_15_i_0[1]_net_1 , \temp_data_2_15_i_7[7]_net_1 , 
        \temp_data_2_15_i_5[7]_net_1 , \temp_data_2_15_i_4[7]_net_1 , 
        \temp_data_2_15_i_3[7]_net_1 , \temp_data_2_15_i_2[7]_net_1 , 
        \temp_data_2_15_i_1[7]_net_1 , \temp_data_2_15_i_0[7]_net_1 , 
        \temp_data_2_15_i_7[6]_net_1 , \temp_data_2_15_i_5[6]_net_1 , 
        \temp_data_2_15_i_4[6]_net_1 , \temp_data_2_15_i_3[6]_net_1 , 
        \temp_data_2_15_i_2[6]_net_1 , \temp_data_2_15_i_1[6]_net_1 , 
        \temp_data_2_15_i_0[6]_net_1 , \temp_data_2_15_i_7[2]_net_1 , 
        \temp_data_2_15_i_5[2]_net_1 , \temp_data_2_15_i_4[2]_net_1 , 
        \temp_data_2_15_i_3[2]_net_1 , \temp_data_2_15_i_2[2]_net_1 , 
        \temp_data_2_15_i_1[2]_net_1 , \temp_data_2_15_i_0[2]_net_1 , 
        \temp_data_2_15_i_11[3]_net_1 , \temp_data_2_15_i_11[4]_net_1 , 
        \temp_data_2_15_i_11[0]_net_1 , \temp_data_2_15_i_11[5]_net_1 , 
        \temp_data_2_15_i_11[1]_net_1 , \temp_data_2_15_i_11[7]_net_1 , 
        \temp_data_2_15_i_11[6]_net_1 , \temp_data_2_15_i_11[2]_net_1 , 
        \temp_data_2_15_i_12[3]_net_1 , \temp_data_2_15_i_12[4]_net_1 , 
        \temp_data_2_15_i_12[0]_net_1 , \temp_data_2_15_i_12[5]_net_1 , 
        \temp_data_2_15_i_12[1]_net_1 , \temp_data_2_15_i_12[7]_net_1 , 
        \temp_data_2_15_i_12[6]_net_1 , \temp_data_2_15_i_12[2]_net_1 ;
    
    CFG3 #( .INIT(8'hF2) )  un1_mem_0_5_145 (.A(\mem_2_[1]_net_1 ), .B(
        N_478), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_145_i));
    CFG4 #( .INIT(16'hFFFE) )  \temp_data_2_15_i_12[0]  (.A(
        \temp_data_2_15_i_3[0]_net_1 ), .B(
        \temp_data_2_15_i_2[0]_net_1 ), .C(
        \temp_data_2_15_i_1[0]_net_1 ), .D(
        \temp_data_2_15_i_0[0]_net_1 ), .Y(
        \temp_data_2_15_i_12[0]_net_1 ));
    SLE \mem_13_[4]  (.D(CoreAPB3_0_APBmslave2_PWDATA[4]), .CLK(
        FCCC_0_GL1), .EN(mem_13__1_sqmuxa), .ALn(un1_mem_0_5_236_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_13_rs[4] ));
    SLE un1_mem_0_5_215_rs (.D(VCC_net_1), .CLK(un1_mem_0_5_3_net_1), 
        .EN(VCC_net_1), .ALn(un1_mem_0_5_215_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(VCC_net_1), .Q(
        un1_mem_0_5_215_rs_net_1));
    SLE un1_mem_0_5_109_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_13__1_sqmuxa), .ALn(un1_mem_0_5_109_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_mem_0_5_109_set_net_1));
    SLE \mem_4_[5]  (.D(CoreAPB3_0_APBmslave2_PWDATA[5]), .CLK(
        FCCC_0_GL1), .EN(mem_4__1_sqmuxa), .ALn(un1_mem_0_5_166_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_4_rs[5] ));
    SLE \mem_12_[2]  (.D(CoreAPB3_0_APBmslave2_PWDATA[2]), .CLK(
        FCCC_0_GL1), .EN(mem_12__1_sqmuxa), .ALn(un1_mem_0_5_226_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_12_rs[2] ));
    SLE un1_mem_0_5_130_rs (.D(VCC_net_1), .CLK(un1_mem_0_5_84_net_1), 
        .EN(VCC_net_1), .ALn(un1_mem_0_5_130_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(VCC_net_1), .Q(
        un1_mem_0_5_130_rs_net_1));
    SLE un1_mem_0_5_193_rs (.D(VCC_net_1), .CLK(un1_mem_0_5_98_net_1), 
        .EN(VCC_net_1), .ALn(un1_mem_0_5_193_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(VCC_net_1), .Q(
        un1_mem_0_5_193_rs_net_1));
    CFG3 #( .INIT(8'hF2) )  un1_mem_0_5_251 (.A(\mem_15_[3]_net_1 ), 
        .B(N_474), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_251_i));
    CFG1 #( .INIT(2'h1) )  un1_mem_0_5_17_set_RNO (.A(
        un1_mem_0_5_17_net_1), .Y(un1_mem_0_5_17_i));
    CFG2 #( .INIT(4'h8) )  mem_15__1_sqmuxa_0_a2 (.A(N_474), .B(
        wr_enable), .Y(mem_15__1_sqmuxa));
    SLE un1_mem_0_5_107_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_13__1_sqmuxa), .ALn(un1_mem_0_5_107_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_mem_0_5_107_set_net_1));
    CFG3 #( .INIT(8'hF2) )  un1_mem_0_5_189 (.A(\mem_9_[7]_net_1 ), .B(
        N_467), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_189_i));
    CFG1 #( .INIT(2'h1) )  un1_mem_0_5_15_set_RNO (.A(
        un1_mem_0_5_15_net_1), .Y(un1_mem_0_5_15_i));
    SLE \mem_11_[4]  (.D(CoreAPB3_0_APBmslave2_PWDATA[4]), .CLK(
        FCCC_0_GL1), .EN(mem_11__1_sqmuxa), .ALn(un1_mem_0_5_214_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_11_rs[4] ));
    CFG3 #( .INIT(8'hF2) )  un1_mem_0_5_187 (.A(\mem_9_[6]_net_1 ), .B(
        N_467), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_187_i));
    CFG3 #( .INIT(8'hF8) )  un1_mem_0_5_198_rs_RNIA7I5 (.A(
        un1_mem_0_5_39_set_net_1), .B(un1_mem_0_5_198_rs_net_1), .C(
        \mem_6_rs[5] ), .Y(\mem_6_[5]_net_1 ));
    SLE \mem_13_[6]  (.D(CoreAPB3_0_APBmslave2_PWDATA[6]), .CLK(
        FCCC_0_GL1), .EN(mem_13__1_sqmuxa), .ALn(un1_mem_0_5_238_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_13_rs[6] ));
    CFG3 #( .INIT(8'h02) )  un1_mem_0_5_82 (.A(\mem_0_[2]_net_1 ), .B(
        N_473), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_82_net_1));
    CFG3 #( .INIT(8'hF2) )  un1_mem_0_5_199 (.A(\mem_10_[4]_net_1 ), 
        .B(N_471), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_199_i));
    SLE \mem_1_[2]  (.D(CoreAPB3_0_APBmslave2_PWDATA[2]), .CLK(
        FCCC_0_GL1), .EN(mem_1__1_sqmuxa), .ALn(un1_mem_0_5_138_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_1_rs[2] ));
    CFG3 #( .INIT(8'hF2) )  un1_mem_0_5_197 (.A(\mem_10_[3]_net_1 ), 
        .B(N_471), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_197_i));
    CFG4 #( .INIT(16'h7530) )  \temp_data_2_15_i_7[4]  (.A(
        \mem_12_[4]_net_1 ), .B(\mem_8_[4]_net_1 ), .C(N_479), .D(
        N_469), .Y(\temp_data_2_15_i_7[4]_net_1 ));
    SLE \mem_9_[2]  (.D(CoreAPB3_0_APBmslave2_PWDATA[2]), .CLK(
        FCCC_0_GL1), .EN(mem_9__1_sqmuxa), .ALn(un1_mem_0_5_179_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_9_rs[2] ));
    SLE \mem_6_[1]  (.D(CoreAPB3_0_APBmslave2_PWDATA[1]), .CLK(
        FCCC_0_GL1), .EN(mem_6__1_sqmuxa), .ALn(un1_mem_0_5_190_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_6_rs[1] ));
    SLE un1_mem_0_5_99_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_10__1_sqmuxa), .ALn(un1_mem_0_5_99_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_mem_0_5_99_set_net_1));
    CFG3 #( .INIT(8'hF2) )  un1_mem_0_5_135 (.A(\mem_0_[7]_net_1 ), .B(
        N_473), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_135_i));
    SLE un1_mem_0_5_203_rs (.D(VCC_net_1), .CLK(un1_mem_0_5_103_net_1), 
        .EN(VCC_net_1), .ALn(un1_mem_0_5_203_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(VCC_net_1), .Q(
        un1_mem_0_5_203_rs_net_1));
    CFG3 #( .INIT(8'hF8) )  \mem_15__RNIL8TK[1]  (.A(
        un1_mem_0_5_59_set_net_1), .B(un1_mem_0_5_249_rs_net_1), .C(
        \mem_15_rs[1] ), .Y(\mem_15_[1]_net_1 ));
    CFG3 #( .INIT(8'h02) )  un1_mem_0_5_41 (.A(\mem_1_[4]_net_1 ), .B(
        N_481), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_41_net_1));
    SLE un1_mem_0_5_29_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_6__1_sqmuxa), .ALn(un1_mem_0_5_29_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_mem_0_5_29_set_net_1));
    CFG3 #( .INIT(8'hF2) )  un1_mem_0_5_241 (.A(\mem_14_[1]_net_1 ), 
        .B(N_482), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_241_i));
    CFG3 #( .INIT(8'h02) )  un1_mem_0_5_65 (.A(\mem_4_[4]_net_1 ), .B(
        N_476), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_65_net_1));
    CFG3 #( .INIT(8'hF2) )  un1_mem_0_5_168 (.A(\mem_4_[6]_net_1 ), .B(
        N_476), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_168_i));
    CFG3 #( .INIT(8'hF2) )  un1_mem_0_5_174 (.A(\mem_5_[1]_net_1 ), .B(
        N_472), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_174_i));
    CFG1 #( .INIT(2'h1) )  un1_mem_0_5_80_set_RNO (.A(
        un1_mem_0_5_80_net_1), .Y(un1_mem_0_5_80_i));
    CFG4 #( .INIT(16'h7350) )  \temp_data_2_15_i_1[3]  (.A(
        \mem_11_[3]_net_1 ), .B(\mem_3_[3]_net_1 ), .C(N_475), .D(
        N_470), .Y(\temp_data_2_15_i_1[3]_net_1 ));
    SLE \mem_11_[6]  (.D(CoreAPB3_0_APBmslave2_PWDATA[6]), .CLK(
        FCCC_0_GL1), .EN(mem_11__1_sqmuxa), .ALn(un1_mem_0_5_218_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_11_rs[6] ));
    SLE \mem_0_[1]  (.D(CoreAPB3_0_APBmslave2_PWDATA[1]), .CLK(
        FCCC_0_GL1), .EN(mem_0__1_sqmuxa), .ALn(un1_mem_0_5_128_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_0_rs[1] ));
    SLE un1_mem_0_5_187_rs (.D(VCC_net_1), .CLK(un1_mem_0_5_78_net_1), 
        .EN(VCC_net_1), .ALn(un1_mem_0_5_187_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(VCC_net_1), .Q(
        un1_mem_0_5_187_rs_net_1));
    CFG3 #( .INIT(8'hF2) )  un1_mem_0_5_247 (.A(\mem_14_[7]_net_1 ), 
        .B(N_482), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_247_i));
    SLE un1_mem_0_5_168_rs (.D(VCC_net_1), .CLK(un1_mem_0_5_9_net_1), 
        .EN(VCC_net_1), .ALn(un1_mem_0_5_168_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(VCC_net_1), .Q(
        un1_mem_0_5_168_rs_net_1));
    CFG1 #( .INIT(2'h1) )  un1_mem_0_5_63_set_RNO (.A(
        un1_mem_0_5_63_net_1), .Y(un1_mem_0_5_63_i));
    CFG3 #( .INIT(8'hF8) )  \mem_11__RNICVCQ[7]  (.A(
        un1_mem_0_5_95_set_net_1), .B(un1_mem_0_5_220_rs_net_1), .C(
        \mem_11_rs[7] ), .Y(\mem_11_[7]_net_1 ));
    CFG3 #( .INIT(8'h02) )  un1_mem_0_5_64 (.A(\mem_8_[2]_net_1 ), .B(
        N_479), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_64_net_1));
    SLE un1_mem_0_5_220_rs (.D(VCC_net_1), .CLK(un1_mem_0_5_95_net_1), 
        .EN(VCC_net_1), .ALn(un1_mem_0_5_220_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(VCC_net_1), .Q(
        un1_mem_0_5_220_rs_net_1));
    CFG3 #( .INIT(8'hF2) )  un1_mem_0_5_153 (.A(\mem_3_[1]_net_1 ), .B(
        N_470), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_153_i));
    CFG3 #( .INIT(8'hF2) )  un1_mem_0_5_231 (.A(\mem_12_[7]_net_1 ), 
        .B(N_469), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_231_i));
    CFG4 #( .INIT(16'h0001) )  \temp_data_RNO[4]  (.A(
        \temp_data_2_15_i_4[4]_net_1 ), .B(
        \temp_data_2_15_i_5[4]_net_1 ), .C(
        \temp_data_2_15_i_11[4]_net_1 ), .D(
        \temp_data_2_15_i_12[4]_net_1 ), .Y(N_16_i_0));
    SLE un1_mem_0_5_48_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_3__1_sqmuxa), .ALn(un1_mem_0_5_48_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_mem_0_5_48_set_net_1));
    CFG3 #( .INIT(8'hF2) )  un1_mem_0_5_222 (.A(\mem_12_[0]_net_1 ), 
        .B(N_469), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_222_i));
    CFG1 #( .INIT(2'h1) )  un1_mem_0_5_19_set_RNO (.A(
        un1_mem_0_5_19_net_1), .Y(un1_mem_0_5_19_i));
    SLE un1_mem_0_5_51_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_7__1_sqmuxa), .ALn(un1_mem_0_5_51_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_mem_0_5_51_set_net_1));
    CFG3 #( .INIT(8'hF8) )  un1_mem_0_5_74_set_RNI8B5V (.A(
        un1_mem_0_5_74_set_net_1), .B(un1_mem_0_5_179_rs_net_1), .C(
        \mem_9_rs[2] ), .Y(\mem_9_[2]_net_1 ));
    CFG3 #( .INIT(8'h02) )  un1_mem_0_5_105 (.A(\mem_13_[1]_net_1 ), 
        .B(N_477), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_105_net_1));
    CFG3 #( .INIT(8'hF2) )  un1_mem_0_5_237 (.A(\mem_13_[5]_net_1 ), 
        .B(N_477), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_237_i));
    CFG1 #( .INIT(2'h1) )  un1_mem_0_5_8_set_RNO (.A(
        un1_mem_0_5_8_net_1), .Y(un1_mem_0_5_8_i));
    SLE un1_mem_0_5_178_rs (.D(VCC_net_1), .CLK(un1_mem_0_5_42_net_1), 
        .EN(VCC_net_1), .ALn(un1_mem_0_5_178_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(VCC_net_1), .Q(
        un1_mem_0_5_178_rs_net_1));
    CFG4 #( .INIT(16'h1000) )  \WRITE_GEN.mem_3__2_i_a2[1]  (.A(
        CoreAPB3_0_APBmslave2_PADDR[3]), .B(
        CoreAPB3_0_APBmslave2_PADDR[2]), .C(
        CoreAPB3_0_APBmslave2_PADDR[0]), .D(
        CoreAPB3_0_APBmslave2_PADDR[1]), .Y(N_470));
    CFG3 #( .INIT(8'hF8) )  un1_mem_0_5_175_rs_RNI0LC21 (.A(
        un1_mem_0_5_72_set_net_1), .B(un1_mem_0_5_175_rs_net_1), .C(
        \mem_9_rs[0] ), .Y(\mem_9_[0]_net_1 ));
    SLE un1_mem_0_5_250_rs (.D(VCC_net_1), .CLK(un1_mem_0_5_56_net_1), 
        .EN(VCC_net_1), .ALn(un1_mem_0_5_250_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(VCC_net_1), .Q(
        un1_mem_0_5_250_rs_net_1));
    CFG4 #( .INIT(16'h7350) )  \temp_data_2_15_i_4[5]  (.A(
        \mem_10_[5]_net_1 ), .B(\mem_6_[5]_net_1 ), .C(N_471), .D(
        N_468), .Y(\temp_data_2_15_i_4[5]_net_1 ));
    SLE \mem_8_[3]  (.D(CoreAPB3_0_APBmslave2_PWDATA[3]), .CLK(
        FCCC_0_GL1), .EN(mem_8__1_sqmuxa), .ALn(un1_mem_0_5_225_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_8_rs[3] ));
    CFG3 #( .INIT(8'hF2) )  un1_mem_0_5_143 (.A(\mem_1_[7]_net_1 ), .B(
        N_481), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_143_i));
    CFG3 #( .INIT(8'h02) )  un1_mem_0_5_63 (.A(\mem_15_[6]_net_1 ), .B(
        N_474), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_63_net_1));
    CFG3 #( .INIT(8'hF8) )  un1_mem_0_5_204_rs_RNI6O5C (.A(
        un1_mem_0_5_125_set_net_1), .B(un1_mem_0_5_204_rs_net_1), .C(
        \mem_7_rs[0] ), .Y(\mem_7_[0]_net_1 ));
    CFG3 #( .INIT(8'hF8) )  un1_mem_0_5_172_rs_RNIK1KK (.A(
        un1_mem_0_5_13_set_net_1), .B(un1_mem_0_5_172_rs_net_1), .C(
        \mem_5_rs[0] ), .Y(\mem_5_[0]_net_1 ));
    CFG1 #( .INIT(2'h1) )  un1_mem_0_5_117_set_RNO (.A(
        un1_mem_0_5_117_net_1), .Y(un1_mem_0_5_117_i));
    CFG3 #( .INIT(8'hF2) )  un1_mem_0_5_184 (.A(\mem_5_[6]_net_1 ), .B(
        N_472), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_184_i));
    CFG3 #( .INIT(8'hF2) )  un1_mem_0_5_159 (.A(\mem_3_[6]_net_1 ), .B(
        N_470), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_159_i));
    CFG3 #( .INIT(8'hF2) )  un1_mem_0_5_157 (.A(\mem_3_[5]_net_1 ), .B(
        N_470), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_157_i));
    CFG1 #( .INIT(2'h1) )  un1_mem_0_5_114_set_RNO (.A(
        un1_mem_0_5_114_net_1), .Y(un1_mem_0_5_114_i));
    CFG1 #( .INIT(2'h1) )  un1_mem_0_5_77_set_RNO (.A(
        un1_mem_0_5_77_net_1), .Y(un1_mem_0_5_77_i));
    CFG3 #( .INIT(8'hF8) )  un1_mem_0_5_35_set_RNI09DG (.A(
        un1_mem_0_5_35_set_net_1), .B(un1_mem_0_5_194_rs_net_1), .C(
        \mem_6_rs[3] ), .Y(\mem_6_[3]_net_1 ));
    CFG3 #( .INIT(8'hF8) )  un1_mem_0_5_243_rs_RNIP2DD (.A(
        un1_mem_0_5_115_set_net_1), .B(un1_mem_0_5_243_rs_net_1), .C(
        \mem_14_rs[3] ), .Y(\mem_14_[3]_net_1 ));
    SLE \mem_1_[1]  (.D(CoreAPB3_0_APBmslave2_PWDATA[1]), .CLK(
        FCCC_0_GL1), .EN(mem_1__1_sqmuxa), .ALn(un1_mem_0_5_137_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_1_rs[1] ));
    CFG3 #( .INIT(8'hF2) )  un1_mem_0_5_194 (.A(\mem_6_[3]_net_1 ), .B(
        N_468), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_194_i));
    SLE \mem_9_[1]  (.D(CoreAPB3_0_APBmslave2_PWDATA[1]), .CLK(
        FCCC_0_GL1), .EN(mem_9__1_sqmuxa), .ALn(un1_mem_0_5_177_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_9_rs[1] ));
    CFG3 #( .INIT(8'h02) )  un1_mem_0_5_12 (.A(\mem_1_[1]_net_1 ), .B(
        N_481), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_12_net_1));
    CFG4 #( .INIT(16'h0001) )  \temp_data_RNO[6]  (.A(
        \temp_data_2_15_i_4[6]_net_1 ), .B(
        \temp_data_2_15_i_5[6]_net_1 ), .C(
        \temp_data_2_15_i_11[6]_net_1 ), .D(
        \temp_data_2_15_i_12[6]_net_1 ), .Y(N_47_i_0));
    CFG1 #( .INIT(2'h1) )  un1_mem_0_5_125_set_RNO (.A(
        un1_mem_0_5_125_net_1), .Y(un1_mem_0_5_125_i));
    SLE \mem_12_[7]  (.D(CoreAPB3_0_APBmslave2_PWDATA[7]), .CLK(
        FCCC_0_GL1), .EN(mem_12__1_sqmuxa), .ALn(un1_mem_0_5_231_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_12_rs[7] ));
    CFG3 #( .INIT(8'hF8) )  \mem_3__RNIU02R[3]  (.A(
        un1_mem_0_5_48_set_net_1), .B(un1_mem_0_5_155_rs_net_1), .C(
        \mem_3_rs[3] ), .Y(\mem_3_[3]_net_1 ));
    CFG1 #( .INIT(2'h1) )  un1_mem_0_5_75_set_RNO (.A(
        un1_mem_0_5_75_net_1), .Y(un1_mem_0_5_75_i));
    CFG1 #( .INIT(2'h1) )  un1_mem_0_5_120_set_RNO (.A(
        un1_mem_0_5_120_net_1), .Y(un1_mem_0_5_120_i));
    CFG3 #( .INIT(8'h02) )  un1_mem_0_5_9 (.A(\mem_4_[6]_net_1 ), .B(
        N_476), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_9_net_1));
    CFG3 #( .INIT(8'h02) )  un1_mem_0_5_126 (.A(\mem_3_[2]_net_1 ), .B(
        N_470), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_126_net_1));
    SLE \mem_14_[0]  (.D(CoreAPB3_0_APBmslave2_PWDATA[0]), .CLK(
        FCCC_0_GL1), .EN(mem_14__1_sqmuxa), .ALn(un1_mem_0_5_240_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_14_rs[0] ));
    CFG3 #( .INIT(8'hF8) )  un1_mem_0_5_set_RNIEHIN (.A(
        un1_mem_0_5_set_net_1), .B(un1_mem_0_5_161_rs_net_1), .C(
        \mem_4_rs[0] ), .Y(\mem_4_[0]_net_1 ));
    SLE un1_mem_0_5_223_rs (.D(VCC_net_1), .CLK(un1_mem_0_5_64_net_1), 
        .EN(VCC_net_1), .ALn(un1_mem_0_5_223_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(VCC_net_1), .Q(
        un1_mem_0_5_223_rs_net_1));
    CFG3 #( .INIT(8'hF8) )  un1_mem_0_5_142_rs_RNIO2KU (.A(
        un1_mem_0_5_45_set_net_1), .B(un1_mem_0_5_142_rs_net_1), .C(
        \mem_1_rs[6] ), .Y(\mem_1_[6]_net_1 ));
    SLE \mem_10_[5]  (.D(CoreAPB3_0_APBmslave2_PWDATA[5]), .CLK(
        FCCC_0_GL1), .EN(mem_10__1_sqmuxa), .ALn(un1_mem_0_5_201_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_10_rs[5] ));
    CFG3 #( .INIT(8'hF2) )  un1_mem_0_5_201 (.A(\mem_10_[5]_net_1 ), 
        .B(N_471), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_201_i));
    CFG3 #( .INIT(8'hF2) )  un1_mem_0_5_133 (.A(\mem_0_[5]_net_1 ), .B(
        N_473), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_133_i));
    SLE un1_mem_0_5_249_rs (.D(VCC_net_1), .CLK(un1_mem_0_5_59_net_1), 
        .EN(VCC_net_1), .ALn(un1_mem_0_5_249_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(VCC_net_1), .Q(
        un1_mem_0_5_249_rs_net_1));
    CFG3 #( .INIT(8'hF2) )  un1_mem_0_5_149 (.A(\mem_2_[5]_net_1 ), .B(
        N_478), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_149_i));
    SLE un1_mem_0_5_114_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_14__1_sqmuxa), .ALn(un1_mem_0_5_114_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_mem_0_5_114_set_net_1));
    CFG3 #( .INIT(8'h02) )  un1_mem_0_5_47 (.A(\mem_1_[5]_net_1 ), .B(
        N_481), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_47_net_1));
    CFG3 #( .INIT(8'hF8) )  un1_mem_0_5_113_set_RNIJIQI (.A(
        un1_mem_0_5_113_set_net_1), .B(un1_mem_0_5_241_rs_net_1), .C(
        \mem_14_rs[1] ), .Y(\mem_14_[1]_net_1 ));
    CFG3 #( .INIT(8'hF2) )  un1_mem_0_5_147 (.A(\mem_2_[3]_net_1 ), .B(
        N_478), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_147_i));
    CFG4 #( .INIT(16'h7350) )  \temp_data_2_15_i_5[1]  (.A(
        \mem_7_[1]_net_1 ), .B(\mem_5_[1]_net_1 ), .C(N_480), .D(N_472)
        , .Y(\temp_data_2_15_i_5[1]_net_1 ));
    SLE \data_out[5]  (.D(\temp_data[5]_net_1 ), .CLK(FCCC_0_GL1), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(
        CoreAPB3_0_APBmslave3_PRDATA[5]));
    CFG1 #( .INIT(2'h1) )  un1_mem_0_5_10_set_RNO (.A(
        un1_mem_0_5_10_net_1), .Y(un1_mem_0_5_10_i));
    SLE \mem_5_[2]  (.D(CoreAPB3_0_APBmslave2_PWDATA[2]), .CLK(
        FCCC_0_GL1), .EN(mem_5__1_sqmuxa), .ALn(un1_mem_0_5_176_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_5_rs[2] ));
    CFG1 #( .INIT(2'h1) )  un1_mem_0_5_107_set_RNO (.A(
        un1_mem_0_5_107_net_1), .Y(un1_mem_0_5_107_i));
    CFG3 #( .INIT(8'hF2) )  un1_mem_0_5_207 (.A(\mem_11_[0]_net_1 ), 
        .B(N_475), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_207_i));
    SLE un1_mem_0_5_106_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_13__1_sqmuxa), .ALn(un1_mem_0_5_106_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_mem_0_5_106_set_net_1));
    SLE un1_mem_0_5_10_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_1__1_sqmuxa), .ALn(un1_mem_0_5_10_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_mem_0_5_10_set_net_1));
    SLE \mem_6_[6]  (.D(CoreAPB3_0_APBmslave2_PWDATA[6]), .CLK(
        FCCC_0_GL1), .EN(mem_6__1_sqmuxa), .ALn(un1_mem_0_5_200_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_6_rs[6] ));
    CFG1 #( .INIT(2'h1) )  un1_mem_0_5_64_set_RNO (.A(
        un1_mem_0_5_64_net_1), .Y(un1_mem_0_5_64_i));
    CFG1 #( .INIT(2'h1) )  un1_mem_0_5_104_set_RNO (.A(
        un1_mem_0_5_104_net_1), .Y(un1_mem_0_5_104_i));
    CFG3 #( .INIT(8'hF8) )  \mem_3__RNISIGN[7]  (.A(
        un1_mem_0_5_55_set_net_1), .B(un1_mem_0_5_160_rs_net_1), .C(
        \mem_3_rs[7] ), .Y(\mem_3_[7]_net_1 ));
    SLE un1_mem_0_5_61_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_15__1_sqmuxa), .ALn(un1_mem_0_5_61_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_mem_0_5_61_set_net_1));
    SLE un1_mem_0_5_253_rs (.D(VCC_net_1), .CLK(un1_mem_0_5_58_net_1), 
        .EN(VCC_net_1), .ALn(un1_mem_0_5_253_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(VCC_net_1), .Q(
        un1_mem_0_5_253_rs_net_1));
    SLE \mem_10_[1]  (.D(CoreAPB3_0_APBmslave2_PWDATA[1]), .CLK(
        FCCC_0_GL1), .EN(mem_10__1_sqmuxa), .ALn(un1_mem_0_5_193_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_10_rs[1] ));
    CFG1 #( .INIT(2'h1) )  un1_mem_0_5_96_set_RNO (.A(
        un1_mem_0_5_96_net_1), .Y(un1_mem_0_5_96_i));
    CFG3 #( .INIT(8'hF8) )  un1_mem_0_5_183_rs_RNI77551 (.A(
        un1_mem_0_5_76_set_net_1), .B(un1_mem_0_5_183_rs_net_1), .C(
        \mem_9_rs[4] ), .Y(\mem_9_[4]_net_1 ));
    CFG4 #( .INIT(16'h7530) )  \temp_data_2_15_i_7[6]  (.A(
        \mem_12_[6]_net_1 ), .B(\mem_8_[6]_net_1 ), .C(N_479), .D(
        N_469), .Y(\temp_data_2_15_i_7[6]_net_1 ));
    CFG3 #( .INIT(8'hF8) )  \mem_2__RNI4TJP[7]  (.A(
        un1_mem_0_5_120_set_net_1), .B(un1_mem_0_5_151_rs_net_1), .C(
        \mem_2_rs[7] ), .Y(\mem_2_[7]_net_1 ));
    CFG3 #( .INIT(8'hF8) )  un1_mem_0_5_43_set_RNIP8NP (.A(
        un1_mem_0_5_43_set_net_1), .B(un1_mem_0_5_139_rs_net_1), .C(
        \mem_1_rs[3] ), .Y(\mem_1_[3]_net_1 ));
    CFG4 #( .INIT(16'h0008) )  \WRITE_GEN.mem_12__2_i_a2[4]  (.A(
        CoreAPB3_0_APBmslave2_PADDR[3]), .B(
        CoreAPB3_0_APBmslave2_PADDR[2]), .C(
        CoreAPB3_0_APBmslave2_PADDR[0]), .D(
        CoreAPB3_0_APBmslave2_PADDR[1]), .Y(N_469));
    CFG3 #( .INIT(8'h02) )  un1_mem_0_5_60 (.A(\mem_15_[7]_net_1 ), .B(
        N_474), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_60_net_1));
    CFG3 #( .INIT(8'h02) )  un1_mem_0_5_3 (.A(\mem_7_[6]_net_1 ), .B(
        N_480), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_3_net_1));
    CFG4 #( .INIT(16'h7530) )  \temp_data_2_15_i_0[3]  (.A(
        \mem_9_[3]_net_1 ), .B(\mem_1_[3]_net_1 ), .C(N_481), .D(N_467)
        , .Y(\temp_data_2_15_i_0[3]_net_1 ));
    CFG1 #( .INIT(2'h1) )  un1_mem_0_5_98_set_RNO (.A(
        un1_mem_0_5_98_net_1), .Y(un1_mem_0_5_98_i));
    SLE un1_mem_0_5_208_rs (.D(VCC_net_1), .CLK(un1_mem_0_5_49_net_1), 
        .EN(VCC_net_1), .ALn(un1_mem_0_5_208_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(VCC_net_1), .Q(
        un1_mem_0_5_208_rs_net_1));
    SLE un1_mem_0_5_70_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_8__1_sqmuxa), .ALn(un1_mem_0_5_70_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_mem_0_5_70_set_net_1));
    CFG3 #( .INIT(8'hF2) )  un1_mem_0_5_139 (.A(\mem_1_[3]_net_1 ), .B(
        N_481), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_139_i));
    CFG3 #( .INIT(8'hF2) )  un1_mem_0_5_137 (.A(\mem_1_[1]_net_1 ), .B(
        N_481), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_137_i));
    SLE un1_mem_0_5_146_rs (.D(VCC_net_1), .CLK(un1_mem_0_5_30_net_1), 
        .EN(VCC_net_1), .ALn(un1_mem_0_5_146_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(VCC_net_1), .Q(
        un1_mem_0_5_146_rs_net_1));
    SLE \mem_0_[6]  (.D(CoreAPB3_0_APBmslave2_PWDATA[6]), .CLK(
        FCCC_0_GL1), .EN(mem_0__1_sqmuxa), .ALn(un1_mem_0_5_134_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_0_rs[6] ));
    SLE un1_mem_0_5_207_rs (.D(VCC_net_1), .CLK(un1_mem_0_5_88_net_1), 
        .EN(VCC_net_1), .ALn(un1_mem_0_5_207_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(VCC_net_1), .Q(
        un1_mem_0_5_207_rs_net_1));
    SLE \temp_data[5]  (.D(N_39_i_0), .CLK(FCCC_0_GL1), .EN(rd_enable), 
        .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\temp_data[5]_net_1 ));
    SLE un1_mem_0_5_157_rs (.D(VCC_net_1), .CLK(un1_mem_0_5_52_net_1), 
        .EN(VCC_net_1), .ALn(un1_mem_0_5_157_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(VCC_net_1), .Q(
        un1_mem_0_5_157_rs_net_1));
    CFG1 #( .INIT(2'h1) )  un1_mem_0_5_79_set_RNO (.A(
        un1_mem_0_5_79_net_1), .Y(un1_mem_0_5_79_i));
    CFG3 #( .INIT(8'hF8) )  un1_mem_0_5_132_rs_RNIOCGF (.A(
        un1_mem_0_5_85_set_net_1), .B(un1_mem_0_5_132_rs_net_1), .C(
        \mem_0_rs[4] ), .Y(\mem_0_[4]_net_1 ));
    CFG3 #( .INIT(8'h02) )  un1_mem_0_5_21 (.A(\mem_12_[5]_net_1 ), .B(
        N_469), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_21_net_1));
    CFG3 #( .INIT(8'hF2) )  un1_mem_0_5_246 (.A(\mem_14_[6]_net_1 ), 
        .B(N_482), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_246_i));
    SLE un1_mem_0_5_43_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_1__1_sqmuxa), .ALn(un1_mem_0_5_43_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_mem_0_5_43_set_net_1));
    SLE un1_mem_0_5_112_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_14__1_sqmuxa), .ALn(un1_mem_0_5_112_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_mem_0_5_112_set_net_1));
    CFG3 #( .INIT(8'h02) )  un1_mem_0_5_103 (.A(\mem_10_[6]_net_1 ), 
        .B(N_471), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_103_net_1));
    CFG3 #( .INIT(8'h02) )  un1_mem_0_5_48 (.A(\mem_3_[3]_net_1 ), .B(
        N_470), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_48_net_1));
    CFG3 #( .INIT(8'hF2) )  un1_mem_0_5_154 (.A(\mem_3_[2]_net_1 ), .B(
        N_470), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_154_i));
    CFG4 #( .INIT(16'h7530) )  \temp_data_2_15_i_7[3]  (.A(
        \mem_12_[3]_net_1 ), .B(\mem_8_[3]_net_1 ), .C(N_479), .D(
        N_469), .Y(\temp_data_2_15_i_7[3]_net_1 ));
    SLE un1_mem_0_5_54_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_7__1_sqmuxa), .ALn(un1_mem_0_5_54_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_mem_0_5_54_set_net_1));
    SLE un1_mem_0_5_80_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_0__1_sqmuxa), .ALn(un1_mem_0_5_80_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_mem_0_5_80_set_net_1));
    CFG3 #( .INIT(8'h02) )  un1_mem_0_5_49 (.A(\mem_7_[2]_net_1 ), .B(
        N_480), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_49_net_1));
    CFG4 #( .INIT(16'h7350) )  \temp_data_2_15_i_2[6]  (.A(
        \mem_13_[6]_net_1 ), .B(\mem_15_[6]_net_1 ), .C(N_477), .D(
        N_474), .Y(\temp_data_2_15_i_2[6]_net_1 ));
    CFG3 #( .INIT(8'h02) )  un1_mem_0_5_86 (.A(\mem_0_[5]_net_1 ), .B(
        N_473), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_86_net_1));
    CFG1 #( .INIT(2'h1) )  un1_mem_0_5_1_set_RNO (.A(
        un1_mem_0_5_1_net_1), .Y(un1_mem_0_5_1_i));
    CFG4 #( .INIT(16'h7350) )  \temp_data_2_15_i_3[4]  (.A(
        \mem_14_[4]_net_1 ), .B(\mem_2_[4]_net_1 ), .C(N_482), .D(
        N_478), .Y(\temp_data_2_15_i_3[4]_net_1 ));
    CFG3 #( .INIT(8'hF2) )  un1_mem_0_5_220 (.A(\mem_11_[7]_net_1 ), 
        .B(N_475), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_220_i));
    CFG3 #( .INIT(8'h02) )  un1_mem_0_5_72 (.A(\mem_9_[0]_net_1 ), .B(
        N_467), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_72_net_1));
    CFG3 #( .INIT(8'h02) )  un1_mem_0_5_51 (.A(\mem_7_[3]_net_1 ), .B(
        N_480), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_51_net_1));
    CFG1 #( .INIT(2'h1) )  un1_mem_0_5_86_set_RNO (.A(
        un1_mem_0_5_86_net_1), .Y(un1_mem_0_5_86_i));
    CFG1 #( .INIT(2'h1) )  un1_mem_0_5_92_set_RNO (.A(
        un1_mem_0_5_92_net_1), .Y(un1_mem_0_5_92_i));
    SLE un1_mem_0_5_124_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_3__1_sqmuxa), .ALn(un1_mem_0_5_124_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_mem_0_5_124_set_net_1));
    CFG3 #( .INIT(8'hF2) )  un1_mem_0_5_236 (.A(\mem_13_[4]_net_1 ), 
        .B(N_477), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_236_i));
    CFG3 #( .INIT(8'hF2) )  un1_mem_0_5_144 (.A(\mem_2_[0]_net_1 ), .B(
        N_478), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_144_i));
    SLE un1_mem_0_5_239_rs (.D(VCC_net_1), .CLK(un1_mem_0_5_111_net_1), 
        .EN(VCC_net_1), .ALn(un1_mem_0_5_239_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(VCC_net_1), .Q(
        un1_mem_0_5_239_rs_net_1));
    CFG1 #( .INIT(2'h1) )  un1_mem_0_5_88_set_RNO (.A(
        un1_mem_0_5_88_net_1), .Y(un1_mem_0_5_88_i));
    CFG4 #( .INIT(16'h7350) )  \temp_data_2_15_i_4[2]  (.A(
        \mem_10_[2]_net_1 ), .B(\mem_6_[2]_net_1 ), .C(N_471), .D(
        N_468), .Y(\temp_data_2_15_i_4[2]_net_1 ));
    SLE \mem_5_[1]  (.D(CoreAPB3_0_APBmslave2_PWDATA[1]), .CLK(
        FCCC_0_GL1), .EN(mem_5__1_sqmuxa), .ALn(un1_mem_0_5_174_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_5_rs[1] ));
    SLE un1_mem_0_5_214_rs (.D(VCC_net_1), .CLK(un1_mem_0_5_92_net_1), 
        .EN(VCC_net_1), .ALn(un1_mem_0_5_214_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(VCC_net_1), .Q(
        un1_mem_0_5_214_rs_net_1));
    SLE un1_mem_0_5_47_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_1__1_sqmuxa), .ALn(un1_mem_0_5_47_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_mem_0_5_47_set_net_1));
    CFG3 #( .INIT(8'h02) )  un1_mem_0_5_109 (.A(\mem_13_[5]_net_1 ), 
        .B(N_477), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_109_net_1));
    GND GND (.Y(GND_net_1));
    CFG3 #( .INIT(8'h02) )  un1_mem_0_5_107 (.A(\mem_13_[3]_net_1 ), 
        .B(N_477), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_107_net_1));
    CFG2 #( .INIT(4'h8) )  mem_4__1_sqmuxa_0_a2 (.A(N_476), .B(
        wr_enable), .Y(mem_4__1_sqmuxa));
    SLE \mem_15_[2]  (.D(CoreAPB3_0_APBmslave2_PWDATA[2]), .CLK(
        FCCC_0_GL1), .EN(mem_15__1_sqmuxa), .ALn(un1_mem_0_5_250_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_15_rs[2] ));
    SLE \mem_1_[6]  (.D(CoreAPB3_0_APBmslave2_PWDATA[6]), .CLK(
        FCCC_0_GL1), .EN(mem_1__1_sqmuxa), .ALn(un1_mem_0_5_142_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_1_rs[6] ));
    SLE \mem_9_[6]  (.D(CoreAPB3_0_APBmslave2_PWDATA[6]), .CLK(
        FCCC_0_GL1), .EN(mem_9__1_sqmuxa), .ALn(un1_mem_0_5_187_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_9_rs[6] ));
    CFG3 #( .INIT(8'hF8) )  \mem_14__RNI2R8D[6]  (.A(
        un1_mem_0_5_118_set_net_1), .B(un1_mem_0_5_246_rs_net_1), .C(
        \mem_14_rs[6] ), .Y(\mem_14_[6]_net_1 ));
    SLE \mem_8_[4]  (.D(CoreAPB3_0_APBmslave2_PWDATA[4]), .CLK(
        FCCC_0_GL1), .EN(mem_8__1_sqmuxa), .ALn(un1_mem_0_5_167_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_8_rs[4] ));
    CFG2 #( .INIT(4'h8) )  mem_7__1_sqmuxa_0_a2 (.A(N_480), .B(
        wr_enable), .Y(mem_7__1_sqmuxa));
    CFG1 #( .INIT(2'h1) )  un1_mem_0_5_70_set_RNO (.A(
        un1_mem_0_5_70_net_1), .Y(un1_mem_0_5_70_i));
    CFG4 #( .INIT(16'hEFEE) )  \temp_data_2_15_i_11[3]  (.A(N_377), .B(
        \temp_data_2_15_i_7[3]_net_1 ), .C(\mem_0_[3]_net_1 ), .D(
        N_473), .Y(\temp_data_2_15_i_11[3]_net_1 ));
    SLE \mem_13_[3]  (.D(CoreAPB3_0_APBmslave2_PWDATA[3]), .CLK(
        FCCC_0_GL1), .EN(mem_13__1_sqmuxa), .ALn(un1_mem_0_5_235_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_13_rs[3] ));
    CFG4 #( .INIT(16'h7530) )  \temp_data_2_15_i_0[7]  (.A(
        \mem_9_[7]_net_1 ), .B(\mem_1_[7]_net_1 ), .C(N_481), .D(N_467)
        , .Y(\temp_data_2_15_i_0[7]_net_1 ));
    CFG3 #( .INIT(8'h02) )  un1_mem_0_5_121 (.A(\mem_6_[6]_net_1 ), .B(
        N_468), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_121_net_1));
    SLE un1_mem_0_5_12_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_1__1_sqmuxa), .ALn(un1_mem_0_5_12_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_mem_0_5_12_set_net_1));
    SLE un1_mem_0_5_46_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_5__1_sqmuxa), .ALn(un1_mem_0_5_46_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_mem_0_5_46_set_net_1));
    CFG3 #( .INIT(8'hF8) )  un1_mem_0_5_203_rs_RNIHO59 (.A(
        un1_mem_0_5_103_set_net_1), .B(un1_mem_0_5_203_rs_net_1), .C(
        \mem_10_rs[6] ), .Y(\mem_10_[6]_net_1 ));
    CFG3 #( .INIT(8'hF2) )  un1_mem_0_5_134 (.A(\mem_0_[6]_net_1 ), .B(
        N_473), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_134_i));
    CFG3 #( .INIT(8'hF8) )  \mem_15__RNIIISL[6]  (.A(
        un1_mem_0_5_63_set_net_1), .B(un1_mem_0_5_255_rs_net_1), .C(
        \mem_15_rs[6] ), .Y(\mem_15_[6]_net_1 ));
    SLE un1_mem_0_5_197_rs (.D(VCC_net_1), .CLK(un1_mem_0_5_96_net_1), 
        .EN(VCC_net_1), .ALn(un1_mem_0_5_197_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(VCC_net_1), .Q(
        un1_mem_0_5_197_rs_net_1));
    SLE un1_mem_0_5_228_rs (.D(VCC_net_1), .CLK(un1_mem_0_5_20_net_1), 
        .EN(VCC_net_1), .ALn(un1_mem_0_5_228_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(VCC_net_1), .Q(
        un1_mem_0_5_228_rs_net_1));
    CFG3 #( .INIT(8'hF8) )  un1_mem_0_5_66_set_RNI1G0Q (.A(
        un1_mem_0_5_66_set_net_1), .B(un1_mem_0_5_225_rs_net_1), .C(
        \mem_8_rs[3] ), .Y(\mem_8_[3]_net_1 ));
    SLE un1_mem_0_5_136_rs (.D(VCC_net_1), .CLK(un1_mem_0_5_10_net_1), 
        .EN(VCC_net_1), .ALn(un1_mem_0_5_136_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(VCC_net_1), .Q(
        un1_mem_0_5_136_rs_net_1));
    SLE \temp_data[7]  (.D(N_64_i_0), .CLK(FCCC_0_GL1), .EN(rd_enable), 
        .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\temp_data[7]_net_1 ));
    SLE un1_mem_0_5_185_rs (.D(VCC_net_1), .CLK(un1_mem_0_5_77_net_1), 
        .EN(VCC_net_1), .ALn(un1_mem_0_5_185_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(VCC_net_1), .Q(
        un1_mem_0_5_185_rs_net_1));
    SLE \mem_11_[3]  (.D(CoreAPB3_0_APBmslave2_PWDATA[3]), .CLK(
        FCCC_0_GL1), .EN(mem_11__1_sqmuxa), .ALn(un1_mem_0_5_212_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_11_rs[3] ));
    SLE un1_mem_0_5_227_rs (.D(VCC_net_1), .CLK(un1_mem_0_5_19_net_1), 
        .EN(VCC_net_1), .ALn(un1_mem_0_5_227_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(VCC_net_1), .Q(
        un1_mem_0_5_227_rs_net_1));
    SLE un1_mem_0_5_72_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_9__1_sqmuxa), .ALn(un1_mem_0_5_72_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_mem_0_5_72_set_net_1));
    SLE un1_mem_0_5_64_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_8__1_sqmuxa), .ALn(un1_mem_0_5_64_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_mem_0_5_64_set_net_1));
    CFG3 #( .INIT(8'hF2) )  un1_mem_0_5_214 (.A(\mem_11_[4]_net_1 ), 
        .B(N_475), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_214_i));
    CFG4 #( .INIT(16'hEFEE) )  \temp_data_2_15_i_11[7]  (.A(N_455), .B(
        \temp_data_2_15_i_7[7]_net_1 ), .C(\mem_0_[7]_net_1 ), .D(
        N_473), .Y(\temp_data_2_15_i_11[7]_net_1 ));
    SLE un1_mem_0_5_15_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_5__1_sqmuxa), .ALn(un1_mem_0_5_15_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_mem_0_5_15_set_net_1));
    SLE \mem_7_[3]  (.D(CoreAPB3_0_APBmslave2_PWDATA[3]), .CLK(
        FCCC_0_GL1), .EN(mem_7__1_sqmuxa), .ALn(un1_mem_0_5_210_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_7_rs[3] ));
    CFG3 #( .INIT(8'hF8) )  un1_mem_0_5_117_set_RNIVIV7 (.A(
        un1_mem_0_5_117_set_net_1), .B(un1_mem_0_5_245_rs_net_1), .C(
        \mem_14_rs[5] ), .Y(\mem_14_[5]_net_1 ));
    SLE un1_mem_0_5_122_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_3__1_sqmuxa), .ALn(un1_mem_0_5_122_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_mem_0_5_122_set_net_1));
    CFG1 #( .INIT(2'h1) )  un1_mem_0_5_37_set_RNO (.A(
        un1_mem_0_5_37_net_1), .Y(un1_mem_0_5_37_i));
    CFG3 #( .INIT(8'h02) )  un1_mem_0_5_118 (.A(\mem_14_[6]_net_1 ), 
        .B(N_482), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_118_net_1));
    SLE un1_mem_0_5_181_rs (.D(VCC_net_1), .CLK(un1_mem_0_5_75_net_1), 
        .EN(VCC_net_1), .ALn(un1_mem_0_5_181_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(VCC_net_1), .Q(
        un1_mem_0_5_181_rs_net_1));
    CFG4 #( .INIT(16'h7350) )  \temp_data_2_15_i_2[3]  (.A(
        \mem_13_[3]_net_1 ), .B(\mem_15_[3]_net_1 ), .C(N_477), .D(
        N_474), .Y(\temp_data_2_15_i_2[3]_net_1 ));
    CFG1 #( .INIT(2'h1) )  un1_mem_0_5_82_set_RNO (.A(
        un1_mem_0_5_82_net_1), .Y(un1_mem_0_5_82_i));
    CFG3 #( .INIT(8'hF2) )  un1_mem_0_5_206 (.A(\mem_7_[1]_net_1 ), .B(
        N_480), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_206_i));
    SLE \mem_2_[3]  (.D(CoreAPB3_0_APBmslave2_PWDATA[3]), .CLK(
        FCCC_0_GL1), .EN(mem_2__1_sqmuxa), .ALn(un1_mem_0_5_147_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_2_rs[3] ));
    CFG1 #( .INIT(2'h1) )  un1_mem_0_5_51_set_RNO (.A(
        un1_mem_0_5_51_net_1), .Y(un1_mem_0_5_51_i));
    SLE \temp_data[6]  (.D(N_47_i_0), .CLK(FCCC_0_GL1), .EN(rd_enable), 
        .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\temp_data[6]_net_1 ));
    CFG1 #( .INIT(2'h1) )  un1_mem_0_5_35_set_RNO (.A(
        un1_mem_0_5_35_net_1), .Y(un1_mem_0_5_35_i));
    CFG3 #( .INIT(8'h02) )  un1_mem_0_5_45 (.A(\mem_1_[6]_net_1 ), .B(
        N_481), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_45_net_1));
    CFG3 #( .INIT(8'h02) )  un1_mem_0_5_27 (.A(\mem_5_[7]_net_1 ), .B(
        N_472), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_27_net_1));
    SLE un1_mem_0_5_75_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_9__1_sqmuxa), .ALn(un1_mem_0_5_75_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_mem_0_5_75_set_net_1));
    CFG4 #( .INIT(16'hEFEE) )  \temp_data_2_15_i_11[0]  (.A(N_329), .B(
        \temp_data_2_15_i_7[0]_net_1 ), .C(\mem_0_[0]_net_1 ), .D(
        N_473), .Y(\temp_data_2_15_i_11[0]_net_1 ));
    CFG3 #( .INIT(8'h02) )  un1_mem_0_5_16 (.A(\mem_12_[0]_net_1 ), .B(
        N_469), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_16_net_1));
    SLE \mem_8_[0]  (.D(CoreAPB3_0_APBmslave2_PWDATA[0]), .CLK(
        FCCC_0_GL1), .EN(mem_8__1_sqmuxa), .ALn(un1_mem_0_5_219_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_8_rs[0] ));
    SLE \mem_4_[3]  (.D(CoreAPB3_0_APBmslave2_PWDATA[3]), .CLK(
        FCCC_0_GL1), .EN(mem_4__1_sqmuxa), .ALn(un1_mem_0_5_164_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_4_rs[3] ));
    CFG4 #( .INIT(16'h4000) )  \WRITE_GEN.mem_7__2_i_a2[6]  (.A(
        CoreAPB3_0_APBmslave2_PADDR[3]), .B(
        CoreAPB3_0_APBmslave2_PADDR[2]), .C(
        CoreAPB3_0_APBmslave2_PADDR[0]), .D(
        CoreAPB3_0_APBmslave2_PADDR[1]), .Y(N_480));
    CFG1 #( .INIT(2'h1) )  un1_mem_0_5_47_set_RNO (.A(
        un1_mem_0_5_47_net_1), .Y(un1_mem_0_5_47_i));
    CFG3 #( .INIT(8'hF8) )  un1_mem_0_5_140_rs_RNIGALR (.A(
        un1_mem_0_5_41_set_net_1), .B(un1_mem_0_5_140_rs_net_1), .C(
        \mem_1_rs[4] ), .Y(\mem_1_[4]_net_1 ));
    CFG1 #( .INIT(2'h1) )  un1_mem_0_5_112_set_RNO (.A(
        un1_mem_0_5_112_net_1), .Y(un1_mem_0_5_112_i));
    CFG3 #( .INIT(8'hF8) )  un1_mem_0_5_40_set_RNIQICR (.A(
        un1_mem_0_5_40_set_net_1), .B(un1_mem_0_5_176_rs_net_1), .C(
        \mem_5_rs[2] ), .Y(\mem_5_[2]_net_1 ));
    CFG3 #( .INIT(8'hF2) )  un1_mem_0_5_166 (.A(\mem_4_[5]_net_1 ), .B(
        N_476), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_166_i));
    SLE un1_mem_0_5_111_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_13__1_sqmuxa), .ALn(un1_mem_0_5_111_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_mem_0_5_111_set_net_1));
    SLE un1_mem_0_5_82_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_0__1_sqmuxa), .ALn(un1_mem_0_5_82_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_mem_0_5_82_set_net_1));
    SLE un1_mem_0_5_160_rs (.D(VCC_net_1), .CLK(un1_mem_0_5_55_net_1), 
        .EN(VCC_net_1), .ALn(un1_mem_0_5_160_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(VCC_net_1), .Q(
        un1_mem_0_5_160_rs_net_1));
    SLE un1_mem_0_5_91_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_11__1_sqmuxa), .ALn(un1_mem_0_5_91_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_mem_0_5_91_set_net_1));
    CFG1 #( .INIT(2'h1) )  un1_mem_0_5_45_set_RNO (.A(
        un1_mem_0_5_45_net_1), .Y(un1_mem_0_5_45_i));
    CFG4 #( .INIT(16'h7350) )  \temp_data_2_15_i_1[5]  (.A(
        \mem_11_[5]_net_1 ), .B(\mem_3_[5]_net_1 ), .C(N_475), .D(
        N_470), .Y(\temp_data_2_15_i_1[5]_net_1 ));
    CFG1 #( .INIT(2'h1) )  un1_mem_0_5_16_set_RNO (.A(
        un1_mem_0_5_16_net_1), .Y(un1_mem_0_5_16_i));
    SLE un1_mem_0_5_21_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_12__1_sqmuxa), .ALn(un1_mem_0_5_21_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_mem_0_5_21_set_net_1));
    CFG3 #( .INIT(8'h02) )  un1_mem_0_5_44 (.A(\mem_5_[4]_net_1 ), .B(
        N_472), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_44_net_1));
    CFG4 #( .INIT(16'h0001) )  \WRITE_GEN.mem_0__2_i_a2[6]  (.A(
        CoreAPB3_0_APBmslave2_PADDR[3]), .B(
        CoreAPB3_0_APBmslave2_PADDR[2]), .C(
        CoreAPB3_0_APBmslave2_PADDR[0]), .D(
        CoreAPB3_0_APBmslave2_PADDR[1]), .Y(N_473));
    CFG4 #( .INIT(16'h0001) )  \temp_data_RNO[1]  (.A(
        \temp_data_2_15_i_4[1]_net_1 ), .B(
        \temp_data_2_15_i_5[1]_net_1 ), .C(
        \temp_data_2_15_i_11[1]_net_1 ), .D(
        \temp_data_2_15_i_12[1]_net_1 ), .Y(N_8_i_0));
    CFG3 #( .INIT(8'h02) )  un1_mem_0_5_57 (.A(\mem_15_[0]_net_1 ), .B(
        N_474), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_57_net_1));
    CFG3 #( .INIT(8'h02) )  un1_mem_0_5_104 (.A(\mem_13_[0]_net_1 ), 
        .B(N_477), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_104_net_1));
    CFG1 #( .INIT(2'h1) )  un1_mem_0_5_18_set_RNO (.A(
        un1_mem_0_5_18_net_1), .Y(un1_mem_0_5_18_i));
    CFG4 #( .INIT(16'h7350) )  \temp_data_2_15_i_5[5]  (.A(
        \mem_7_[5]_net_1 ), .B(\mem_5_[5]_net_1 ), .C(N_480), .D(N_472)
        , .Y(\temp_data_2_15_i_5[5]_net_1 ));
    SLE un1_mem_0_5_85_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_0__1_sqmuxa), .ALn(un1_mem_0_5_85_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_mem_0_5_85_set_net_1));
    SLE un1_mem_0_5_216_rs (.D(VCC_net_1), .CLK(un1_mem_0_5_93_net_1), 
        .EN(VCC_net_1), .ALn(un1_mem_0_5_216_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(VCC_net_1), .Q(
        un1_mem_0_5_216_rs_net_1));
    SLE un1_mem_0_5_110_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_13__1_sqmuxa), .ALn(un1_mem_0_5_110_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_mem_0_5_110_set_net_1));
    CFG1 #( .INIT(2'h1) )  un1_mem_0_5_2_set_RNO (.A(
        un1_mem_0_5_2_net_1), .Y(un1_mem_0_5_2_i));
    SLE un1_mem_0_5_182_rs (.D(VCC_net_1), .CLK(un1_mem_0_5_46_net_1), 
        .EN(VCC_net_1), .ALn(un1_mem_0_5_182_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(VCC_net_1), .Q(
        un1_mem_0_5_182_rs_net_1));
    CFG3 #( .INIT(8'hF2) )  un1_mem_0_5_215 (.A(\mem_7_[6]_net_1 ), .B(
        N_480), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_215_i));
    SLE un1_mem_0_5_189_rs (.D(VCC_net_1), .CLK(un1_mem_0_5_79_net_1), 
        .EN(VCC_net_1), .ALn(un1_mem_0_5_189_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(VCC_net_1), .Q(
        un1_mem_0_5_189_rs_net_1));
    CFG2 #( .INIT(4'h8) )  mem_14__1_sqmuxa_0_a2 (.A(N_482), .B(
        wr_enable), .Y(mem_14__1_sqmuxa));
    CFG1 #( .INIT(2'h1) )  un1_mem_0_5_102_set_RNO (.A(
        un1_mem_0_5_102_net_1), .Y(un1_mem_0_5_102_i));
    SLE un1_mem_0_5_170_rs (.D(VCC_net_1), .CLK(un1_mem_0_5_11_net_1), 
        .EN(VCC_net_1), .ALn(un1_mem_0_5_170_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(VCC_net_1), .Q(
        un1_mem_0_5_170_rs_net_1));
    CFG1 #( .INIT(2'h1) )  un1_mem_0_5_39_set_RNO (.A(
        un1_mem_0_5_39_net_1), .Y(un1_mem_0_5_39_i));
    CFG4 #( .INIT(16'h7350) )  \temp_data_2_15_i_1[4]  (.A(
        \mem_11_[4]_net_1 ), .B(\mem_3_[4]_net_1 ), .C(N_475), .D(
        N_470), .Y(\temp_data_2_15_i_1[4]_net_1 ));
    CFG1 #( .INIT(2'h1) )  un1_mem_0_5_set_RNO (.A(un1_mem_0_5_net_1), 
        .Y(un1_mem_0_5_i));
    SLE \mem_5_[6]  (.D(CoreAPB3_0_APBmslave2_PWDATA[6]), .CLK(
        FCCC_0_GL1), .EN(mem_5__1_sqmuxa), .ALn(un1_mem_0_5_184_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_5_rs[6] ));
    CFG3 #( .INIT(8'h02) )  un1_mem_0_5_28 (.A(\mem_2_[1]_net_1 ), .B(
        N_478), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_28_net_1));
    CFG3 #( .INIT(8'h02) )  un1_mem_0_5_43 (.A(\mem_1_[3]_net_1 ), .B(
        N_481), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_43_net_1));
    SLE un1_mem_0_5_119_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_14__1_sqmuxa), .ALn(un1_mem_0_5_119_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_mem_0_5_119_set_net_1));
    SLE \mem_15_[7]  (.D(CoreAPB3_0_APBmslave2_PWDATA[7]), .CLK(
        FCCC_0_GL1), .EN(mem_15__1_sqmuxa), .ALn(un1_mem_0_5_252_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_15_rs[7] ));
    CFG3 #( .INIT(8'h02) )  un1_mem_0_5_29 (.A(\mem_6_[0]_net_1 ), .B(
        N_468), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_29_net_1));
    CFG3 #( .INIT(8'hF2) )  un1_mem_0_5_228 (.A(\mem_12_[4]_net_1 ), 
        .B(N_469), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_228_i));
    SLE un1_mem_0_5_143_rs (.D(VCC_net_1), .CLK(un1_mem_0_5_24_net_1), 
        .EN(VCC_net_1), .ALn(un1_mem_0_5_143_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(VCC_net_1), .Q(
        un1_mem_0_5_143_rs_net_1));
    SLE un1_mem_0_5_117_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_14__1_sqmuxa), .ALn(un1_mem_0_5_117_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_mem_0_5_117_set_net_1));
    CFG1 #( .INIT(2'h1) )  un1_mem_0_5_49_set_RNO (.A(
        un1_mem_0_5_49_net_1), .Y(un1_mem_0_5_49_i));
    SLE un1_mem_0_5_19_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_12__1_sqmuxa), .ALn(un1_mem_0_5_19_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_mem_0_5_19_set_net_1));
    CFG3 #( .INIT(8'hF8) )  un1_mem_0_5_186_rs_RNI5E981 (.A(
        un1_mem_0_5_27_set_net_1), .B(un1_mem_0_5_186_rs_net_1), .C(
        \mem_5_rs[7] ), .Y(\mem_5_[7]_net_1 ));
    CFG1 #( .INIT(2'h1) )  un1_mem_0_5_12_set_RNO (.A(
        un1_mem_0_5_12_net_1), .Y(un1_mem_0_5_12_i));
    CFG1 #( .INIT(2'h1) )  un1_mem_0_5_119_set_RNO (.A(
        un1_mem_0_5_119_net_1), .Y(un1_mem_0_5_119_i));
    CFG3 #( .INIT(8'h02) )  un1_mem_0_5_58 (.A(\mem_15_[4]_net_1 ), .B(
        N_474), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_58_net_1));
    SLE \mem_12_[5]  (.D(CoreAPB3_0_APBmslave2_PWDATA[5]), .CLK(
        FCCC_0_GL1), .EN(mem_12__1_sqmuxa), .ALn(un1_mem_0_5_229_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_12_rs[5] ));
    CFG4 #( .INIT(16'h0080) )  \WRITE_GEN.mem_13__2_i_a2[5]  (.A(
        CoreAPB3_0_APBmslave2_PADDR[3]), .B(
        CoreAPB3_0_APBmslave2_PADDR[2]), .C(
        CoreAPB3_0_APBmslave2_PADDR[0]), .D(
        CoreAPB3_0_APBmslave2_PADDR[1]), .Y(N_477));
    CFG3 #( .INIT(8'hF8) )  un1_mem_0_5_137_rs_RNIHDC41 (.A(
        un1_mem_0_5_12_set_net_1), .B(un1_mem_0_5_137_rs_net_1), .C(
        \mem_1_rs[1] ), .Y(\mem_1_[1]_net_1 ));
    CFG3 #( .INIT(8'hF2) )  un1_mem_0_5_178 (.A(\mem_5_[3]_net_1 ), .B(
        N_472), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_178_i));
    SLE \mem_13_[0]  (.D(CoreAPB3_0_APBmslave2_PWDATA[0]), .CLK(
        FCCC_0_GL1), .EN(mem_13__1_sqmuxa), .ALn(un1_mem_0_5_232_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_13_rs[0] ));
    SLE un1_mem_0_5_8_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_0__1_sqmuxa), .ALn(un1_mem_0_5_8_i), .ADn(GND_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_mem_0_5_8_set_net_1));
    CFG3 #( .INIT(8'h02) )  un1_mem_0_5_59 (.A(\mem_15_[1]_net_1 ), .B(
        N_474), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_59_net_1));
    CFG3 #( .INIT(8'hF2) )  un1_mem_0_5_229 (.A(\mem_12_[5]_net_1 ), 
        .B(N_469), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_229_i));
    SLE un1_mem_0_5_212_rs (.D(VCC_net_1), .CLK(un1_mem_0_5_91_net_1), 
        .EN(VCC_net_1), .ALn(un1_mem_0_5_212_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(VCC_net_1), .Q(
        un1_mem_0_5_212_rs_net_1));
    CFG4 #( .INIT(16'hFFFE) )  \temp_data_2_15_i_12[7]  (.A(
        \temp_data_2_15_i_3[7]_net_1 ), .B(
        \temp_data_2_15_i_2[7]_net_1 ), .C(
        \temp_data_2_15_i_1[7]_net_1 ), .D(
        \temp_data_2_15_i_0[7]_net_1 ), .Y(
        \temp_data_2_15_i_12[7]_net_1 ));
    SLE un1_mem_0_5_121_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_6__1_sqmuxa), .ALn(un1_mem_0_5_121_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_mem_0_5_121_set_net_1));
    SLE un1_mem_0_5_58_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_15__1_sqmuxa), .ALn(un1_mem_0_5_58_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_mem_0_5_58_set_net_1));
    SLE un1_mem_0_5_30_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_2__1_sqmuxa), .ALn(un1_mem_0_5_30_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_mem_0_5_30_set_net_1));
    SLE un1_mem_0_5_79_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_9__1_sqmuxa), .ALn(un1_mem_0_5_79_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_mem_0_5_79_set_net_1));
    CFG3 #( .INIT(8'hF8) )  \mem_10__RNILCFV[2]  (.A(
        un1_mem_0_5_99_set_net_1), .B(un1_mem_0_5_195_rs_net_1), .C(
        \mem_10_rs[2] ), .Y(\mem_10_[2]_net_1 ));
    CFG3 #( .INIT(8'h02) )  un1_mem_0_5_76 (.A(\mem_9_[4]_net_1 ), .B(
        N_467), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_76_net_1));
    SLE un1_mem_0_5_155_rs (.D(VCC_net_1), .CLK(un1_mem_0_5_48_net_1), 
        .EN(VCC_net_1), .ALn(un1_mem_0_5_155_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(VCC_net_1), .Q(
        un1_mem_0_5_155_rs_net_1));
    CFG3 #( .INIT(8'hF8) )  \mem_2__RNIJLTN[2]  (.A(
        un1_mem_0_5_30_set_net_1), .B(un1_mem_0_5_146_rs_net_1), .C(
        \mem_2_rs[2] ), .Y(\mem_2_[2]_net_1 ));
    SLE un1_mem_0_5_201_rs (.D(VCC_net_1), .CLK(un1_mem_0_5_102_net_1), 
        .EN(VCC_net_1), .ALn(un1_mem_0_5_201_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(VCC_net_1), .Q(
        un1_mem_0_5_201_rs_net_1));
    SLE \mem_12_[1]  (.D(CoreAPB3_0_APBmslave2_PWDATA[1]), .CLK(
        FCCC_0_GL1), .EN(mem_12__1_sqmuxa), .ALn(un1_mem_0_5_224_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_12_rs[1] ));
    SLE un1_mem_0_5_151_rs (.D(VCC_net_1), .CLK(un1_mem_0_5_120_net_1), 
        .EN(VCC_net_1), .ALn(un1_mem_0_5_151_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(VCC_net_1), .Q(
        un1_mem_0_5_151_rs_net_1));
    CFG3 #( .INIT(8'h02) )  un1_mem_0_5_122 (.A(\mem_3_[0]_net_1 ), .B(
        N_470), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_122_net_1));
    SLE un1_mem_0_5_105_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_13__1_sqmuxa), .ALn(un1_mem_0_5_105_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_mem_0_5_105_set_net_1));
    SLE \mem_11_[0]  (.D(CoreAPB3_0_APBmslave2_PWDATA[0]), .CLK(
        FCCC_0_GL1), .EN(mem_11__1_sqmuxa), .ALn(un1_mem_0_5_207_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_11_rs[0] ));
    CFG1 #( .INIT(2'h1) )  un1_mem_0_5_30_set_RNO (.A(
        un1_mem_0_5_30_net_1), .Y(un1_mem_0_5_30_i));
    CFG3 #( .INIT(8'h02) )  un1_mem_0_5_40 (.A(\mem_5_[2]_net_1 ), .B(
        N_472), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_40_net_1));
    CFG3 #( .INIT(8'hF8) )  un1_mem_0_5_164_rs_RNI9DOL (.A(
        un1_mem_0_5_6_set_net_1), .B(un1_mem_0_5_164_rs_net_1), .C(
        \mem_4_rs[3] ), .Y(\mem_4_[3]_net_1 ));
    SLE un1_mem_0_5_120_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_2__1_sqmuxa), .ALn(un1_mem_0_5_120_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_mem_0_5_120_set_net_1));
    CFG3 #( .INIT(8'hF8) )  \mem_6__RNI5OVQ[4]  (.A(
        un1_mem_0_5_37_set_net_1), .B(un1_mem_0_5_196_rs_net_1), .C(
        \mem_6_rs[4] ), .Y(\mem_6_[4]_net_1 ));
    CFG1 #( .INIT(2'h1) )  un1_mem_0_5_76_set_RNO (.A(
        un1_mem_0_5_76_net_1), .Y(un1_mem_0_5_76_i));
    SLE un1_mem_0_5_205_rs (.D(VCC_net_1), .CLK(un1_mem_0_5_100_net_1), 
        .EN(VCC_net_1), .ALn(un1_mem_0_5_205_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(VCC_net_1), .Q(
        un1_mem_0_5_205_rs_net_1));
    CFG2 #( .INIT(4'h8) )  mem_5__1_sqmuxa_0_a2 (.A(N_472), .B(
        wr_enable), .Y(mem_5__1_sqmuxa));
    SLE \mem_3_[7]  (.D(CoreAPB3_0_APBmslave2_PWDATA[7]), .CLK(
        FCCC_0_GL1), .EN(mem_3__1_sqmuxa), .ALn(un1_mem_0_5_160_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_3_rs[7] ));
    SLE \mem_7_[4]  (.D(CoreAPB3_0_APBmslave2_PWDATA[4]), .CLK(
        FCCC_0_GL1), .EN(mem_7__1_sqmuxa), .ALn(un1_mem_0_5_158_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_7_rs[4] ));
    CFG1 #( .INIT(2'h1) )  un1_mem_0_5_109_set_RNO (.A(
        un1_mem_0_5_109_net_1), .Y(un1_mem_0_5_109_i));
    CFG1 #( .INIT(2'h1) )  un1_mem_0_5_78_set_RNO (.A(
        un1_mem_0_5_78_net_1), .Y(un1_mem_0_5_78_i));
    SLE un1_mem_0_5_184_rs (.D(VCC_net_1), .CLK(un1_mem_0_5_25_net_1), 
        .EN(VCC_net_1), .ALn(un1_mem_0_5_184_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(VCC_net_1), .Q(
        un1_mem_0_5_184_rs_net_1));
    SLE un1_mem_0_5_89_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_11__1_sqmuxa), .ALn(un1_mem_0_5_89_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_mem_0_5_89_set_net_1));
    SLE un1_mem_0_5_94_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_11__1_sqmuxa), .ALn(un1_mem_0_5_94_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_mem_0_5_94_set_net_1));
    CFG3 #( .INIT(8'hF8) )  un1_mem_0_5_78_set_RNIFTT11 (.A(
        un1_mem_0_5_78_set_net_1), .B(un1_mem_0_5_187_rs_net_1), .C(
        \mem_9_rs[6] ), .Y(\mem_9_[6]_net_1 ));
    CFG3 #( .INIT(8'hF8) )  un1_mem_0_5_178_rs_RNIV1V51 (.A(
        un1_mem_0_5_42_set_net_1), .B(un1_mem_0_5_178_rs_net_1), .C(
        \mem_5_rs[3] ), .Y(\mem_5_[3]_net_1 ));
    CFG3 #( .INIT(8'hF2) )  un1_mem_0_5_161 (.A(\mem_4_[0]_net_1 ), .B(
        N_476), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_161_i));
    SLE \mem_2_[4]  (.D(CoreAPB3_0_APBmslave2_PWDATA[4]), .CLK(
        FCCC_0_GL1), .EN(mem_2__1_sqmuxa), .ALn(un1_mem_0_5_148_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_2_rs[4] ));
    CFG1 #( .INIT(2'h1) )  un1_mem_0_5_40_set_RNO (.A(
        un1_mem_0_5_40_net_1), .Y(un1_mem_0_5_40_i));
    SLE \mem_3_[5]  (.D(CoreAPB3_0_APBmslave2_PWDATA[5]), .CLK(
        FCCC_0_GL1), .EN(mem_3__1_sqmuxa), .ALn(un1_mem_0_5_157_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_3_rs[5] ));
    SLE un1_mem_0_5_24_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_1__1_sqmuxa), .ALn(un1_mem_0_5_24_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_mem_0_5_24_set_net_1));
    CFG3 #( .INIT(8'hF8) )  \mem_6__RNI3P1N[0]  (.A(
        un1_mem_0_5_29_set_net_1), .B(un1_mem_0_5_188_rs_net_1), .C(
        \mem_6_rs[0] ), .Y(\mem_6_[0]_net_1 ));
    SLE un1_mem_0_5_129_rs (.D(VCC_net_1), .CLK(un1_mem_0_5_82_net_1), 
        .EN(VCC_net_1), .ALn(un1_mem_0_5_129_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(VCC_net_1), .Q(
        un1_mem_0_5_129_rs_net_1));
    CFG4 #( .INIT(16'hFFFE) )  \temp_data_2_15_i_12[2]  (.A(
        \temp_data_2_15_i_3[2]_net_1 ), .B(
        \temp_data_2_15_i_2[2]_net_1 ), .C(
        \temp_data_2_15_i_1[2]_net_1 ), .D(
        \temp_data_2_15_i_0[2]_net_1 ), .Y(
        \temp_data_2_15_i_12[2]_net_1 ));
    CFG2 #( .INIT(4'h2) )  \temp_data_2_15_i_a2_13[7]  (.A(N_476), .B(
        \mem_4_[7]_net_1 ), .Y(N_455));
    CFG3 #( .INIT(8'hF8) )  un1_mem_0_5_58_set_RNIIPAE (.A(
        un1_mem_0_5_58_set_net_1), .B(un1_mem_0_5_253_rs_net_1), .C(
        \mem_15_rs[4] ), .Y(\mem_15_[4]_net_1 ));
    CFG3 #( .INIT(8'h02) )  un1_mem_0_5_25 (.A(\mem_5_[6]_net_1 ), .B(
        N_472), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_25_net_1));
    CFG3 #( .INIT(8'hF2) )  un1_mem_0_5_223 (.A(\mem_8_[2]_net_1 ), .B(
        N_479), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_223_i));
    CFG3 #( .INIT(8'h02) )  un1_mem_0_5_81 (.A(\mem_0_[1]_net_1 ), .B(
        N_473), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_81_net_1));
    CFG3 #( .INIT(8'hF2) )  un1_mem_0_5_188 (.A(\mem_6_[0]_net_1 ), .B(
        N_468), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_188_i));
    CFG4 #( .INIT(16'h7350) )  \temp_data_2_15_i_5[0]  (.A(
        \mem_7_[0]_net_1 ), .B(\mem_5_[0]_net_1 ), .C(N_480), .D(N_472)
        , .Y(\temp_data_2_15_i_5[0]_net_1 ));
    SLE \mem_4_[4]  (.D(CoreAPB3_0_APBmslave2_PWDATA[4]), .CLK(
        FCCC_0_GL1), .EN(mem_4__1_sqmuxa), .ALn(un1_mem_0_5_165_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_4_rs[4] ));
    CFG3 #( .INIT(8'hF8) )  \mem_11__RNID3DK[5]  (.A(
        un1_mem_0_5_93_set_net_1), .B(un1_mem_0_5_216_rs_net_1), .C(
        \mem_11_rs[5] ), .Y(\mem_11_[5]_net_1 ));
    CFG3 #( .INIT(8'hF2) )  un1_mem_0_5_198 (.A(\mem_6_[5]_net_1 ), .B(
        N_468), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_198_i));
    SLE un1_mem_0_5_133_rs (.D(VCC_net_1), .CLK(un1_mem_0_5_86_net_1), 
        .EN(VCC_net_1), .ALn(un1_mem_0_5_133_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(VCC_net_1), .Q(
        un1_mem_0_5_133_rs_net_1));
    CFG4 #( .INIT(16'h7530) )  \temp_data_2_15_i_0[6]  (.A(
        \mem_9_[6]_net_1 ), .B(\mem_1_[6]_net_1 ), .C(N_481), .D(N_467)
        , .Y(\temp_data_2_15_i_0[6]_net_1 ));
    SLE un1_mem_0_5_127_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_7__1_sqmuxa), .ALn(un1_mem_0_5_127_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_mem_0_5_127_set_net_1));
    CFG2 #( .INIT(4'h8) )  mem_12__1_sqmuxa_0_a2 (.A(N_469), .B(
        wr_enable), .Y(mem_12__1_sqmuxa));
    CFG3 #( .INIT(8'h02) )  un1_mem_0_5_92 (.A(\mem_11_[4]_net_1 ), .B(
        N_475), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_92_net_1));
    SLE un1_mem_0_5_152_rs (.D(VCC_net_1), .CLK(un1_mem_0_5_122_net_1), 
        .EN(VCC_net_1), .ALn(un1_mem_0_5_152_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(VCC_net_1), .Q(
        un1_mem_0_5_152_rs_net_1));
    SLE un1_mem_0_5_68_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_8__1_sqmuxa), .ALn(un1_mem_0_5_68_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_mem_0_5_68_set_net_1));
    SLE un1_mem_0_5_159_rs (.D(VCC_net_1), .CLK(un1_mem_0_5_83_net_1), 
        .EN(VCC_net_1), .ALn(un1_mem_0_5_159_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(VCC_net_1), .Q(
        un1_mem_0_5_159_rs_net_1));
    CFG3 #( .INIT(8'hF8) )  un1_mem_0_5_109_set_RNI0KRF (.A(
        un1_mem_0_5_109_set_net_1), .B(un1_mem_0_5_237_rs_net_1), .C(
        \mem_13_rs[5] ), .Y(\mem_13_[5]_net_1 ));
    CFG1 #( .INIT(2'h1) )  un1_mem_0_5_53_set_RNO (.A(
        un1_mem_0_5_53_net_1), .Y(un1_mem_0_5_53_i));
    CFG3 #( .INIT(8'h02) )  un1_mem_0_5_24 (.A(\mem_1_[7]_net_1 ), .B(
        N_481), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_24_net_1));
    CFG2 #( .INIT(4'h2) )  \temp_data_2_15_i_a2_13[2]  (.A(N_476), .B(
        \mem_4_[2]_net_1 ), .Y(N_361));
    CFG3 #( .INIT(8'h02) )  un1_mem_0_5_55 (.A(\mem_3_[7]_net_1 ), .B(
        N_470), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_55_net_1));
    CFG4 #( .INIT(16'h7350) )  \temp_data_2_15_i_2[1]  (.A(
        \mem_13_[1]_net_1 ), .B(\mem_15_[1]_net_1 ), .C(N_477), .D(
        N_474), .Y(\temp_data_2_15_i_2[1]_net_1 ));
    SLE \mem_10_[4]  (.D(CoreAPB3_0_APBmslave2_PWDATA[4]), .CLK(
        FCCC_0_GL1), .EN(mem_10__1_sqmuxa), .ALn(un1_mem_0_5_199_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_10_rs[4] ));
    CFG1 #( .INIT(2'h1) )  un1_mem_0_5_21_set_RNO (.A(
        un1_mem_0_5_21_net_1), .Y(un1_mem_0_5_21_i));
    CFG3 #( .INIT(8'hF8) )  un1_mem_0_5_62_set_RNIFAJG (.A(
        un1_mem_0_5_62_set_net_1), .B(un1_mem_0_5_254_rs_net_1), .C(
        \mem_15_rs[5] ), .Y(\mem_15_[5]_net_1 ));
    SLE \mem_7_[0]  (.D(CoreAPB3_0_APBmslave2_PWDATA[0]), .CLK(
        FCCC_0_GL1), .EN(mem_7__1_sqmuxa), .ALn(un1_mem_0_5_204_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_7_rs[0] ));
    SLE un1_mem_0_5_195_rs (.D(VCC_net_1), .CLK(un1_mem_0_5_99_net_1), 
        .EN(VCC_net_1), .ALn(un1_mem_0_5_195_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(VCC_net_1), .Q(
        un1_mem_0_5_195_rs_net_1));
    SLE un1_mem_0_5_5_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_8__1_sqmuxa), .ALn(un1_mem_0_5_5_i), .ADn(GND_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_mem_0_5_5_set_net_1));
    CFG1 #( .INIT(2'h1) )  un1_mem_0_5_72_set_RNO (.A(
        un1_mem_0_5_72_net_1), .Y(un1_mem_0_5_72_i));
    SLE \mem_14_[2]  (.D(CoreAPB3_0_APBmslave2_PWDATA[2]), .CLK(
        FCCC_0_GL1), .EN(mem_14__1_sqmuxa), .ALn(un1_mem_0_5_242_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_14_rs[2] ));
    CFG1 #( .INIT(2'h1) )  un1_mem_0_5_67_set_RNO (.A(
        un1_mem_0_5_67_net_1), .Y(un1_mem_0_5_67_i));
    SLE \mem_2_[0]  (.D(CoreAPB3_0_APBmslave2_PWDATA[0]), .CLK(
        FCCC_0_GL1), .EN(mem_2__1_sqmuxa), .ALn(un1_mem_0_5_144_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_2_rs[0] ));
    SLE un1_mem_0_5_191_rs (.D(VCC_net_1), .CLK(un1_mem_0_5_97_net_1), 
        .EN(VCC_net_1), .ALn(un1_mem_0_5_191_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(VCC_net_1), .Q(
        un1_mem_0_5_191_rs_net_1));
    CFG3 #( .INIT(8'h02) )  un1_mem_0_5_32 (.A(\mem_2_[3]_net_1 ), .B(
        N_478), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_32_net_1));
    CFG4 #( .INIT(16'h7350) )  \temp_data_2_15_i_3[6]  (.A(
        \mem_14_[6]_net_1 ), .B(\mem_2_[6]_net_1 ), .C(N_482), .D(
        N_478), .Y(\temp_data_2_15_i_3[6]_net_1 ));
    CFG3 #( .INIT(8'hF2) )  un1_mem_0_5_212 (.A(\mem_11_[3]_net_1 ), 
        .B(N_475), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_212_i));
    CFG4 #( .INIT(16'h7350) )  \temp_data_2_15_i_1[0]  (.A(
        \mem_11_[0]_net_1 ), .B(\mem_3_[0]_net_1 ), .C(N_475), .D(
        N_470), .Y(\temp_data_2_15_i_1[0]_net_1 ));
    SLE un1_mem_0_5_32_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_2__1_sqmuxa), .ALn(un1_mem_0_5_32_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_mem_0_5_32_set_net_1));
    CFG1 #( .INIT(2'h1) )  un1_mem_0_5_65_set_RNO (.A(
        un1_mem_0_5_65_net_1), .Y(un1_mem_0_5_65_i));
    SLE un1_mem_0_5_221_rs (.D(VCC_net_1), .CLK(un1_mem_0_5_5_net_1), 
        .EN(VCC_net_1), .ALn(un1_mem_0_5_221_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(VCC_net_1), .Q(
        un1_mem_0_5_221_rs_net_1));
    CFG3 #( .INIT(8'h02) )  un1_mem_0_5_54 (.A(\mem_7_[5]_net_1 ), .B(
        N_480), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_54_net_1));
    SLE \mem_4_[0]  (.D(CoreAPB3_0_APBmslave2_PWDATA[0]), .CLK(
        FCCC_0_GL1), .EN(mem_4__1_sqmuxa), .ALn(un1_mem_0_5_161_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_4_rs[0] ));
    SLE \mem_10_[6]  (.D(CoreAPB3_0_APBmslave2_PWDATA[6]), .CLK(
        FCCC_0_GL1), .EN(mem_10__1_sqmuxa), .ALn(un1_mem_0_5_203_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_10_rs[6] ));
    CFG3 #( .INIT(8'h02) )  un1_mem_0_5_23 (.A(\mem_12_[7]_net_1 ), .B(
        N_469), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_23_net_1));
    SLE un1_mem_0_5_116_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_14__1_sqmuxa), .ALn(un1_mem_0_5_116_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_mem_0_5_116_set_net_1));
    CFG4 #( .INIT(16'hFFFE) )  \temp_data_2_15_i_12[5]  (.A(
        \temp_data_2_15_i_3[5]_net_1 ), .B(
        \temp_data_2_15_i_2[5]_net_1 ), .C(
        \temp_data_2_15_i_1[5]_net_1 ), .D(
        \temp_data_2_15_i_0[5]_net_1 ), .Y(
        \temp_data_2_15_i_12[5]_net_1 ));
    CFG3 #( .INIT(8'h02) )  un1_mem_0_5_6 (.A(\mem_4_[3]_net_1 ), .B(
        N_476), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_6_net_1));
    CFG4 #( .INIT(16'h7350) )  \temp_data_2_15_i_3[0]  (.A(
        \mem_14_[0]_net_1 ), .B(\mem_2_[0]_net_1 ), .C(N_482), .D(
        N_478), .Y(\temp_data_2_15_i_3[0]_net_1 ));
    SLE un1_mem_0_5_53_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_7__1_sqmuxa), .ALn(un1_mem_0_5_53_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_mem_0_5_53_set_net_1));
    CFG4 #( .INIT(16'h7350) )  \temp_data_2_15_i_1[2]  (.A(
        \mem_11_[2]_net_1 ), .B(\mem_3_[2]_net_1 ), .C(N_475), .D(
        N_470), .Y(\temp_data_2_15_i_1[2]_net_1 ));
    SLE un1_mem_0_5_225_rs (.D(VCC_net_1), .CLK(un1_mem_0_5_66_net_1), 
        .EN(VCC_net_1), .ALn(un1_mem_0_5_225_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(VCC_net_1), .Q(
        un1_mem_0_5_225_rs_net_1));
    SLE un1_mem_0_5_35_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_6__1_sqmuxa), .ALn(un1_mem_0_5_35_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_mem_0_5_35_set_net_1));
    CFG4 #( .INIT(16'hFFFE) )  \temp_data_2_15_i_12[3]  (.A(
        \temp_data_2_15_i_3[3]_net_1 ), .B(
        \temp_data_2_15_i_2[3]_net_1 ), .C(
        \temp_data_2_15_i_1[3]_net_1 ), .D(
        \temp_data_2_15_i_0[3]_net_1 ), .Y(
        \temp_data_2_15_i_12[3]_net_1 ));
    CFG4 #( .INIT(16'h7350) )  \temp_data_2_15_i_5[7]  (.A(
        \mem_7_[7]_net_1 ), .B(\mem_5_[7]_net_1 ), .C(N_480), .D(N_472)
        , .Y(\temp_data_2_15_i_5[7]_net_1 ));
    CFG3 #( .INIT(8'hF8) )  un1_mem_0_5_79_set_RNIJ8A81 (.A(
        un1_mem_0_5_79_set_net_1), .B(un1_mem_0_5_189_rs_net_1), .C(
        \mem_9_rs[7] ), .Y(\mem_9_[7]_net_1 ));
    SLE un1_mem_0_5_251_rs (.D(VCC_net_1), .CLK(un1_mem_0_5_61_net_1), 
        .EN(VCC_net_1), .ALn(un1_mem_0_5_251_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(VCC_net_1), .Q(
        un1_mem_0_5_251_rs_net_1));
    CFG3 #( .INIT(8'hF2) )  un1_mem_0_5_254 (.A(\mem_15_[5]_net_1 ), 
        .B(N_474), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_254_i));
    CFG3 #( .INIT(8'hF8) )  \mem_2__RNIN1DH[3]  (.A(
        un1_mem_0_5_32_set_net_1), .B(un1_mem_0_5_147_rs_net_1), .C(
        \mem_2_rs[3] ), .Y(\mem_2_[3]_net_1 ));
    SLE un1_mem_0_5_6_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_4__1_sqmuxa), .ALn(un1_mem_0_5_6_i), .ADn(GND_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_mem_0_5_6_set_net_1));
    CFG3 #( .INIT(8'h02) )  un1_mem_0_5_53 (.A(\mem_7_[4]_net_1 ), .B(
        N_480), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_53_net_1));
    SLE un1_mem_0_5_240_rs (.D(VCC_net_1), .CLK(un1_mem_0_5_112_net_1), 
        .EN(VCC_net_1), .ALn(un1_mem_0_5_240_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(VCC_net_1), .Q(
        un1_mem_0_5_240_rs_net_1));
    CFG3 #( .INIT(8'h02) )  un1_mem_0_5_11 (.A(\mem_4_[7]_net_1 ), .B(
        N_476), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_11_net_1));
    CFG3 #( .INIT(8'hF2) )  un1_mem_0_5_158 (.A(\mem_7_[4]_net_1 ), .B(
        N_480), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_158_i));
    CFG4 #( .INIT(16'h7350) )  \temp_data_2_15_i_3[2]  (.A(
        \mem_14_[2]_net_1 ), .B(\mem_2_[2]_net_1 ), .C(N_482), .D(
        N_478), .Y(\temp_data_2_15_i_3[2]_net_1 ));
    SLE un1_mem_0_5_255_rs (.D(VCC_net_1), .CLK(un1_mem_0_5_63_net_1), 
        .EN(VCC_net_1), .ALn(un1_mem_0_5_255_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(VCC_net_1), .Q(
        un1_mem_0_5_255_rs_net_1));
    CFG2 #( .INIT(4'h2) )  \temp_data_2_15_i_a2_13[3]  (.A(N_476), .B(
        \mem_4_[3]_net_1 ), .Y(N_377));
    CFG3 #( .INIT(8'h02) )  un1_mem_0_5_116 (.A(\mem_14_[4]_net_1 ), 
        .B(N_482), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_116_net_1));
    SLE un1_mem_0_5_192_rs (.D(VCC_net_1), .CLK(un1_mem_0_5_33_net_1), 
        .EN(VCC_net_1), .ALn(un1_mem_0_5_192_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(VCC_net_1), .Q(
        un1_mem_0_5_192_rs_net_1));
    CFG3 #( .INIT(8'h02) )  un1_mem_0_5_87 (.A(\mem_0_[6]_net_1 ), .B(
        N_473), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_87_net_1));
    SLE un1_mem_0_5_199_rs (.D(VCC_net_1), .CLK(un1_mem_0_5_101_net_1), 
        .EN(VCC_net_1), .ALn(un1_mem_0_5_199_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(VCC_net_1), .Q(
        un1_mem_0_5_199_rs_net_1));
    CFG4 #( .INIT(16'hEFEE) )  \temp_data_2_15_i_11[1]  (.A(N_345), .B(
        \temp_data_2_15_i_7[1]_net_1 ), .C(\mem_0_[1]_net_1 ), .D(
        N_473), .Y(\temp_data_2_15_i_11[1]_net_1 ));
    SLE un1_mem_0_5_57_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_15__1_sqmuxa), .ALn(un1_mem_0_5_57_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_mem_0_5_57_set_net_1));
    CFG3 #( .INIT(8'hF8) )  \mem_12__RNI3NVT[6]  (.A(
        un1_mem_0_5_22_set_net_1), .B(un1_mem_0_5_230_rs_net_1), .C(
        \mem_12_rs[6] ), .Y(\mem_12_[6]_net_1 ));
    SLE \data_out[4]  (.D(\temp_data[4]_net_1 ), .CLK(FCCC_0_GL1), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(
        CoreAPB3_0_APBmslave3_PRDATA[4]));
    CFG1 #( .INIT(2'h1) )  un1_mem_0_5_121_set_RNO (.A(
        un1_mem_0_5_121_net_1), .Y(un1_mem_0_5_121_i));
    SLE un1_mem_0_5_154_rs (.D(VCC_net_1), .CLK(un1_mem_0_5_126_net_1), 
        .EN(VCC_net_1), .ALn(un1_mem_0_5_154_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(VCC_net_1), .Q(
        un1_mem_0_5_154_rs_net_1));
    CFG2 #( .INIT(4'h8) )  mem_2__1_sqmuxa_0_a2 (.A(N_478), .B(
        wr_enable), .Y(mem_2__1_sqmuxa));
    CFG3 #( .INIT(8'hF2) )  un1_mem_0_5_244 (.A(\mem_14_[4]_net_1 ), 
        .B(N_482), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_244_i));
    CFG4 #( .INIT(16'h7350) )  \temp_data_2_15_i_2[0]  (.A(
        \mem_13_[0]_net_1 ), .B(\mem_15_[0]_net_1 ), .C(N_477), .D(
        N_474), .Y(\temp_data_2_15_i_2[0]_net_1 ));
    CFG1 #( .INIT(2'h1) )  un1_mem_0_5_69_set_RNO (.A(
        un1_mem_0_5_69_net_1), .Y(un1_mem_0_5_69_i));
    CFG1 #( .INIT(2'h1) )  un1_mem_0_5_4_set_RNO (.A(
        un1_mem_0_5_4_net_1), .Y(un1_mem_0_5_4_i));
    CFG1 #( .INIT(2'h1) )  un1_mem_0_5_9_set_RNO (.A(
        un1_mem_0_5_9_net_1), .Y(un1_mem_0_5_9_i));
    CFG1 #( .INIT(2'h1) )  un1_mem_0_5_116_set_RNO (.A(
        un1_mem_0_5_116_net_1), .Y(un1_mem_0_5_116_i));
    CFG4 #( .INIT(16'h0010) )  \WRITE_GEN.mem_1__2_i_a2[5]  (.A(
        CoreAPB3_0_APBmslave2_PADDR[3]), .B(
        CoreAPB3_0_APBmslave2_PADDR[2]), .C(
        CoreAPB3_0_APBmslave2_PADDR[0]), .D(
        CoreAPB3_0_APBmslave2_PADDR[1]), .Y(N_481));
    CFG4 #( .INIT(16'hFFFE) )  \temp_data_2_15_i_12[6]  (.A(
        \temp_data_2_15_i_3[6]_net_1 ), .B(
        \temp_data_2_15_i_2[6]_net_1 ), .C(
        \temp_data_2_15_i_1[6]_net_1 ), .D(
        \temp_data_2_15_i_0[6]_net_1 ), .Y(
        \temp_data_2_15_i_12[6]_net_1 ));
    CFG3 #( .INIT(8'hF2) )  un1_mem_0_5_148 (.A(\mem_2_[4]_net_1 ), .B(
        N_478), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_148_i));
    CFG1 #( .INIT(2'h1) )  un1_mem_0_5_54_set_RNO (.A(
        un1_mem_0_5_54_net_1), .Y(un1_mem_0_5_54_i));
    CFG3 #( .INIT(8'h02) )  un1_mem_0_5_20 (.A(\mem_12_[4]_net_1 ), .B(
        N_469), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_20_net_1));
    SLE \data_out[3]  (.D(\temp_data[3]_net_1 ), .CLK(FCCC_0_GL1), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(
        CoreAPB3_0_APBmslave3_PRDATA[3]));
    SLE un1_mem_0_5_188_rs (.D(VCC_net_1), .CLK(un1_mem_0_5_29_net_1), 
        .EN(VCC_net_1), .ALn(un1_mem_0_5_188_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(VCC_net_1), .Q(
        un1_mem_0_5_188_rs_net_1));
    SLE un1_mem_0_5_108_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_13__1_sqmuxa), .ALn(un1_mem_0_5_108_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_mem_0_5_108_set_net_1));
    CFG3 #( .INIT(8'hF8) )  un1_mem_0_5_181_rs_RNI3SOU (.A(
        un1_mem_0_5_75_set_net_1), .B(un1_mem_0_5_181_rs_net_1), .C(
        \mem_9_rs[3] ), .Y(\mem_9_[3]_net_1 ));
    SLE un1_mem_0_5_166_rs (.D(VCC_net_1), .CLK(un1_mem_0_5_67_net_1), 
        .EN(VCC_net_1), .ALn(un1_mem_0_5_166_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(VCC_net_1), .Q(
        un1_mem_0_5_166_rs_net_1));
    CFG3 #( .INIT(8'hF8) )  un1_mem_0_5_17_set_RNI59QO (.A(
        un1_mem_0_5_17_set_net_1), .B(un1_mem_0_5_224_rs_net_1), .C(
        \mem_12_rs[1] ), .Y(\mem_12_[1]_net_1 ));
    CFG2 #( .INIT(4'h2) )  \temp_data_2_15_i_a2_13[5]  (.A(N_476), .B(
        \mem_4_[5]_net_1 ), .Y(N_416));
    SLE un1_mem_0_5_56_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_15__1_sqmuxa), .ALn(un1_mem_0_5_56_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_mem_0_5_56_set_net_1));
    CFG3 #( .INIT(8'hF8) )  un1_mem_0_5_170_rs_RNIMMRL (.A(
        un1_mem_0_5_11_set_net_1), .B(un1_mem_0_5_170_rs_net_1), .C(
        \mem_4_rs[7] ), .Y(\mem_4_[7]_net_1 ));
    CFG2 #( .INIT(4'h2) )  \temp_data_2_15_i_a2_13[6]  (.A(N_476), .B(
        \mem_4_[6]_net_1 ), .Y(N_434));
    CFG3 #( .INIT(8'hF8) )  \mem_10__RNIH13P[1]  (.A(
        un1_mem_0_5_98_set_net_1), .B(un1_mem_0_5_193_rs_net_1), .C(
        \mem_10_rs[1] ), .Y(\mem_10_[1]_net_1 ));
    SLE un1_mem_0_5_63_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_15__1_sqmuxa), .ALn(un1_mem_0_5_63_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_mem_0_5_63_set_net_1));
    CFG1 #( .INIT(2'h1) )  un1_mem_0_5_36_set_RNO (.A(
        un1_mem_0_5_36_net_1), .Y(un1_mem_0_5_36_i));
    CFG4 #( .INIT(16'h0001) )  \temp_data_RNO[0]  (.A(
        \temp_data_2_15_i_4[0]_net_1 ), .B(
        \temp_data_2_15_i_5[0]_net_1 ), .C(
        \temp_data_2_15_i_11[0]_net_1 ), .D(
        \temp_data_2_15_i_12[0]_net_1 ), .Y(N_4_i_0));
    CFG2 #( .INIT(4'h2) )  \temp_data_2_15_i_a2_13[0]  (.A(N_476), .B(
        \mem_4_[0]_net_1 ), .Y(N_329));
    CFG3 #( .INIT(8'hF2) )  un1_mem_0_5_162 (.A(\mem_4_[1]_net_1 ), .B(
        N_476), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_162_i));
    SLE un1_mem_0_5_126_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_3__1_sqmuxa), .ALn(un1_mem_0_5_126_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_mem_0_5_126_set_net_1));
    CFG1 #( .INIT(2'h1) )  un1_mem_0_5_38_set_RNO (.A(
        un1_mem_0_5_38_net_1), .Y(un1_mem_0_5_38_i));
    SLE un1_mem_0_5_243_rs (.D(VCC_net_1), .CLK(un1_mem_0_5_115_net_1), 
        .EN(VCC_net_1), .ALn(un1_mem_0_5_243_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(VCC_net_1), .Q(
        un1_mem_0_5_243_rs_net_1));
    CFG3 #( .INIT(8'hF2) )  un1_mem_0_5_234 (.A(\mem_13_[2]_net_1 ), 
        .B(N_477), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_234_i));
    CFG3 #( .INIT(8'h02) )  un1_mem_0_5_50 (.A(\mem_3_[4]_net_1 ), .B(
        N_470), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_50_net_1));
    CFG3 #( .INIT(8'hF2) )  un1_mem_0_5_255 (.A(\mem_15_[6]_net_1 ), 
        .B(N_474), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_255_i));
    CFG3 #( .INIT(8'hF8) )  \mem_2__RNIQB2N[6]  (.A(
        un1_mem_0_5_38_set_net_1), .B(un1_mem_0_5_150_rs_net_1), .C(
        \mem_2_rs[6] ), .Y(\mem_2_[6]_net_1 ));
    SLE \mem_8_[2]  (.D(CoreAPB3_0_APBmslave2_PWDATA[2]), .CLK(
        FCCC_0_GL1), .EN(mem_8__1_sqmuxa), .ALn(un1_mem_0_5_223_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_8_rs[2] ));
    CFG3 #( .INIT(8'hF2) )  un1_mem_0_5_138 (.A(\mem_1_[2]_net_1 ), .B(
        N_481), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_138_i));
    CFG1 #( .INIT(2'h1) )  un1_mem_0_5_106_set_RNO (.A(
        un1_mem_0_5_106_net_1), .Y(un1_mem_0_5_106_i));
    CFG4 #( .INIT(16'hEFEE) )  \temp_data_2_15_i_11[5]  (.A(N_416), .B(
        \temp_data_2_15_i_7[5]_net_1 ), .C(\mem_0_[5]_net_1 ), .D(
        N_473), .Y(\temp_data_2_15_i_11[5]_net_1 ));
    SLE \mem_6_[7]  (.D(CoreAPB3_0_APBmslave2_PWDATA[7]), .CLK(
        FCCC_0_GL1), .EN(mem_6__1_sqmuxa), .ALn(un1_mem_0_5_202_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_6_rs[7] ));
    CFG1 #( .INIT(2'h1) )  un1_mem_0_5_46_set_RNO (.A(
        un1_mem_0_5_46_net_1), .Y(un1_mem_0_5_46_i));
    SLE un1_mem_0_5_176_rs (.D(VCC_net_1), .CLK(un1_mem_0_5_40_net_1), 
        .EN(VCC_net_1), .ALn(un1_mem_0_5_176_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(VCC_net_1), .Q(
        un1_mem_0_5_176_rs_net_1));
    SLE \mem_14_[7]  (.D(CoreAPB3_0_APBmslave2_PWDATA[7]), .CLK(
        FCCC_0_GL1), .EN(mem_14__1_sqmuxa), .ALn(un1_mem_0_5_247_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_14_rs[7] ));
    CFG3 #( .INIT(8'h02) )  un1_mem_0_5_88 (.A(\mem_11_[0]_net_1 ), .B(
        N_475), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_88_net_1));
    CFG3 #( .INIT(8'hF8) )  \mem_10__RNIHJPE[7]  (.A(
        un1_mem_0_5_100_set_net_1), .B(un1_mem_0_5_205_rs_net_1), .C(
        \mem_10_rs[7] ), .Y(\mem_10_[7]_net_1 ));
    CFG2 #( .INIT(4'h8) )  mem_3__1_sqmuxa_0_a2 (.A(N_470), .B(
        wr_enable), .Y(mem_3__1_sqmuxa));
    CFG1 #( .INIT(2'h1) )  un1_mem_0_5_48_set_RNO (.A(
        un1_mem_0_5_48_net_1), .Y(un1_mem_0_5_48_i));
    SLE \mem_6_[5]  (.D(CoreAPB3_0_APBmslave2_PWDATA[5]), .CLK(
        FCCC_0_GL1), .EN(mem_6__1_sqmuxa), .ALn(un1_mem_0_5_198_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_6_rs[5] ));
    CFG3 #( .INIT(8'h02) )  un1_mem_0_5_89 (.A(\mem_11_[1]_net_1 ), .B(
        N_475), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_89_net_1));
    SLE un1_mem_0_5_39_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_6__1_sqmuxa), .ALn(un1_mem_0_5_39_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_mem_0_5_39_set_net_1));
    SLE \mem_15_[5]  (.D(CoreAPB3_0_APBmslave2_PWDATA[5]), .CLK(
        FCCC_0_GL1), .EN(mem_15__1_sqmuxa), .ALn(un1_mem_0_5_254_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_15_rs[5] ));
    SLE un1_mem_0_5_147_rs (.D(VCC_net_1), .CLK(un1_mem_0_5_32_net_1), 
        .EN(VCC_net_1), .ALn(un1_mem_0_5_147_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(VCC_net_1), .Q(
        un1_mem_0_5_147_rs_net_1));
    CFG1 #( .INIT(2'h1) )  un1_mem_0_5_60_set_RNO (.A(
        un1_mem_0_5_60_net_1), .Y(un1_mem_0_5_60_i));
    CFG3 #( .INIT(8'hF8) )  un1_mem_0_5_233_rs_RNIKJMA1 (.A(
        un1_mem_0_5_105_set_net_1), .B(un1_mem_0_5_233_rs_net_1), .C(
        \mem_13_rs[1] ), .Y(\mem_13_[1]_net_1 ));
    SLE un1_mem_0_5_98_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_10__1_sqmuxa), .ALn(un1_mem_0_5_98_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_mem_0_5_98_set_net_1));
    CFG3 #( .INIT(8'hF2) )  un1_mem_0_5_245 (.A(\mem_14_[5]_net_1 ), 
        .B(N_482), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_245_i));
    SLE un1_mem_0_5_67_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_4__1_sqmuxa), .ALn(un1_mem_0_5_67_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_mem_0_5_67_set_net_1));
    CFG4 #( .INIT(16'hEFEE) )  \temp_data_2_15_i_11[6]  (.A(N_434), .B(
        \temp_data_2_15_i_7[6]_net_1 ), .C(\mem_0_[6]_net_1 ), .D(
        N_473), .Y(\temp_data_2_15_i_11[6]_net_1 ));
    SLE \mem_0_[7]  (.D(CoreAPB3_0_APBmslave2_PWDATA[7]), .CLK(
        FCCC_0_GL1), .EN(mem_0__1_sqmuxa), .ALn(un1_mem_0_5_135_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_0_rs[7] ));
    SLE un1_mem_0_5_28_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_2__1_sqmuxa), .ALn(un1_mem_0_5_28_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_mem_0_5_28_set_net_1));
    SLE un1_mem_0_5_230_rs (.D(VCC_net_1), .CLK(un1_mem_0_5_22_net_1), 
        .EN(VCC_net_1), .ALn(un1_mem_0_5_230_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(VCC_net_1), .Q(
        un1_mem_0_5_230_rs_net_1));
    CFG3 #( .INIT(8'hF2) )  un1_mem_0_5_210 (.A(\mem_7_[3]_net_1 ), .B(
        N_480), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_210_i));
    SLE un1_mem_0_5_219_rs (.D(VCC_net_1), .CLK(un1_mem_0_5_7_net_1), 
        .EN(VCC_net_1), .ALn(un1_mem_0_5_219_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(VCC_net_1), .Q(
        un1_mem_0_5_219_rs_net_1));
    CFG3 #( .INIT(8'h02) )  un1_mem_0_5_71 (.A(\mem_8_[7]_net_1 ), .B(
        N_479), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_71_net_1));
    SLE un1_mem_0_5_9_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_4__1_sqmuxa), .ALn(un1_mem_0_5_9_i), .ADn(GND_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_mem_0_5_9_set_net_1));
    CFG3 #( .INIT(8'hF8) )  un1_mem_0_5_239_rs_RNIT0RQ (.A(
        un1_mem_0_5_111_set_net_1), .B(un1_mem_0_5_239_rs_net_1), .C(
        \mem_13_rs[7] ), .Y(\mem_13_[7]_net_1 ));
    CFG3 #( .INIT(8'hF8) )  un1_mem_0_5_92_set_RNI9O0E (.A(
        un1_mem_0_5_92_set_net_1), .B(un1_mem_0_5_214_rs_net_1), .C(
        \mem_11_rs[4] ), .Y(\mem_11_[4]_net_1 ));
    SLE un1_mem_0_5_194_rs (.D(VCC_net_1), .CLK(un1_mem_0_5_35_net_1), 
        .EN(VCC_net_1), .ALn(un1_mem_0_5_194_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(VCC_net_1), .Q(
        un1_mem_0_5_194_rs_net_1));
    CFG3 #( .INIT(8'h02) )  un1_mem_0_5_96 (.A(\mem_10_[3]_net_1 ), .B(
        N_471), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_96_net_1));
    SLE \mem_0_[5]  (.D(CoreAPB3_0_APBmslave2_PWDATA[5]), .CLK(
        FCCC_0_GL1), .EN(mem_0__1_sqmuxa), .ALn(un1_mem_0_5_133_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_0_rs[5] ));
    CFG3 #( .INIT(8'h02) )  un1_mem_0_5_17 (.A(\mem_12_[1]_net_1 ), .B(
        N_469), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_17_net_1));
    SLE \mem_15_[1]  (.D(CoreAPB3_0_APBmslave2_PWDATA[1]), .CLK(
        FCCC_0_GL1), .EN(mem_15__1_sqmuxa), .ALn(un1_mem_0_5_249_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_15_rs[1] ));
    CFG3 #( .INIT(8'hF8) )  un1_mem_0_5_88_set_RNICCUB (.A(
        un1_mem_0_5_88_set_net_1), .B(un1_mem_0_5_207_rs_net_1), .C(
        \mem_11_rs[0] ), .Y(\mem_11_[0]_net_1 ));
    CFG1 #( .INIT(2'h1) )  un1_mem_0_5_32_set_RNO (.A(
        un1_mem_0_5_32_net_1), .Y(un1_mem_0_5_32_i));
    CFG3 #( .INIT(8'hF2) )  un1_mem_0_5_176 (.A(\mem_5_[2]_net_1 ), .B(
        N_472), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_176_i));
    SLE un1_mem_0_5_66_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_8__1_sqmuxa), .ALn(un1_mem_0_5_66_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_mem_0_5_66_set_net_1));
    SLE un1_mem_0_5_204_rs (.D(VCC_net_1), .CLK(un1_mem_0_5_125_net_1), 
        .EN(VCC_net_1), .ALn(un1_mem_0_5_204_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(VCC_net_1), .Q(
        un1_mem_0_5_204_rs_net_1));
    CFG3 #( .INIT(8'hF2) )  un1_mem_0_5_204 (.A(\mem_7_[0]_net_1 ), .B(
        N_480), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_204_i));
    SLE un1_mem_0_5_11_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_4__1_sqmuxa), .ALn(un1_mem_0_5_11_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_mem_0_5_11_set_net_1));
    CFG3 #( .INIT(8'hF2) )  un1_mem_0_5_235 (.A(\mem_13_[3]_net_1 ), 
        .B(N_477), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_235_i));
    CFG3 #( .INIT(8'h02) )  un1_mem_0_5_108 (.A(\mem_13_[4]_net_1 ), 
        .B(N_477), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_108_net_1));
    CFG1 #( .INIT(2'h1) )  un1_mem_0_5_23_set_RNO (.A(
        un1_mem_0_5_23_net_1), .Y(un1_mem_0_5_23_i));
    CFG4 #( .INIT(16'h7350) )  \temp_data_2_15_i_3[3]  (.A(
        \mem_14_[3]_net_1 ), .B(\mem_2_[3]_net_1 ), .C(N_482), .D(
        N_478), .Y(\temp_data_2_15_i_3[3]_net_1 ));
    SLE \data_out[6]  (.D(\temp_data[6]_net_1 ), .CLK(FCCC_0_GL1), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(
        CoreAPB3_0_APBmslave3_PRDATA[6]));
    SLE \data_out[0]  (.D(\temp_data[0]_net_1 ), .CLK(FCCC_0_GL1), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(
        CoreAPB3_0_APBmslave3_PRDATA[0]));
    CFG3 #( .INIT(8'h02) )  un1_mem_0_5_120 (.A(\mem_2_[7]_net_1 ), .B(
        N_478), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_120_net_1));
    CFG3 #( .INIT(8'h02) )  un1_mem_0_5_111 (.A(\mem_13_[7]_net_1 ), 
        .B(N_477), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_111_net_1));
    CFG1 #( .INIT(2'h1) )  un1_mem_0_5_42_set_RNO (.A(
        un1_mem_0_5_42_net_1), .Y(un1_mem_0_5_42_i));
    SLE un1_mem_0_5_128_rs (.D(VCC_net_1), .CLK(un1_mem_0_5_81_net_1), 
        .EN(VCC_net_1), .ALn(un1_mem_0_5_128_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(VCC_net_1), .Q(
        un1_mem_0_5_128_rs_net_1));
    CFG1 #( .INIT(2'h1) )  un1_mem_0_5_7_set_RNO (.A(
        un1_mem_0_5_7_net_1), .Y(un1_mem_0_5_7_i));
    CFG3 #( .INIT(8'h02) )  un1_mem_0_5_36 (.A(\mem_2_[5]_net_1 ), .B(
        N_478), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_36_net_1));
    SLE un1_mem_0_5_71_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_8__1_sqmuxa), .ALn(un1_mem_0_5_71_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_mem_0_5_71_set_net_1));
    CFG3 #( .INIT(8'hF8) )  \mem_3__RNI5HO01[1]  (.A(
        un1_mem_0_5_124_set_net_1), .B(un1_mem_0_5_153_rs_net_1), .C(
        \mem_3_rs[1] ), .Y(\mem_3_[1]_net_1 ));
    CFG4 #( .INIT(16'h0800) )  \WRITE_GEN.mem_14__2_i_a2[5]  (.A(
        CoreAPB3_0_APBmslave2_PADDR[3]), .B(
        CoreAPB3_0_APBmslave2_PADDR[2]), .C(
        CoreAPB3_0_APBmslave2_PADDR[0]), .D(
        CoreAPB3_0_APBmslave2_PADDR[1]), .Y(N_482));
    SLE \mem_8_[1]  (.D(CoreAPB3_0_APBmslave2_PWDATA[1]), .CLK(
        FCCC_0_GL1), .EN(mem_8__1_sqmuxa), .ALn(un1_mem_0_5_221_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_8_rs[1] ));
    SLE un1_mem_0_5_233_rs (.D(VCC_net_1), .CLK(un1_mem_0_5_105_net_1), 
        .EN(VCC_net_1), .ALn(un1_mem_0_5_233_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(VCC_net_1), .Q(
        un1_mem_0_5_233_rs_net_1));
    SLE \mem_1_[7]  (.D(CoreAPB3_0_APBmslave2_PWDATA[7]), .CLK(
        FCCC_0_GL1), .EN(mem_1__1_sqmuxa), .ALn(un1_mem_0_5_143_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_1_rs[7] ));
    CFG3 #( .INIT(8'hF8) )  un1_mem_0_5_223_rs_RNIS0EV (.A(
        un1_mem_0_5_64_set_net_1), .B(un1_mem_0_5_223_rs_net_1), .C(
        \mem_8_rs[2] ), .Y(\mem_8_[2]_net_1 ));
    SLE \mem_9_[7]  (.D(CoreAPB3_0_APBmslave2_PWDATA[7]), .CLK(
        FCCC_0_GL1), .EN(mem_9__1_sqmuxa), .ALn(un1_mem_0_5_189_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_9_rs[7] ));
    SLE un1_mem_0_5_158_rs (.D(VCC_net_1), .CLK(un1_mem_0_5_53_net_1), 
        .EN(VCC_net_1), .ALn(un1_mem_0_5_158_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(VCC_net_1), .Q(
        un1_mem_0_5_158_rs_net_1));
    SLE \mem_1_[5]  (.D(CoreAPB3_0_APBmslave2_PWDATA[5]), .CLK(
        FCCC_0_GL1), .EN(mem_1__1_sqmuxa), .ALn(un1_mem_0_5_141_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_1_rs[5] ));
    CFG3 #( .INIT(8'h02) )  un1_mem_0_5_85 (.A(\mem_0_[4]_net_1 ), .B(
        N_473), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_85_net_1));
    CFG3 #( .INIT(8'h02) )  un1_mem_0_5 (.A(\mem_4_[0]_net_1 ), .B(
        N_476), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_net_1));
    SLE \temp_data[4]  (.D(N_16_i_0), .CLK(FCCC_0_GL1), .EN(rd_enable), 
        .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\temp_data[4]_net_1 ));
    CFG3 #( .INIT(8'h02) )  un1_mem_0_5_18 (.A(\mem_12_[2]_net_1 ), .B(
        N_469), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_18_net_1));
    SLE \mem_9_[5]  (.D(CoreAPB3_0_APBmslave2_PWDATA[5]), .CLK(
        FCCC_0_GL1), .EN(mem_9__1_sqmuxa), .ALn(un1_mem_0_5_185_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_9_rs[5] ));
    CFG1 #( .INIT(2'h1) )  un1_mem_0_5_6_set_RNO (.A(
        un1_mem_0_5_6_net_1), .Y(un1_mem_0_5_6_i));
    SLE un1_mem_0_5_81_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_0__1_sqmuxa), .ALn(un1_mem_0_5_81_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_mem_0_5_81_set_net_1));
    CFG3 #( .INIT(8'h02) )  un1_mem_0_5_19 (.A(\mem_12_[3]_net_1 ), .B(
        N_469), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_19_net_1));
    CFG3 #( .INIT(8'hF2) )  un1_mem_0_5_186 (.A(\mem_5_[7]_net_1 ), .B(
        N_472), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_186_i));
    SLE un1_mem_0_5_137_rs (.D(VCC_net_1), .CLK(un1_mem_0_5_12_net_1), 
        .EN(VCC_net_1), .ALn(un1_mem_0_5_137_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(VCC_net_1), .Q(
        un1_mem_0_5_137_rs_net_1));
    CFG4 #( .INIT(16'h0001) )  \temp_data_RNO[5]  (.A(
        \temp_data_2_15_i_4[5]_net_1 ), .B(
        \temp_data_2_15_i_5[5]_net_1 ), .C(
        \temp_data_2_15_i_11[5]_net_1 ), .D(
        \temp_data_2_15_i_12[5]_net_1 ), .Y(N_39_i_0));
    CFG3 #( .INIT(8'hF8) )  un1_mem_0_5_14_set_RNILPRT (.A(
        un1_mem_0_5_14_set_net_1), .B(un1_mem_0_5_138_rs_net_1), .C(
        \mem_1_rs[2] ), .Y(\mem_1_[2]_net_1 ));
    CFG1 #( .INIT(2'h1) )  un1_mem_0_5_91_set_RNO (.A(
        un1_mem_0_5_91_net_1), .Y(un1_mem_0_5_91_i));
    CFG3 #( .INIT(8'hF2) )  un1_mem_0_5_196 (.A(\mem_6_[4]_net_1 ), .B(
        N_468), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_196_i));
    CFG3 #( .INIT(8'hF2) )  un1_mem_0_5_205 (.A(\mem_10_[7]_net_1 ), 
        .B(N_471), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_205_i));
    CFG3 #( .INIT(8'hF8) )  un1_mem_0_5_159_rs_RNI4GOJ (.A(
        un1_mem_0_5_83_set_net_1), .B(un1_mem_0_5_159_rs_net_1), .C(
        \mem_3_rs[6] ), .Y(\mem_3_[6]_net_1 ));
    CFG1 #( .INIT(2'h1) )  un1_mem_0_5_115_set_RNO (.A(
        un1_mem_0_5_115_net_1), .Y(un1_mem_0_5_115_i));
    CFG3 #( .INIT(8'hF8) )  un1_mem_0_5_106_set_RNINRVV (.A(
        un1_mem_0_5_106_set_net_1), .B(un1_mem_0_5_234_rs_net_1), .C(
        \mem_13_rs[2] ), .Y(\mem_13_[2]_net_1 ));
    SLE \mem_12_[4]  (.D(CoreAPB3_0_APBmslave2_PWDATA[4]), .CLK(
        FCCC_0_GL1), .EN(mem_12__1_sqmuxa), .ALn(un1_mem_0_5_228_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_12_rs[4] ));
    SLE \mem_10_[3]  (.D(CoreAPB3_0_APBmslave2_PWDATA[3]), .CLK(
        FCCC_0_GL1), .EN(mem_10__1_sqmuxa), .ALn(un1_mem_0_5_197_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_10_rs[3] ));
    CFG3 #( .INIT(8'h02) )  un1_mem_0_5_84 (.A(\mem_0_[3]_net_1 ), .B(
        N_473), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_84_net_1));
    CFG3 #( .INIT(8'hF8) )  un1_mem_0_5_131_rs_RNIEHEP (.A(
        un1_mem_0_5_80_set_net_1), .B(un1_mem_0_5_131_rs_net_1), .C(
        \mem_0_rs[0] ), .Y(\mem_0_[0]_net_1 ));
    CFG1 #( .INIT(2'h1) )  un1_mem_0_5_110_set_RNO (.A(
        un1_mem_0_5_110_net_1), .Y(un1_mem_0_5_110_i));
    CFG1 #( .INIT(2'h1) )  un1_mem_0_5_118_set_RNO (.A(
        un1_mem_0_5_118_net_1), .Y(un1_mem_0_5_118_i));
    SLE un1_mem_0_5_248_rs (.D(VCC_net_1), .CLK(un1_mem_0_5_57_net_1), 
        .EN(VCC_net_1), .ALn(un1_mem_0_5_248_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(VCC_net_1), .Q(
        un1_mem_0_5_248_rs_net_1));
    SLE \mem_3_[3]  (.D(CoreAPB3_0_APBmslave2_PWDATA[3]), .CLK(
        FCCC_0_GL1), .EN(mem_3__1_sqmuxa), .ALn(un1_mem_0_5_155_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_3_rs[3] ));
    CFG3 #( .INIT(8'h02) )  un1_mem_0_5_77 (.A(\mem_9_[5]_net_1 ), .B(
        N_467), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_77_net_1));
    SLE un1_mem_0_5_40_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_5__1_sqmuxa), .ALn(un1_mem_0_5_40_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_mem_0_5_40_set_net_1));
    CFG3 #( .INIT(8'hF8) )  \mem_11__RNIHEPQ[6]  (.A(
        un1_mem_0_5_94_set_net_1), .B(un1_mem_0_5_218_rs_net_1), .C(
        \mem_11_rs[6] ), .Y(\mem_11_[6]_net_1 ));
    CFG2 #( .INIT(4'h8) )  mem_10__1_sqmuxa_0_a2 (.A(N_471), .B(
        wr_enable), .Y(mem_10__1_sqmuxa));
    SLE un1_mem_0_5_93_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_11__1_sqmuxa), .ALn(un1_mem_0_5_93_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_mem_0_5_93_set_net_1));
    SLE un1_mem_0_5_247_rs (.D(VCC_net_1), .CLK(un1_mem_0_5_119_net_1), 
        .EN(VCC_net_1), .ALn(un1_mem_0_5_247_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(VCC_net_1), .Q(
        un1_mem_0_5_247_rs_net_1));
    SLE un1_mem_0_5_23_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_12__1_sqmuxa), .ALn(un1_mem_0_5_23_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_mem_0_5_23_set_net_1));
    SLE \mem_13_[2]  (.D(CoreAPB3_0_APBmslave2_PWDATA[2]), .CLK(
        FCCC_0_GL1), .EN(mem_13__1_sqmuxa), .ALn(un1_mem_0_5_234_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_13_rs[2] ));
    SLE un1_mem_0_5_224_rs (.D(VCC_net_1), .CLK(un1_mem_0_5_17_net_1), 
        .EN(VCC_net_1), .ALn(un1_mem_0_5_224_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(VCC_net_1), .Q(
        un1_mem_0_5_224_rs_net_1));
    SLE un1_mem_0_5_206_rs (.D(VCC_net_1), .CLK(un1_mem_0_5_127_net_1), 
        .EN(VCC_net_1), .ALn(un1_mem_0_5_206_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(VCC_net_1), .Q(
        un1_mem_0_5_206_rs_net_1));
    CFG3 #( .INIT(8'hF2) )  un1_mem_0_5_252 (.A(\mem_15_[7]_net_1 ), 
        .B(N_474), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_252_i));
    CFG4 #( .INIT(16'h7530) )  \temp_data_2_15_i_7[0]  (.A(
        \mem_12_[0]_net_1 ), .B(\mem_8_[0]_net_1 ), .C(N_479), .D(
        N_469), .Y(\temp_data_2_15_i_7[0]_net_1 ));
    CFG1 #( .INIT(2'h1) )  un1_mem_0_5_24_set_RNO (.A(
        un1_mem_0_5_24_net_1), .Y(un1_mem_0_5_24_i));
    CFG3 #( .INIT(8'hF8) )  un1_mem_0_5_236_rs_RNITBIQ (.A(
        un1_mem_0_5_108_set_net_1), .B(un1_mem_0_5_236_rs_net_1), .C(
        \mem_13_rs[4] ), .Y(\mem_13_[4]_net_1 ));
    SLE \mem_12_[6]  (.D(CoreAPB3_0_APBmslave2_PWDATA[6]), .CLK(
        FCCC_0_GL1), .EN(mem_12__1_sqmuxa), .ALn(un1_mem_0_5_230_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_12_rs[6] ));
    SLE un1_mem_0_5_163_rs (.D(VCC_net_1), .CLK(un1_mem_0_5_4_net_1), 
        .EN(VCC_net_1), .ALn(un1_mem_0_5_163_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(VCC_net_1), .Q(
        un1_mem_0_5_163_rs_net_1));
    CFG3 #( .INIT(8'h02) )  un1_mem_0_5_4 (.A(\mem_4_[2]_net_1 ), .B(
        N_476), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_4_net_1));
    CFG3 #( .INIT(8'hF8) )  un1_mem_0_5_250_rs_RNIB6LI (.A(
        un1_mem_0_5_56_set_net_1), .B(un1_mem_0_5_250_rs_net_1), .C(
        \mem_15_rs[2] ), .Y(\mem_15_[2]_net_1 ));
    CFG3 #( .INIT(8'h02) )  un1_mem_0_5_83 (.A(\mem_3_[6]_net_1 ), .B(
        N_470), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_83_net_1));
    SLE un1_mem_0_5_115_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_14__1_sqmuxa), .ALn(un1_mem_0_5_115_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_mem_0_5_115_set_net_1));
    CFG1 #( .INIT(2'h1) )  un1_mem_0_5_105_set_RNO (.A(
        un1_mem_0_5_105_net_1), .Y(un1_mem_0_5_105_i));
    CFG3 #( .INIT(8'hF8) )  un1_mem_0_5_197_rs_RNIL735 (.A(
        un1_mem_0_5_96_set_net_1), .B(un1_mem_0_5_197_rs_net_1), .C(
        \mem_10_rs[3] ), .Y(\mem_10_[3]_net_1 ));
    CFG1 #( .INIT(2'h1) )  un1_mem_0_5_100_set_RNO (.A(
        un1_mem_0_5_100_net_1), .Y(un1_mem_0_5_100_i));
    SLE \mem_11_[2]  (.D(CoreAPB3_0_APBmslave2_PWDATA[2]), .CLK(
        FCCC_0_GL1), .EN(mem_11__1_sqmuxa), .ALn(un1_mem_0_5_211_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_11_rs[2] ));
    CFG1 #( .INIT(2'h1) )  un1_mem_0_5_108_set_RNO (.A(
        un1_mem_0_5_108_net_1), .Y(un1_mem_0_5_108_i));
    CFG3 #( .INIT(8'h02) )  un1_mem_0_5_125 (.A(\mem_7_[0]_net_1 ), .B(
        N_480), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_125_net_1));
    CFG3 #( .INIT(8'hF2) )  un1_mem_0_5_171 (.A(\mem_8_[6]_net_1 ), .B(
        N_479), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_171_i));
    SLE un1_mem_0_5_254_rs (.D(VCC_net_1), .CLK(un1_mem_0_5_62_net_1), 
        .EN(VCC_net_1), .ALn(un1_mem_0_5_254_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(VCC_net_1), .Q(
        un1_mem_0_5_254_rs_net_1));
    CFG1 #( .INIT(2'h1) )  un1_mem_0_5_123_set_RNO (.A(
        un1_mem_0_5_123_net_1), .Y(un1_mem_0_5_123_i));
    CFG3 #( .INIT(8'hF8) )  \mem_8__RNICUH51[0]  (.A(
        un1_mem_0_5_7_set_net_1), .B(un1_mem_0_5_219_rs_net_1), .C(
        \mem_8_rs[0] ), .Y(\mem_8_[0]_net_1 ));
    SLE un1_mem_0_5_14_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_1__1_sqmuxa), .ALn(un1_mem_0_5_14_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_mem_0_5_14_set_net_1));
    CFG3 #( .INIT(8'hF2) )  un1_mem_0_5_242 (.A(\mem_14_[2]_net_1 ), 
        .B(N_482), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_242_i));
    CFG3 #( .INIT(8'hF2) )  un1_mem_0_5_218 (.A(\mem_11_[6]_net_1 ), 
        .B(N_475), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_218_i));
    CFG4 #( .INIT(16'h7350) )  \temp_data_2_15_i_3[7]  (.A(
        \mem_14_[7]_net_1 ), .B(\mem_2_[7]_net_1 ), .C(N_482), .D(
        N_478), .Y(\temp_data_2_15_i_3[7]_net_1 ));
    SLE \mem_7_[2]  (.D(CoreAPB3_0_APBmslave2_PWDATA[2]), .CLK(
        FCCC_0_GL1), .EN(mem_7__1_sqmuxa), .ALn(un1_mem_0_5_208_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_7_rs[2] ));
    SLE un1_mem_0_5_97_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_10__1_sqmuxa), .ALn(un1_mem_0_5_97_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_mem_0_5_97_set_net_1));
    CFG1 #( .INIT(2'h1) )  un1_mem_0_5_81_set_RNO (.A(
        un1_mem_0_5_81_net_1), .Y(un1_mem_0_5_81_i));
    SLE un1_mem_0_5_198_rs (.D(VCC_net_1), .CLK(un1_mem_0_5_39_net_1), 
        .EN(VCC_net_1), .ALn(un1_mem_0_5_198_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(VCC_net_1), .Q(
        un1_mem_0_5_198_rs_net_1));
    SLE un1_mem_0_5_27_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_5__1_sqmuxa), .ALn(un1_mem_0_5_27_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_mem_0_5_27_set_net_1));
    CFG4 #( .INIT(16'h0002) )  \WRITE_GEN.mem_8__2_i_a2[7]  (.A(
        CoreAPB3_0_APBmslave2_PADDR[3]), .B(
        CoreAPB3_0_APBmslave2_PADDR[2]), .C(
        CoreAPB3_0_APBmslave2_PADDR[0]), .D(
        CoreAPB3_0_APBmslave2_PADDR[1]), .Y(N_479));
    SLE un1_mem_0_5_103_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_10__1_sqmuxa), .ALn(un1_mem_0_5_103_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_mem_0_5_103_set_net_1));
    SLE \mem_2_[2]  (.D(CoreAPB3_0_APBmslave2_PWDATA[2]), .CLK(
        FCCC_0_GL1), .EN(mem_2__1_sqmuxa), .ALn(un1_mem_0_5_146_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_2_rs[2] ));
    CFG1 #( .INIT(2'h1) )  un1_mem_0_5_66_set_RNO (.A(
        un1_mem_0_5_66_net_1), .Y(un1_mem_0_5_66_i));
    CFG3 #( .INIT(8'hF8) )  un1_mem_0_5_21_set_RNI99FV (.A(
        un1_mem_0_5_21_set_net_1), .B(un1_mem_0_5_229_rs_net_1), .C(
        \mem_12_rs[5] ), .Y(\mem_12_[5]_net_1 ));
    CFG3 #( .INIT(8'h02) )  un1_mem_0_5_15 (.A(\mem_5_[1]_net_1 ), .B(
        N_472), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_15_net_1));
    SLE un1_mem_0_5_74_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_9__1_sqmuxa), .ALn(un1_mem_0_5_74_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_mem_0_5_74_set_net_1));
    CFG3 #( .INIT(8'hF8) )  un1_mem_0_5_242_rs_RNIMQ38 (.A(
        un1_mem_0_5_114_set_net_1), .B(un1_mem_0_5_242_rs_net_1), .C(
        \mem_14_rs[2] ), .Y(\mem_14_[2]_net_1 ));
    SLE un1_mem_0_5_173_rs (.D(VCC_net_1), .CLK(un1_mem_0_5_71_net_1), 
        .EN(VCC_net_1), .ALn(un1_mem_0_5_173_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(VCC_net_1), .Q(
        un1_mem_0_5_173_rs_net_1));
    CFG3 #( .INIT(8'h02) )  un1_mem_0_5_78 (.A(\mem_9_[6]_net_1 ), .B(
        N_467), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_78_net_1));
    CFG3 #( .INIT(8'hF2) )  un1_mem_0_5_156 (.A(\mem_3_[4]_net_1 ), .B(
        N_470), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_156_i));
    SLE \mem_5_[7]  (.D(CoreAPB3_0_APBmslave2_PWDATA[7]), .CLK(
        FCCC_0_GL1), .EN(mem_5__1_sqmuxa), .ALn(un1_mem_0_5_186_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_5_rs[7] ));
    CFG1 #( .INIT(2'h1) )  un1_mem_0_5_68_set_RNO (.A(
        un1_mem_0_5_68_net_1), .Y(un1_mem_0_5_68_i));
    SLE \mem_4_[2]  (.D(CoreAPB3_0_APBmslave2_PWDATA[2]), .CLK(
        FCCC_0_GL1), .EN(mem_4__1_sqmuxa), .ALn(un1_mem_0_5_163_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_4_rs[2] ));
    CFG3 #( .INIT(8'hF8) )  \mem_2__RNIVPBK[5]  (.A(
        un1_mem_0_5_36_set_net_1), .B(un1_mem_0_5_149_rs_net_1), .C(
        \mem_2_rs[5] ), .Y(\mem_2_[5]_net_1 ));
    SLE un1_mem_0_5_1_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_7__1_sqmuxa), .ALn(un1_mem_0_5_1_i), .ADn(GND_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_mem_0_5_1_set_net_1));
    SLE un1_mem_0_5_96_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_10__1_sqmuxa), .ALn(un1_mem_0_5_96_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_mem_0_5_96_set_net_1));
    CFG3 #( .INIT(8'h02) )  un1_mem_0_5_79 (.A(\mem_9_[7]_net_1 ), .B(
        N_467), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_79_net_1));
    SLE \mem_8_[6]  (.D(CoreAPB3_0_APBmslave2_PWDATA[6]), .CLK(
        FCCC_0_GL1), .EN(mem_8__1_sqmuxa), .ALn(un1_mem_0_5_171_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_8_rs[6] ));
    CFG3 #( .INIT(8'hF2) )  un1_mem_0_5_219 (.A(\mem_8_[0]_net_1 ), .B(
        N_479), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_219_i));
    SLE un1_mem_0_5_26_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_2__1_sqmuxa), .ALn(un1_mem_0_5_26_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_mem_0_5_26_set_net_1));
    SLE un1_mem_0_5_202_rs (.D(VCC_net_1), .CLK(un1_mem_0_5_123_net_1), 
        .EN(VCC_net_1), .ALn(un1_mem_0_5_202_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(VCC_net_1), .Q(
        un1_mem_0_5_202_rs_net_1));
    CFG3 #( .INIT(8'hF2) )  un1_mem_0_5_221 (.A(\mem_8_[1]_net_1 ), .B(
        N_479), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_221_i));
    CFG3 #( .INIT(8'hF2) )  un1_mem_0_5_232 (.A(\mem_13_[0]_net_1 ), 
        .B(N_477), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_232_i));
    SLE \mem_5_[5]  (.D(CoreAPB3_0_APBmslave2_PWDATA[5]), .CLK(
        FCCC_0_GL1), .EN(mem_5__1_sqmuxa), .ALn(un1_mem_0_5_182_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_5_rs[5] ));
    CFG4 #( .INIT(16'h7350) )  \temp_data_2_15_i_4[4]  (.A(
        \mem_10_[4]_net_1 ), .B(\mem_6_[4]_net_1 ), .C(N_471), .D(
        N_468), .Y(\temp_data_2_15_i_4[4]_net_1 ));
    CFG3 #( .INIT(8'h02) )  un1_mem_0_5_14 (.A(\mem_1_[2]_net_1 ), .B(
        N_481), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_14_net_1));
    CFG4 #( .INIT(16'h7350) )  \temp_data_2_15_i_4[7]  (.A(
        \mem_10_[7]_net_1 ), .B(\mem_6_[7]_net_1 ), .C(N_471), .D(
        N_468), .Y(\temp_data_2_15_i_4[7]_net_1 ));
    CFG3 #( .INIT(8'h02) )  un1_mem_0_5_80 (.A(\mem_0_[0]_net_1 ), .B(
        N_473), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_80_net_1));
    SLE un1_mem_0_5_180_rs (.D(VCC_net_1), .CLK(un1_mem_0_5_44_net_1), 
        .EN(VCC_net_1), .ALn(un1_mem_0_5_180_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(VCC_net_1), .Q(
        un1_mem_0_5_180_rs_net_1));
    SLE un1_mem_0_5_238_rs (.D(VCC_net_1), .CLK(un1_mem_0_5_110_net_1), 
        .EN(VCC_net_1), .ALn(un1_mem_0_5_238_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(VCC_net_1), .Q(
        un1_mem_0_5_238_rs_net_1));
    CFG3 #( .INIT(8'hF2) )  un1_mem_0_5_146 (.A(\mem_2_[2]_net_1 ), .B(
        N_478), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_146_i));
    CFG3 #( .INIT(8'h02) )  un1_mem_0_5_112 (.A(\mem_14_[0]_net_1 ), 
        .B(N_482), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_112_net_1));
    SLE un1_mem_0_5_84_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_0__1_sqmuxa), .ALn(un1_mem_0_5_84_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_mem_0_5_84_set_net_1));
    SLE un1_mem_0_5_237_rs (.D(VCC_net_1), .CLK(un1_mem_0_5_109_net_1), 
        .EN(VCC_net_1), .ALn(un1_mem_0_5_237_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(VCC_net_1), .Q(
        un1_mem_0_5_237_rs_net_1));
    CFG3 #( .INIT(8'hF2) )  un1_mem_0_5_227 (.A(\mem_12_[3]_net_1 ), 
        .B(N_469), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_227_i));
    CFG2 #( .INIT(4'h8) )  mem_13__1_sqmuxa_0_a2 (.A(N_477), .B(
        wr_enable), .Y(mem_13__1_sqmuxa));
    CFG3 #( .INIT(8'hF2) )  un1_mem_0_5_181 (.A(\mem_9_[3]_net_1 ), .B(
        N_467), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_181_i));
    SLE un1_mem_0_5_145_rs (.D(VCC_net_1), .CLK(un1_mem_0_5_28_net_1), 
        .EN(VCC_net_1), .ALn(un1_mem_0_5_145_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(VCC_net_1), .Q(
        un1_mem_0_5_145_rs_net_1));
    CFG3 #( .INIT(8'h02) )  un1_mem_0_5_62 (.A(\mem_15_[5]_net_1 ), .B(
        N_474), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_62_net_1));
    CFG3 #( .INIT(8'hF8) )  un1_mem_0_5_84_set_RNIK14P (.A(
        un1_mem_0_5_84_set_net_1), .B(un1_mem_0_5_130_rs_net_1), .C(
        \mem_0_rs[3] ), .Y(\mem_0_[3]_net_1 ));
    SLE un1_mem_0_5_42_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_5__1_sqmuxa), .ALn(un1_mem_0_5_42_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_mem_0_5_42_set_net_1));
    SLE un1_mem_0_5_226_rs (.D(VCC_net_1), .CLK(un1_mem_0_5_18_net_1), 
        .EN(VCC_net_1), .ALn(un1_mem_0_5_226_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(VCC_net_1), .Q(
        un1_mem_0_5_226_rs_net_1));
    CFG3 #( .INIT(8'hF2) )  un1_mem_0_5_191 (.A(\mem_10_[0]_net_1 ), 
        .B(N_471), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_191_i));
    CFG3 #( .INIT(8'hF8) )  un1_mem_0_5_73_set_RNI40PO (.A(
        un1_mem_0_5_73_set_net_1), .B(un1_mem_0_5_177_rs_net_1), .C(
        \mem_9_rs[1] ), .Y(\mem_9_[1]_net_1 ));
    CFG3 #( .INIT(8'hF8) )  un1_mem_0_5_251_rs_RNI9R3P (.A(
        un1_mem_0_5_61_set_net_1), .B(un1_mem_0_5_251_rs_net_1), .C(
        \mem_15_rs[3] ), .Y(\mem_15_[3]_net_1 ));
    CFG3 #( .INIT(8'hF2) )  un1_mem_0_5_160 (.A(\mem_3_[7]_net_1 ), .B(
        N_470), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_160_i));
    SLE un1_mem_0_5_141_rs (.D(VCC_net_1), .CLK(un1_mem_0_5_47_net_1), 
        .EN(VCC_net_1), .ALn(un1_mem_0_5_141_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(VCC_net_1), .Q(
        un1_mem_0_5_141_rs_net_1));
    CFG3 #( .INIT(8'hF8) )  \mem_15__RNIHSDR[0]  (.A(
        un1_mem_0_5_57_set_net_1), .B(un1_mem_0_5_248_rs_net_1), .C(
        \mem_15_rs[0] ), .Y(\mem_15_[0]_net_1 ));
    SLE un1_mem_0_5_125_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_7__1_sqmuxa), .ALn(un1_mem_0_5_125_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_mem_0_5_125_set_net_1));
    CFG3 #( .INIT(8'hF8) )  un1_mem_0_5_107_set_RNIQ3951 (.A(
        un1_mem_0_5_107_set_net_1), .B(un1_mem_0_5_235_rs_net_1), .C(
        \mem_13_rs[3] ), .Y(\mem_13_[3]_net_1 ));
    CFG3 #( .INIT(8'h02) )  un1_mem_0_5_13 (.A(\mem_5_[0]_net_1 ), .B(
        N_472), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_13_net_1));
    CFG4 #( .INIT(16'h0004) )  \WRITE_GEN.mem_4__2_i_a2[5]  (.A(
        CoreAPB3_0_APBmslave2_PADDR[3]), .B(
        CoreAPB3_0_APBmslave2_PADDR[2]), .C(
        CoreAPB3_0_APBmslave2_PADDR[0]), .D(
        CoreAPB3_0_APBmslave2_PADDR[1]), .Y(N_476));
    CFG1 #( .INIT(2'h1) )  un1_mem_0_5_62_set_RNO (.A(
        un1_mem_0_5_62_net_1), .Y(un1_mem_0_5_62_i));
    CFG4 #( .INIT(16'h7530) )  \temp_data_2_15_i_0[0]  (.A(
        \mem_9_[0]_net_1 ), .B(\mem_1_[0]_net_1 ), .C(N_481), .D(N_467)
        , .Y(\temp_data_2_15_i_0[0]_net_1 ));
    SLE un1_mem_0_5_45_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_1__1_sqmuxa), .ALn(un1_mem_0_5_45_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_mem_0_5_45_set_net_1));
    CFG3 #( .INIT(8'hF2) )  un1_mem_0_5_213 (.A(\mem_7_[5]_net_1 ), .B(
        N_480), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_213_i));
    CFG3 #( .INIT(8'hF2) )  un1_mem_0_5_136 (.A(\mem_1_[0]_net_1 ), .B(
        N_481), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_136_i));
    SLE \mem_7_[1]  (.D(CoreAPB3_0_APBmslave2_PWDATA[1]), .CLK(
        FCCC_0_GL1), .EN(mem_7__1_sqmuxa), .ALn(un1_mem_0_5_206_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_7_rs[1] ));
    SLE \mem_10_[0]  (.D(CoreAPB3_0_APBmslave2_PWDATA[0]), .CLK(
        FCCC_0_GL1), .EN(mem_10__1_sqmuxa), .ALn(un1_mem_0_5_191_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_10_rs[0] ));
    SLE \mem_13_[7]  (.D(CoreAPB3_0_APBmslave2_PWDATA[7]), .CLK(
        FCCC_0_GL1), .EN(mem_13__1_sqmuxa), .ALn(un1_mem_0_5_239_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_13_rs[7] ));
    SLE \mem_14_[5]  (.D(CoreAPB3_0_APBmslave2_PWDATA[5]), .CLK(
        FCCC_0_GL1), .EN(mem_14__1_sqmuxa), .ALn(un1_mem_0_5_245_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_14_rs[5] ));
    CFG4 #( .INIT(16'h0001) )  \temp_data_RNO[3]  (.A(
        \temp_data_2_15_i_4[3]_net_1 ), .B(
        \temp_data_2_15_i_5[3]_net_1 ), .C(
        \temp_data_2_15_i_11[3]_net_1 ), .D(
        \temp_data_2_15_i_12[3]_net_1 ), .Y(N_12_i_0));
    CFG3 #( .INIT(8'hF2) )  un1_mem_0_5_202 (.A(\mem_6_[7]_net_1 ), .B(
        N_468), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_202_i));
    CFG3 #( .INIT(8'h02) )  un1_mem_0_5_123 (.A(\mem_6_[7]_net_1 ), .B(
        N_468), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_123_net_1));
    CFG1 #( .INIT(2'h1) )  un1_mem_0_5_11_set_RNO (.A(
        un1_mem_0_5_11_net_1), .Y(un1_mem_0_5_11_i));
    CFG4 #( .INIT(16'h7530) )  \temp_data_2_15_i_0[2]  (.A(
        \mem_9_[2]_net_1 ), .B(\mem_1_[2]_net_1 ), .C(N_481), .D(N_467)
        , .Y(\temp_data_2_15_i_0[2]_net_1 ));
    SLE \mem_2_[1]  (.D(CoreAPB3_0_APBmslave2_PWDATA[1]), .CLK(
        FCCC_0_GL1), .EN(mem_2__1_sqmuxa), .ALn(un1_mem_0_5_145_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_2_rs[1] ));
    CFG3 #( .INIT(8'h02) )  un1_mem_0_5_91 (.A(\mem_11_[3]_net_1 ), .B(
        N_475), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_91_net_1));
    CFG3 #( .INIT(8'hF8) )  \mem_7__RNIA31M[7]  (.A(
        un1_mem_0_5_1_set_net_1), .B(un1_mem_0_5_217_rs_net_1), .C(
        \mem_7_rs[7] ), .Y(\mem_7_[7]_net_1 ));
    CFG2 #( .INIT(4'h8) )  mem_0__1_sqmuxa_0_a2 (.A(N_473), .B(
        wr_enable), .Y(mem_0__1_sqmuxa));
    SLE \mem_3_[4]  (.D(CoreAPB3_0_APBmslave2_PWDATA[4]), .CLK(
        FCCC_0_GL1), .EN(mem_3__1_sqmuxa), .ALn(un1_mem_0_5_156_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_3_rs[4] ));
    CFG3 #( .INIT(8'hF2) )  un1_mem_0_5_250 (.A(\mem_15_[2]_net_1 ), 
        .B(N_474), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_250_i));
    CFG4 #( .INIT(16'hFFFE) )  \temp_data_2_15_i_12[1]  (.A(
        \temp_data_2_15_i_3[1]_net_1 ), .B(
        \temp_data_2_15_i_2[1]_net_1 ), .C(
        \temp_data_2_15_i_1[1]_net_1 ), .D(
        \temp_data_2_15_i_0[1]_net_1 ), .Y(
        \temp_data_2_15_i_12[1]_net_1 ));
    SLE \mem_4_[1]  (.D(CoreAPB3_0_APBmslave2_PWDATA[1]), .CLK(
        FCCC_0_GL1), .EN(mem_4__1_sqmuxa), .ALn(un1_mem_0_5_162_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_4_rs[1] ));
    CFG3 #( .INIT(8'h02) )  un1_mem_0_5_75 (.A(\mem_9_[3]_net_1 ), .B(
        N_467), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_75_net_1));
    SLE \mem_11_[7]  (.D(CoreAPB3_0_APBmslave2_PWDATA[7]), .CLK(
        FCCC_0_GL1), .EN(mem_11__1_sqmuxa), .ALn(un1_mem_0_5_220_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_11_rs[7] ));
    CFG4 #( .INIT(16'h7350) )  \temp_data_2_15_i_4[1]  (.A(
        \mem_10_[1]_net_1 ), .B(\mem_6_[1]_net_1 ), .C(N_471), .D(
        N_468), .Y(\temp_data_2_15_i_4[1]_net_1 ));
    SLE \mem_14_[1]  (.D(CoreAPB3_0_APBmslave2_PWDATA[1]), .CLK(
        FCCC_0_GL1), .EN(mem_14__1_sqmuxa), .ALn(un1_mem_0_5_241_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_14_rs[1] ));
    SLE un1_mem_0_5_31_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_6__1_sqmuxa), .ALn(un1_mem_0_5_31_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_mem_0_5_31_set_net_1));
    CFG1 #( .INIT(2'h1) )  un1_mem_0_5_93_set_RNO (.A(
        un1_mem_0_5_93_net_1), .Y(un1_mem_0_5_93_i));
    CFG1 #( .INIT(2'h1) )  un1_mem_0_5_57_set_RNO (.A(
        un1_mem_0_5_57_net_1), .Y(un1_mem_0_5_57_i));
    SLE un1_mem_0_5_142_rs (.D(VCC_net_1), .CLK(un1_mem_0_5_45_net_1), 
        .EN(VCC_net_1), .ALn(un1_mem_0_5_142_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(VCC_net_1), .Q(
        un1_mem_0_5_142_rs_net_1));
    SLE un1_mem_0_5_222_rs (.D(VCC_net_1), .CLK(un1_mem_0_5_16_net_1), 
        .EN(VCC_net_1), .ALn(un1_mem_0_5_222_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(VCC_net_1), .Q(
        un1_mem_0_5_222_rs_net_1));
    SLE un1_mem_0_5_149_rs (.D(VCC_net_1), .CLK(un1_mem_0_5_36_net_1), 
        .EN(VCC_net_1), .ALn(un1_mem_0_5_149_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(VCC_net_1), .Q(
        un1_mem_0_5_149_rs_net_1));
    CFG3 #( .INIT(8'hF8) )  \mem_6__RNI3UQI[6]  (.A(
        un1_mem_0_5_121_set_net_1), .B(un1_mem_0_5_200_rs_net_1), .C(
        \mem_6_rs[6] ), .Y(\mem_6_[6]_net_1 ));
    CFG3 #( .INIT(8'h02) )  un1_mem_0_5_31 (.A(\mem_6_[1]_net_1 ), .B(
        N_468), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_31_net_1));
    CFG1 #( .INIT(2'h1) )  un1_mem_0_5_55_set_RNO (.A(
        un1_mem_0_5_55_net_1), .Y(un1_mem_0_5_55_i));
    CFG4 #( .INIT(16'h7530) )  \temp_data_2_15_i_0[4]  (.A(
        \mem_9_[4]_net_1 ), .B(\mem_1_[4]_net_1 ), .C(N_481), .D(N_467)
        , .Y(\temp_data_2_15_i_0[4]_net_1 ));
    SLE un1_mem_0_5_7_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_8__1_sqmuxa), .ALn(un1_mem_0_5_7_i), .ADn(GND_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_mem_0_5_7_set_net_1));
    CFG3 #( .INIT(8'hF2) )  un1_mem_0_5_240 (.A(\mem_14_[0]_net_1 ), 
        .B(N_482), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_240_i));
    CFG3 #( .INIT(8'hF2) )  un1_mem_0_5_129 (.A(\mem_0_[2]_net_1 ), .B(
        N_473), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_129_i));
    CFG4 #( .INIT(16'h0040) )  \WRITE_GEN.mem_5__2_i_a2[5]  (.A(
        CoreAPB3_0_APBmslave2_PADDR[3]), .B(
        CoreAPB3_0_APBmslave2_PADDR[2]), .C(
        CoreAPB3_0_APBmslave2_PADDR[0]), .D(
        CoreAPB3_0_APBmslave2_PADDR[1]), .Y(N_472));
    CFG3 #( .INIT(8'h02) )  un1_mem_0_5_2 (.A(\mem_4_[1]_net_1 ), .B(
        N_476), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_2_net_1));
    CFG3 #( .INIT(8'h02) )  un1_mem_0_5_127 (.A(\mem_7_[1]_net_1 ), .B(
        N_480), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_127_net_1));
    CFG3 #( .INIT(8'h02) )  un1_mem_0_5_10 (.A(\mem_1_[0]_net_1 ), .B(
        N_481), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_10_net_1));
    CFG3 #( .INIT(8'hF8) )  \mem_4__RNI1LP21[1]  (.A(
        un1_mem_0_5_2_set_net_1), .B(un1_mem_0_5_162_rs_net_1), .C(
        \mem_4_rs[1] ), .Y(\mem_4_[1]_net_1 ));
    CFG4 #( .INIT(16'h0400) )  \WRITE_GEN.mem_6__2_i_a2[5]  (.A(
        CoreAPB3_0_APBmslave2_PADDR[3]), .B(
        CoreAPB3_0_APBmslave2_PADDR[2]), .C(
        CoreAPB3_0_APBmslave2_PADDR[0]), .D(
        CoreAPB3_0_APBmslave2_PADDR[1]), .Y(N_468));
    CFG3 #( .INIT(8'h02) )  un1_mem_0_5_74 (.A(\mem_9_[2]_net_1 ), .B(
        N_467), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_74_net_1));
    SLE \mem_6_[3]  (.D(CoreAPB3_0_APBmslave2_PWDATA[3]), .CLK(
        FCCC_0_GL1), .EN(mem_6__1_sqmuxa), .ALn(un1_mem_0_5_194_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_6_rs[3] ));
    CFG3 #( .INIT(8'hF8) )  un1_mem_0_5_31_set_RNIMA8B (.A(
        un1_mem_0_5_31_set_net_1), .B(un1_mem_0_5_190_rs_net_1), .C(
        \mem_6_rs[1] ), .Y(\mem_6_[1]_net_1 ));
    CFG3 #( .INIT(8'hF8) )  un1_mem_0_5_158_rs_RNI2CFK (.A(
        un1_mem_0_5_53_set_net_1), .B(un1_mem_0_5_158_rs_net_1), .C(
        \mem_7_rs[4] ), .Y(\mem_7_[4]_net_1 ));
    CFG3 #( .INIT(8'h02) )  un1_mem_0_5_106 (.A(\mem_13_[2]_net_1 ), 
        .B(N_477), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_106_net_1));
    CFG3 #( .INIT(8'hF2) )  un1_mem_0_5_151 (.A(\mem_2_[7]_net_1 ), .B(
        N_478), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_151_i));
    SLE un1_mem_0_5_118_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_14__1_sqmuxa), .ALn(un1_mem_0_5_118_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_mem_0_5_118_set_net_1));
    SLE un1_mem_0_5_135_rs (.D(VCC_net_1), .CLK(un1_mem_0_5_8_net_1), 
        .EN(VCC_net_1), .ALn(un1_mem_0_5_135_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(VCC_net_1), .Q(
        un1_mem_0_5_135_rs_net_1));
    CFG3 #( .INIT(8'hF2) )  un1_mem_0_5_172 (.A(\mem_5_[0]_net_1 ), .B(
        N_472), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_172_i));
    SLE un1_mem_0_5_252_rs (.D(VCC_net_1), .CLK(un1_mem_0_5_60_net_1), 
        .EN(VCC_net_1), .ALn(un1_mem_0_5_252_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(VCC_net_1), .Q(
        un1_mem_0_5_252_rs_net_1));
    SLE un1_mem_0_5_131_rs (.D(VCC_net_1), .CLK(un1_mem_0_5_80_net_1), 
        .EN(VCC_net_1), .ALn(un1_mem_0_5_131_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(VCC_net_1), .Q(
        un1_mem_0_5_131_rs_net_1));
    SLE \mem_3_[0]  (.D(CoreAPB3_0_APBmslave2_PWDATA[0]), .CLK(
        FCCC_0_GL1), .EN(mem_3__1_sqmuxa), .ALn(un1_mem_0_5_152_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_3_rs[0] ));
    SLE \mem_0_[3]  (.D(CoreAPB3_0_APBmslave2_PWDATA[3]), .CLK(
        FCCC_0_GL1), .EN(mem_0__1_sqmuxa), .ALn(un1_mem_0_5_130_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_0_rs[3] ));
    CFG3 #( .INIT(8'h02) )  un1_mem_0_5_5 (.A(\mem_8_[1]_net_1 ), .B(
        N_479), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_5_net_1));
    CFG3 #( .INIT(8'hF2) )  un1_mem_0_5_230 (.A(\mem_12_[6]_net_1 ), 
        .B(N_469), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_230_i));
    SLE un1_mem_0_5_150_rs (.D(VCC_net_1), .CLK(un1_mem_0_5_38_net_1), 
        .EN(VCC_net_1), .ALn(un1_mem_0_5_150_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(VCC_net_1), .Q(
        un1_mem_0_5_150_rs_net_1));
    CFG3 #( .INIT(8'hF8) )  \mem_12__RNI6V831[7]  (.A(
        un1_mem_0_5_23_set_net_1), .B(un1_mem_0_5_231_rs_net_1), .C(
        \mem_12_rs[7] ), .Y(\mem_12_[7]_net_1 ));
    CFG3 #( .INIT(8'hF2) )  un1_mem_0_5_141 (.A(\mem_1_[5]_net_1 ), .B(
        N_481), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_141_i));
    CFG4 #( .INIT(16'h7350) )  \temp_data_2_15_i_2[5]  (.A(
        \mem_13_[5]_net_1 ), .B(\mem_15_[5]_net_1 ), .C(N_477), .D(
        N_474), .Y(\temp_data_2_15_i_2[5]_net_1 ));
    CFG3 #( .INIT(8'hF2) )  un1_mem_0_5_165 (.A(\mem_4_[4]_net_1 ), .B(
        N_476), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_165_i));
    CFG3 #( .INIT(8'h02) )  un1_mem_0_5_73 (.A(\mem_9_[1]_net_1 ), .B(
        N_467), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_73_net_1));
    CFG4 #( .INIT(16'h7350) )  \temp_data_2_15_i_2[7]  (.A(
        \mem_13_[7]_net_1 ), .B(\mem_15_[7]_net_1 ), .C(N_477), .D(
        N_474), .Y(\temp_data_2_15_i_2[7]_net_1 ));
    CFG1 #( .INIT(2'h1) )  un1_mem_0_5_83_set_RNO (.A(
        un1_mem_0_5_83_net_1), .Y(un1_mem_0_5_83_i));
    SLE un1_mem_0_5_49_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_7__1_sqmuxa), .ALn(un1_mem_0_5_49_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_mem_0_5_49_set_net_1));
    SLE \mem_15_[4]  (.D(CoreAPB3_0_APBmslave2_PWDATA[4]), .CLK(
        FCCC_0_GL1), .EN(mem_15__1_sqmuxa), .ALn(un1_mem_0_5_253_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_15_rs[4] ));
    CFG3 #( .INIT(8'hF2) )  un1_mem_0_5_226 (.A(\mem_12_[2]_net_1 ), 
        .B(N_469), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_226_i));
    SLE un1_mem_0_5_241_rs (.D(VCC_net_1), .CLK(un1_mem_0_5_113_net_1), 
        .EN(VCC_net_1), .ALn(un1_mem_0_5_241_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(VCC_net_1), .Q(
        un1_mem_0_5_241_rs_net_1));
    CFG3 #( .INIT(8'hF8) )  un1_mem_0_5_173_rs_RNI3EQN (.A(
        un1_mem_0_5_71_set_net_1), .B(un1_mem_0_5_173_rs_net_1), .C(
        \mem_8_rs[7] ), .Y(\mem_8_[7]_net_1 ));
    SLE un1_mem_0_5_18_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_12__1_sqmuxa), .ALn(un1_mem_0_5_18_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_mem_0_5_18_set_net_1));
    CFG3 #( .INIT(8'hF8) )  \mem_3__RNI159N[0]  (.A(
        un1_mem_0_5_122_set_net_1), .B(un1_mem_0_5_152_rs_net_1), .C(
        \mem_3_rs[0] ), .Y(\mem_3_[0]_net_1 ));
    CFG1 #( .INIT(2'h1) )  un1_mem_0_5_59_set_RNO (.A(
        un1_mem_0_5_59_net_1), .Y(un1_mem_0_5_59_i));
    CFG3 #( .INIT(8'hF8) )  un1_mem_0_5_167_rs_RNI9A1R (.A(
        un1_mem_0_5_68_set_net_1), .B(un1_mem_0_5_167_rs_net_1), .C(
        \mem_8_rs[4] ), .Y(\mem_8_[4]_net_1 ));
    CFG3 #( .INIT(8'hF8) )  un1_mem_0_5_134_rs_RNIUS2Q (.A(
        un1_mem_0_5_87_set_net_1), .B(un1_mem_0_5_134_rs_net_1), .C(
        \mem_0_rs[6] ), .Y(\mem_0_[6]_net_1 ));
    CFG1 #( .INIT(2'h1) )  un1_mem_0_5_127_set_RNO (.A(
        un1_mem_0_5_127_net_1), .Y(un1_mem_0_5_127_i));
    SLE \mem_12_[3]  (.D(CoreAPB3_0_APBmslave2_PWDATA[3]), .CLK(
        FCCC_0_GL1), .EN(mem_12__1_sqmuxa), .ALn(un1_mem_0_5_227_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_12_rs[3] ));
    CFG1 #( .INIT(2'h1) )  un1_mem_0_5_71_set_RNO (.A(
        un1_mem_0_5_71_net_1), .Y(un1_mem_0_5_71_i));
    SLE un1_mem_0_5_245_rs (.D(VCC_net_1), .CLK(un1_mem_0_5_117_net_1), 
        .EN(VCC_net_1), .ALn(un1_mem_0_5_245_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(VCC_net_1), .Q(
        un1_mem_0_5_245_rs_net_1));
    CFG3 #( .INIT(8'h02) )  un1_mem_0_5_97 (.A(\mem_10_[0]_net_1 ), .B(
        N_471), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_97_net_1));
    CFG2 #( .INIT(4'h2) )  \temp_data_2_15_i_a2_13[1]  (.A(N_476), .B(
        \mem_4_[1]_net_1 ), .Y(N_345));
    SLE un1_mem_0_5_78_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_9__1_sqmuxa), .ALn(un1_mem_0_5_78_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_mem_0_5_78_set_net_1));
    CFG1 #( .INIT(2'h1) )  un1_mem_0_5_124_set_RNO (.A(
        un1_mem_0_5_124_net_1), .Y(un1_mem_0_5_124_i));
    CFG3 #( .INIT(8'hF8) )  \mem_7__RNI947S[6]  (.A(
        un1_mem_0_5_3_set_net_1), .B(un1_mem_0_5_215_rs_net_1), .C(
        \mem_7_rs[6] ), .Y(\mem_7_[6]_net_1 ));
    SLE \mem_7_[6]  (.D(CoreAPB3_0_APBmslave2_PWDATA[6]), .CLK(
        FCCC_0_GL1), .EN(mem_7__1_sqmuxa), .ALn(un1_mem_0_5_215_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_7_rs[6] ));
    CFG3 #( .INIT(8'hF2) )  un1_mem_0_5_131 (.A(\mem_0_[0]_net_1 ), .B(
        N_473), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_131_i));
    CFG3 #( .INIT(8'hF8) )  un1_mem_0_5_212_rs_RNI5DKN (.A(
        un1_mem_0_5_91_set_net_1), .B(un1_mem_0_5_212_rs_net_1), .C(
        \mem_11_rs[3] ), .Y(\mem_11_[3]_net_1 ));
    CFG3 #( .INIT(8'hF2) )  un1_mem_0_5_182 (.A(\mem_5_[5]_net_1 ), .B(
        N_472), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_182_i));
    SLE un1_mem_0_5_144_rs (.D(VCC_net_1), .CLK(un1_mem_0_5_26_net_1), 
        .EN(VCC_net_1), .ALn(un1_mem_0_5_144_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(VCC_net_1), .Q(
        un1_mem_0_5_144_rs_net_1));
    SLE \mem_15_[6]  (.D(CoreAPB3_0_APBmslave2_PWDATA[6]), .CLK(
        FCCC_0_GL1), .EN(mem_15__1_sqmuxa), .ALn(un1_mem_0_5_255_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_15_rs[6] ));
    CFG1 #( .INIT(2'h1) )  un1_mem_0_5_94_set_RNO (.A(
        un1_mem_0_5_94_net_1), .Y(un1_mem_0_5_94_i));
    SLE un1_mem_0_5_132_rs (.D(VCC_net_1), .CLK(un1_mem_0_5_85_net_1), 
        .EN(VCC_net_1), .ALn(un1_mem_0_5_132_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(VCC_net_1), .Q(
        un1_mem_0_5_132_rs_net_1));
    SLE \temp_data[3]  (.D(N_12_i_0), .CLK(FCCC_0_GL1), .EN(rd_enable), 
        .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\temp_data[3]_net_1 ));
    SLE un1_mem_0_5_139_rs (.D(VCC_net_1), .CLK(un1_mem_0_5_43_net_1), 
        .EN(VCC_net_1), .ALn(un1_mem_0_5_139_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(VCC_net_1), .Q(
        un1_mem_0_5_139_rs_net_1));
    SLE \mem_2_[6]  (.D(CoreAPB3_0_APBmslave2_PWDATA[6]), .CLK(
        FCCC_0_GL1), .EN(mem_2__1_sqmuxa), .ALn(un1_mem_0_5_150_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_2_rs[6] ));
    CFG4 #( .INIT(16'h7350) )  \temp_data_2_15_i_2[4]  (.A(
        \mem_13_[4]_net_1 ), .B(\mem_15_[4]_net_1 ), .C(N_477), .D(
        N_474), .Y(\temp_data_2_15_i_2[4]_net_1 ));
    CFG3 #( .INIT(8'hF2) )  un1_mem_0_5_192 (.A(\mem_6_[2]_net_1 ), .B(
        N_468), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_192_i));
    CFG3 #( .INIT(8'hF8) )  un1_mem_0_5_252_rs_RNIDU0M (.A(
        un1_mem_0_5_60_set_net_1), .B(un1_mem_0_5_252_rs_net_1), .C(
        \mem_15_rs[7] ), .Y(\mem_15_[7]_net_1 ));
    CFG3 #( .INIT(8'h02) )  un1_mem_0_5_124 (.A(\mem_3_[1]_net_1 ), .B(
        N_470), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_124_net_1));
    SLE \mem_1_[3]  (.D(CoreAPB3_0_APBmslave2_PWDATA[3]), .CLK(
        FCCC_0_GL1), .EN(mem_1__1_sqmuxa), .ALn(un1_mem_0_5_139_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_1_rs[3] ));
    SLE \mem_9_[3]  (.D(CoreAPB3_0_APBmslave2_PWDATA[3]), .CLK(
        FCCC_0_GL1), .EN(mem_9__1_sqmuxa), .ALn(un1_mem_0_5_181_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_9_rs[3] ));
    CFG2 #( .INIT(4'h8) )  mem_9__1_sqmuxa_0_a2 (.A(N_467), .B(
        wr_enable), .Y(mem_9__1_sqmuxa));
    CFG3 #( .INIT(8'hF2) )  un1_mem_0_5_200 (.A(\mem_6_[6]_net_1 ), .B(
        N_468), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_200_i));
    SLE \mem_4_[6]  (.D(CoreAPB3_0_APBmslave2_PWDATA[6]), .CLK(
        FCCC_0_GL1), .EN(mem_4__1_sqmuxa), .ALn(un1_mem_0_5_168_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_4_rs[6] ));
    CFG3 #( .INIT(8'h02) )  un1_mem_0_5_70 (.A(\mem_8_[6]_net_1 ), .B(
        N_479), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_70_net_1));
    CFG3 #( .INIT(8'h02) )  un1_mem_0_5_37 (.A(\mem_6_[4]_net_1 ), .B(
        N_468), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_37_net_1));
    SLE un1_mem_0_5_167_rs (.D(VCC_net_1), .CLK(un1_mem_0_5_68_net_1), 
        .EN(VCC_net_1), .ALn(un1_mem_0_5_167_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(VCC_net_1), .Q(
        un1_mem_0_5_167_rs_net_1));
    SLE un1_mem_0_5_34_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_2__1_sqmuxa), .ALn(un1_mem_0_5_34_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_mem_0_5_34_set_net_1));
    SLE un1_mem_0_5_88_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_11__1_sqmuxa), .ALn(un1_mem_0_5_88_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_mem_0_5_88_set_net_1));
    CFG3 #( .INIT(8'h02) )  un1_mem_0_5_66 (.A(\mem_8_[3]_net_1 ), .B(
        N_479), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_66_net_1));
    CFG3 #( .INIT(8'hF8) )  un1_mem_0_5_221_rs_RNI43JO (.A(
        un1_mem_0_5_5_set_net_1), .B(un1_mem_0_5_221_rs_net_1), .C(
        \mem_8_rs[1] ), .Y(\mem_8_[1]_net_1 ));
    CFG4 #( .INIT(16'h7530) )  \temp_data_2_15_i_7[5]  (.A(
        \mem_12_[5]_net_1 ), .B(\mem_8_[5]_net_1 ), .C(N_479), .D(
        N_469), .Y(\temp_data_2_15_i_7[5]_net_1 ));
    CFG3 #( .INIT(8'hF8) )  \mem_10__RNIDMMI[0]  (.A(
        un1_mem_0_5_97_set_net_1), .B(un1_mem_0_5_191_rs_net_1), .C(
        \mem_10_rs[0] ), .Y(\mem_10_[0]_net_1 ));
    CFG3 #( .INIT(8'hF8) )  un1_mem_0_5_238_rs_RNIQOHL (.A(
        un1_mem_0_5_110_set_net_1), .B(un1_mem_0_5_238_rs_net_1), .C(
        \mem_13_rs[6] ), .Y(\mem_13_[6]_net_1 ));
    SLE \data_out[7]  (.D(\temp_data[7]_net_1 ), .CLK(FCCC_0_GL1), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(
        CoreAPB3_0_APBmslave3_PRDATA[7]));
    CFG3 #( .INIT(8'hF8) )  \mem_14__RNIGAHT[0]  (.A(
        un1_mem_0_5_112_set_net_1), .B(un1_mem_0_5_240_rs_net_1), .C(
        \mem_14_rs[0] ), .Y(\mem_14_[0]_net_1 ));
    SLE un1_mem_0_5_210_rs (.D(VCC_net_1), .CLK(un1_mem_0_5_51_net_1), 
        .EN(VCC_net_1), .ALn(un1_mem_0_5_210_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(VCC_net_1), .Q(
        un1_mem_0_5_210_rs_net_1));
    SLE un1_mem_0_5_190_rs (.D(VCC_net_1), .CLK(un1_mem_0_5_31_net_1), 
        .EN(VCC_net_1), .ALn(un1_mem_0_5_190_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(VCC_net_1), .Q(
        un1_mem_0_5_190_rs_net_1));
    CFG1 #( .INIT(2'h1) )  un1_mem_0_5_50_set_RNO (.A(
        un1_mem_0_5_50_net_1), .Y(un1_mem_0_5_50_i));
    CFG2 #( .INIT(4'h8) )  mem_8__1_sqmuxa_0_a2 (.A(N_479), .B(
        wr_enable), .Y(mem_8__1_sqmuxa));
    CFG3 #( .INIT(8'h02) )  un1_mem_0_5_98 (.A(\mem_10_[1]_net_1 ), .B(
        N_471), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_98_net_1));
    CFG3 #( .INIT(8'h02) )  un1_mem_0_5_101 (.A(\mem_10_[4]_net_1 ), 
        .B(N_471), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_101_net_1));
    CFG3 #( .INIT(8'h02) )  un1_mem_0_5_99 (.A(\mem_10_[2]_net_1 ), .B(
        N_471), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_99_net_1));
    SLE un1_mem_0_5_209_rs (.D(VCC_net_1), .CLK(un1_mem_0_5_89_net_1), 
        .EN(VCC_net_1), .ALn(un1_mem_0_5_209_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(VCC_net_1), .Q(
        un1_mem_0_5_209_rs_net_1));
    CFG3 #( .INIT(8'hF8) )  un1_mem_0_5_69_set_RNIDLDH (.A(
        un1_mem_0_5_69_set_net_1), .B(un1_mem_0_5_169_rs_net_1), .C(
        \mem_8_rs[5] ), .Y(\mem_8_[5]_net_1 ));
    SLE un1_mem_0_5_177_rs (.D(VCC_net_1), .CLK(un1_mem_0_5_73_net_1), 
        .EN(VCC_net_1), .ALn(un1_mem_0_5_177_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(VCC_net_1), .Q(
        un1_mem_0_5_177_rs_net_1));
    CFG3 #( .INIT(8'hF2) )  un1_mem_0_5_163 (.A(\mem_4_[2]_net_1 ), .B(
        N_476), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_163_i));
    SLE un1_mem_0_5_50_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_3__1_sqmuxa), .ALn(un1_mem_0_5_50_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_mem_0_5_50_set_net_1));
    CFG1 #( .INIT(2'h1) )  un1_mem_0_5_13_set_RNO (.A(
        un1_mem_0_5_13_net_1), .Y(un1_mem_0_5_13_i));
    CFG1 #( .INIT(2'h1) )  un1_mem_0_5_84_set_RNO (.A(
        un1_mem_0_5_84_net_1), .Y(un1_mem_0_5_84_i));
    SLE un1_mem_0_5_231_rs (.D(VCC_net_1), .CLK(un1_mem_0_5_23_net_1), 
        .EN(VCC_net_1), .ALn(un1_mem_0_5_231_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(VCC_net_1), .Q(
        un1_mem_0_5_231_rs_net_1));
    CFG3 #( .INIT(8'hF2) )  un1_mem_0_5_248 (.A(\mem_15_[0]_net_1 ), 
        .B(N_474), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_248_i));
    CFG4 #( .INIT(16'h7350) )  \temp_data_2_15_i_4[3]  (.A(
        \mem_10_[3]_net_1 ), .B(\mem_6_[3]_net_1 ), .C(N_471), .D(
        N_468), .Y(\temp_data_2_15_i_4[3]_net_1 ));
    CFG4 #( .INIT(16'h7350) )  \temp_data_2_15_i_1[6]  (.A(
        \mem_11_[6]_net_1 ), .B(\mem_3_[6]_net_1 ), .C(N_475), .D(
        N_470), .Y(\temp_data_2_15_i_1[6]_net_1 ));
    SLE \mem_6_[4]  (.D(CoreAPB3_0_APBmslave2_PWDATA[4]), .CLK(
        FCCC_0_GL1), .EN(mem_6__1_sqmuxa), .ALn(un1_mem_0_5_196_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_6_rs[4] ));
    SLE un1_mem_0_5_235_rs (.D(VCC_net_1), .CLK(un1_mem_0_5_107_net_1), 
        .EN(VCC_net_1), .ALn(un1_mem_0_5_235_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(VCC_net_1), .Q(
        un1_mem_0_5_235_rs_net_1));
    CFG3 #( .INIT(8'hF8) )  un1_mem_0_5_24_set_RNINOSM (.A(
        un1_mem_0_5_24_set_net_1), .B(un1_mem_0_5_143_rs_net_1), .C(
        \mem_1_rs[7] ), .Y(\mem_1_[7]_net_1 ));
    CFG3 #( .INIT(8'h02) )  un1_mem_0_5_38 (.A(\mem_2_[6]_net_1 ), .B(
        N_478), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_38_net_1));
    CFG4 #( .INIT(16'h7350) )  \temp_data_2_15_i_2[2]  (.A(
        \mem_13_[2]_net_1 ), .B(\mem_15_[2]_net_1 ), .C(N_477), .D(
        N_474), .Y(\temp_data_2_15_i_2[2]_net_1 ));
    CFG4 #( .INIT(16'h2000) )  \WRITE_GEN.mem_11__2_i_a2[5]  (.A(
        CoreAPB3_0_APBmslave2_PADDR[3]), .B(
        CoreAPB3_0_APBmslave2_PADDR[2]), .C(
        CoreAPB3_0_APBmslave2_PADDR[0]), .D(
        CoreAPB3_0_APBmslave2_PADDR[1]), .Y(N_475));
    CFG3 #( .INIT(8'h02) )  un1_mem_0_5_39 (.A(\mem_6_[5]_net_1 ), .B(
        N_468), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_39_net_1));
    SLE \data_out[2]  (.D(\temp_data[2]_net_1 ), .CLK(FCCC_0_GL1), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(
        CoreAPB3_0_APBmslave3_PRDATA[2]));
    CFG3 #( .INIT(8'hF2) )  un1_mem_0_5_152 (.A(\mem_3_[0]_net_1 ), .B(
        N_470), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_152_i));
    CFG3 #( .INIT(8'h02) )  un1_mem_0_5_110 (.A(\mem_13_[6]_net_1 ), 
        .B(N_477), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_110_net_1));
    SLE un1_mem_0_5_13_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_5__1_sqmuxa), .ALn(un1_mem_0_5_13_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_mem_0_5_13_set_net_1));
    SLE un1_mem_0_5_134_rs (.D(VCC_net_1), .CLK(un1_mem_0_5_87_net_1), 
        .EN(VCC_net_1), .ALn(un1_mem_0_5_134_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(VCC_net_1), .Q(
        un1_mem_0_5_134_rs_net_1));
    CFG3 #( .INIT(8'hF8) )  \mem_3__RNI9T7Q[2]  (.A(
        un1_mem_0_5_126_set_net_1), .B(un1_mem_0_5_154_rs_net_1), .C(
        \mem_3_rs[2] ), .Y(\mem_3_[2]_net_1 ));
    CFG3 #( .INIT(8'hF8) )  \mem_14__RNI53II[7]  (.A(
        un1_mem_0_5_119_set_net_1), .B(un1_mem_0_5_247_rs_net_1), .C(
        \mem_14_rs[7] ), .Y(\mem_14_[7]_net_1 ));
    SLE un1_mem_0_5_186_rs (.D(VCC_net_1), .CLK(un1_mem_0_5_27_net_1), 
        .EN(VCC_net_1), .ALn(un1_mem_0_5_186_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(VCC_net_1), .Q(
        un1_mem_0_5_186_rs_net_1));
    SLE \mem_0_[4]  (.D(CoreAPB3_0_APBmslave2_PWDATA[4]), .CLK(
        FCCC_0_GL1), .EN(mem_0__1_sqmuxa), .ALn(un1_mem_0_5_132_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_0_rs[4] ));
    CFG3 #( .INIT(8'hF8) )  un1_mem_0_5_166_rs_RNI4KVK (.A(
        un1_mem_0_5_67_set_net_1), .B(un1_mem_0_5_166_rs_net_1), .C(
        \mem_4_rs[5] ), .Y(\mem_4_[5]_net_1 ));
    SLE un1_mem_0_5_213_rs (.D(VCC_net_1), .CLK(un1_mem_0_5_54_net_1), 
        .EN(VCC_net_1), .ALn(un1_mem_0_5_213_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(VCC_net_1), .Q(
        un1_mem_0_5_213_rs_net_1));
    CFG1 #( .INIT(2'h1) )  un1_mem_0_5_27_set_RNO (.A(
        un1_mem_0_5_27_net_1), .Y(un1_mem_0_5_27_i));
    CFG3 #( .INIT(8'hF2) )  un1_mem_0_5_249 (.A(\mem_15_[1]_net_1 ), 
        .B(N_474), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_249_i));
    CFG3 #( .INIT(8'h02) )  un1_mem_0_5_42 (.A(\mem_5_[3]_net_1 ), .B(
        N_472), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_42_net_1));
    CFG4 #( .INIT(16'h7350) )  \temp_data_2_15_i_4[0]  (.A(
        \mem_10_[0]_net_1 ), .B(\mem_6_[0]_net_1 ), .C(N_471), .D(
        N_468), .Y(\temp_data_2_15_i_4[0]_net_1 ));
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hF8) )  un1_mem_0_5_174_rs_RNIPG6V (.A(
        un1_mem_0_5_15_set_net_1), .B(un1_mem_0_5_174_rs_net_1), .C(
        \mem_5_rs[1] ), .Y(\mem_5_[1]_net_1 ));
    CFG3 #( .INIT(8'hF2) )  un1_mem_0_5_169 (.A(\mem_8_[5]_net_1 ), .B(
        N_479), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_169_i));
    CFG3 #( .INIT(8'hF2) )  un1_mem_0_5_167 (.A(\mem_8_[4]_net_1 ), .B(
        N_479), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_167_i));
    CFG3 #( .INIT(8'hF2) )  un1_mem_0_5_238 (.A(\mem_13_[6]_net_1 ), 
        .B(N_477), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_238_i));
    CFG1 #( .INIT(2'h1) )  un1_mem_0_5_25_set_RNO (.A(
        un1_mem_0_5_25_net_1), .Y(un1_mem_0_5_25_i));
    SLE un1_mem_0_5_73_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_9__1_sqmuxa), .ALn(un1_mem_0_5_73_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_mem_0_5_73_set_net_1));
    CFG4 #( .INIT(16'h7350) )  \temp_data_2_15_i_1[7]  (.A(
        \mem_11_[7]_net_1 ), .B(\mem_3_[7]_net_1 ), .C(N_475), .D(
        N_470), .Y(\temp_data_2_15_i_1[7]_net_1 ));
    SLE un1_mem_0_5_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_4__1_sqmuxa), .ALn(un1_mem_0_5_i), .ADn(GND_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_mem_0_5_set_net_1));
    CFG3 #( .INIT(8'hF2) )  un1_mem_0_5_142 (.A(\mem_1_[6]_net_1 ), .B(
        N_481), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_142_i));
    SLE \mem_12_[0]  (.D(CoreAPB3_0_APBmslave2_PWDATA[0]), .CLK(
        FCCC_0_GL1), .EN(mem_12__1_sqmuxa), .ALn(un1_mem_0_5_222_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_12_rs[0] ));
    CFG3 #( .INIT(8'hF2) )  un1_mem_0_5_253 (.A(\mem_15_[4]_net_1 ), 
        .B(N_474), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_253_i));
    SLE \mem_5_[3]  (.D(CoreAPB3_0_APBmslave2_PWDATA[3]), .CLK(
        FCCC_0_GL1), .EN(mem_5__1_sqmuxa), .ALn(un1_mem_0_5_178_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_5_rs[3] ));
    CFG4 #( .INIT(16'h0001) )  \temp_data_RNO[7]  (.A(
        \temp_data_2_15_i_4[7]_net_1 ), .B(
        \temp_data_2_15_i_5[7]_net_1 ), .C(
        \temp_data_2_15_i_11[7]_net_1 ), .D(
        \temp_data_2_15_i_12[7]_net_1 ), .Y(N_64_i_0));
    CFG3 #( .INIT(8'hF8) )  un1_mem_0_5_136_rs_RNID1TQ (.A(
        un1_mem_0_5_10_set_net_1), .B(un1_mem_0_5_136_rs_net_1), .C(
        \mem_1_rs[0] ), .Y(\mem_1_[0]_net_1 ));
    CFG4 #( .INIT(16'hFFFE) )  \temp_data_2_15_i_12[4]  (.A(
        \temp_data_2_15_i_3[4]_net_1 ), .B(
        \temp_data_2_15_i_2[4]_net_1 ), .C(
        \temp_data_2_15_i_1[4]_net_1 ), .D(
        \temp_data_2_15_i_0[4]_net_1 ), .Y(
        \temp_data_2_15_i_12[4]_net_1 ));
    SLE \mem_6_[0]  (.D(CoreAPB3_0_APBmslave2_PWDATA[0]), .CLK(
        FCCC_0_GL1), .EN(mem_6__1_sqmuxa), .ALn(un1_mem_0_5_188_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_6_rs[0] ));
    CFG3 #( .INIT(8'hF8) )  \mem_2__RNIOC1E[1]  (.A(
        un1_mem_0_5_28_set_net_1), .B(un1_mem_0_5_145_rs_net_1), .C(
        \mem_2_rs[1] ), .Y(\mem_2_[1]_net_1 ));
    SLE un1_mem_0_5_17_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_12__1_sqmuxa), .ALn(un1_mem_0_5_17_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_mem_0_5_17_set_net_1));
    CFG4 #( .INIT(16'h7350) )  \temp_data_2_15_i_5[2]  (.A(
        \mem_7_[2]_net_1 ), .B(\mem_5_[2]_net_1 ), .C(N_480), .D(N_472)
        , .Y(\temp_data_2_15_i_5[2]_net_1 ));
    SLE un1_mem_0_5_60_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_15__1_sqmuxa), .ALn(un1_mem_0_5_60_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_mem_0_5_60_set_net_1));
    CFG3 #( .INIT(8'hF2) )  un1_mem_0_5_239 (.A(\mem_13_[7]_net_1 ), 
        .B(N_477), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_239_i));
    SLE \mem_13_[5]  (.D(CoreAPB3_0_APBmslave2_PWDATA[5]), .CLK(
        FCCC_0_GL1), .EN(mem_13__1_sqmuxa), .ALn(un1_mem_0_5_237_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_13_rs[5] ));
    CFG4 #( .INIT(16'h7350) )  \temp_data_2_15_i_3[1]  (.A(
        \mem_14_[1]_net_1 ), .B(\mem_2_[1]_net_1 ), .C(N_482), .D(
        N_478), .Y(\temp_data_2_15_i_3[1]_net_1 ));
    CFG3 #( .INIT(8'hF8) )  \mem_10__RNIRVOI[4]  (.A(
        un1_mem_0_5_101_set_net_1), .B(un1_mem_0_5_199_rs_net_1), .C(
        \mem_10_rs[4] ), .Y(\mem_10_[4]_net_1 ));
    CFG3 #( .INIT(8'h02) )  un1_mem_0_5_95 (.A(\mem_11_[7]_net_1 ), .B(
        N_475), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_95_net_1));
    SLE un1_mem_0_5_83_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_3__1_sqmuxa), .ALn(un1_mem_0_5_83_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_mem_0_5_83_set_net_1));
    SLE un1_mem_0_5_148_rs (.D(VCC_net_1), .CLK(un1_mem_0_5_34_net_1), 
        .EN(VCC_net_1), .ALn(un1_mem_0_5_148_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(VCC_net_1), .Q(
        un1_mem_0_5_148_rs_net_1));
    SLE un1_mem_0_5_77_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_9__1_sqmuxa), .ALn(un1_mem_0_5_77_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_mem_0_5_77_set_net_1));
    CFG1 #( .INIT(2'h1) )  un1_mem_0_5_31_set_RNO (.A(
        un1_mem_0_5_31_net_1), .Y(un1_mem_0_5_31_i));
    CFG3 #( .INIT(8'hF2) )  un1_mem_0_5_243 (.A(\mem_14_[3]_net_1 ), 
        .B(N_482), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_243_i));
    SLE un1_mem_0_5_113_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_14__1_sqmuxa), .ALn(un1_mem_0_5_113_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_mem_0_5_113_set_net_1));
    SLE un1_mem_0_5_229_rs (.D(VCC_net_1), .CLK(un1_mem_0_5_21_net_1), 
        .EN(VCC_net_1), .ALn(un1_mem_0_5_229_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(VCC_net_1), .Q(
        un1_mem_0_5_229_rs_net_1));
    SLE \mem_0_[0]  (.D(CoreAPB3_0_APBmslave2_PWDATA[0]), .CLK(
        FCCC_0_GL1), .EN(mem_0__1_sqmuxa), .ALn(un1_mem_0_5_131_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_0_rs[0] ));
    CFG3 #( .INIT(8'hF2) )  un1_mem_0_5_132 (.A(\mem_0_[4]_net_1 ), .B(
        N_473), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_132_i));
    SLE \mem_1_[4]  (.D(CoreAPB3_0_APBmslave2_PWDATA[4]), .CLK(
        FCCC_0_GL1), .EN(mem_1__1_sqmuxa), .ALn(un1_mem_0_5_140_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_1_rs[4] ));
    CFG3 #( .INIT(8'hF8) )  \mem_2__RNIRDSQ[4]  (.A(
        un1_mem_0_5_34_set_net_1), .B(un1_mem_0_5_148_rs_net_1), .C(
        \mem_2_rs[4] ), .Y(\mem_2_[4]_net_1 ));
    SLE un1_mem_0_5_16_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_12__1_sqmuxa), .ALn(un1_mem_0_5_16_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_mem_0_5_16_set_net_1));
    SLE \mem_9_[4]  (.D(CoreAPB3_0_APBmslave2_PWDATA[4]), .CLK(
        FCCC_0_GL1), .EN(mem_9__1_sqmuxa), .ALn(un1_mem_0_5_183_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_9_rs[4] ));
    CFG1 #( .INIT(2'h1) )  un1_mem_0_5_14_set_RNO (.A(
        un1_mem_0_5_14_net_1), .Y(un1_mem_0_5_14_i));
    SLE \mem_13_[1]  (.D(CoreAPB3_0_APBmslave2_PWDATA[1]), .CLK(
        FCCC_0_GL1), .EN(mem_13__1_sqmuxa), .ALn(un1_mem_0_5_233_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_13_rs[1] ));
    SLE \mem_11_[5]  (.D(CoreAPB3_0_APBmslave2_PWDATA[5]), .CLK(
        FCCC_0_GL1), .EN(mem_11__1_sqmuxa), .ALn(un1_mem_0_5_216_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_11_rs[5] ));
    CFG3 #( .INIT(8'hF2) )  un1_mem_0_5_208 (.A(\mem_7_[2]_net_1 ), .B(
        N_480), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_208_i));
    CFG1 #( .INIT(2'h1) )  un1_mem_0_5_111_set_RNO (.A(
        un1_mem_0_5_111_net_1), .Y(un1_mem_0_5_111_i));
    CFG4 #( .INIT(16'h8000) )  \WRITE_GEN.mem_15__2_i_a2[7]  (.A(
        CoreAPB3_0_APBmslave2_PADDR[3]), .B(
        CoreAPB3_0_APBmslave2_PADDR[2]), .C(
        CoreAPB3_0_APBmslave2_PADDR[0]), .D(
        CoreAPB3_0_APBmslave2_PADDR[1]), .Y(N_474));
    CFG3 #( .INIT(8'h02) )  un1_mem_0_5_94 (.A(\mem_11_[6]_net_1 ), .B(
        N_475), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_94_net_1));
    CFG3 #( .INIT(8'hF8) )  un1_mem_0_5_77_set_RNIBIHR (.A(
        un1_mem_0_5_77_set_net_1), .B(un1_mem_0_5_185_rs_net_1), .C(
        \mem_9_rs[5] ), .Y(\mem_9_[5]_net_1 ));
    SLE un1_mem_0_5_52_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_3__1_sqmuxa), .ALn(un1_mem_0_5_52_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_mem_0_5_52_set_net_1));
    CFG1 #( .INIT(2'h1) )  un1_mem_0_5_73_set_RNO (.A(
        un1_mem_0_5_73_net_1), .Y(un1_mem_0_5_73_i));
    CFG3 #( .INIT(8'hF8) )  \mem_12__RNICSF41[3]  (.A(
        un1_mem_0_5_19_set_net_1), .B(un1_mem_0_5_227_rs_net_1), .C(
        \mem_12_rs[3] ), .Y(\mem_12_[3]_net_1 ));
    CFG1 #( .INIT(2'h1) )  un1_mem_0_5_29_set_RNO (.A(
        un1_mem_0_5_29_net_1), .Y(un1_mem_0_5_29_i));
    CFG1 #( .INIT(2'h1) )  un1_mem_0_5_41_set_RNO (.A(
        un1_mem_0_5_41_net_1), .Y(un1_mem_0_5_41_i));
    CFG3 #( .INIT(8'h02) )  un1_mem_0_5_35 (.A(\mem_6_[3]_net_1 ), .B(
        N_468), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_35_net_1));
    SLE un1_mem_0_5_76_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_9__1_sqmuxa), .ALn(un1_mem_0_5_76_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_mem_0_5_76_set_net_1));
    CFG3 #( .INIT(8'h02) )  un1_mem_0_5_8 (.A(\mem_0_[7]_net_1 ), .B(
        N_473), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_8_net_1));
    CFG3 #( .INIT(8'hF8) )  un1_mem_0_5_25_set_RNI0VMT (.A(
        un1_mem_0_5_25_set_net_1), .B(un1_mem_0_5_184_rs_net_1), .C(
        \mem_5_rs[6] ), .Y(\mem_5_[6]_net_1 ));
    SLE un1_mem_0_5_4_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_4__1_sqmuxa), .ALn(un1_mem_0_5_4_i), .ADn(GND_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_mem_0_5_4_set_net_1));
    CFG1 #( .INIT(2'h1) )  un1_mem_0_5_122_set_RNO (.A(
        un1_mem_0_5_122_net_1), .Y(un1_mem_0_5_122_i));
    SLE un1_mem_0_5_87_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_0__1_sqmuxa), .ALn(un1_mem_0_5_87_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_mem_0_5_87_set_net_1));
    SLE \mem_11_[1]  (.D(CoreAPB3_0_APBmslave2_PWDATA[1]), .CLK(
        FCCC_0_GL1), .EN(mem_11__1_sqmuxa), .ALn(un1_mem_0_5_209_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_11_rs[1] ));
    SLE un1_mem_0_5_55_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_3__1_sqmuxa), .ALn(un1_mem_0_5_55_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_mem_0_5_55_set_net_1));
    CFG3 #( .INIT(8'hF2) )  un1_mem_0_5_233 (.A(\mem_13_[1]_net_1 ), 
        .B(N_477), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_233_i));
    CFG3 #( .INIT(8'hF2) )  un1_mem_0_5_164 (.A(\mem_4_[3]_net_1 ), .B(
        N_476), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_164_i));
    CFG3 #( .INIT(8'hF2) )  un1_mem_0_5_209 (.A(\mem_11_[1]_net_1 ), 
        .B(N_475), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_209_i));
    CFG3 #( .INIT(8'hF2) )  un1_mem_0_5_170 (.A(\mem_4_[7]_net_1 ), .B(
        N_476), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_170_i));
    CFG3 #( .INIT(8'h02) )  un1_mem_0_5_115 (.A(\mem_14_[3]_net_1 ), 
        .B(N_482), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_115_net_1));
    CFG3 #( .INIT(8'hF8) )  \mem_7__RNI1ELO[2]  (.A(
        un1_mem_0_5_49_set_net_1), .B(un1_mem_0_5_208_rs_net_1), .C(
        \mem_7_rs[2] ), .Y(\mem_7_[2]_net_1 ));
    CFG4 #( .INIT(16'h7350) )  \temp_data_2_15_i_1[1]  (.A(
        \mem_11_[1]_net_1 ), .B(\mem_3_[1]_net_1 ), .C(N_475), .D(
        N_470), .Y(\temp_data_2_15_i_1[1]_net_1 ));
    CFG3 #( .INIT(8'h02) )  un1_mem_0_5_34 (.A(\mem_2_[4]_net_1 ), .B(
        N_478), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_34_net_1));
    CFG3 #( .INIT(8'h02) )  un1_mem_0_5_93 (.A(\mem_11_[5]_net_1 ), .B(
        N_475), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_93_net_1));
    CFG1 #( .INIT(2'h1) )  un1_mem_0_5_101_set_RNO (.A(
        un1_mem_0_5_101_net_1), .Y(un1_mem_0_5_101_i));
    CFG3 #( .INIT(8'hF8) )  un1_mem_0_5_4_set_RNI519S (.A(
        un1_mem_0_5_4_set_net_1), .B(un1_mem_0_5_163_rs_net_1), .C(
        \mem_4_rs[2] ), .Y(\mem_4_[2]_net_1 ));
    SLE un1_mem_0_5_86_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_0__1_sqmuxa), .ALn(un1_mem_0_5_86_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_mem_0_5_86_set_net_1));
    CFG1 #( .INIT(2'h1) )  un1_mem_0_5_56_set_RNO (.A(
        un1_mem_0_5_56_net_1), .Y(un1_mem_0_5_56_i));
    SLE \mem_1_[0]  (.D(CoreAPB3_0_APBmslave2_PWDATA[0]), .CLK(
        FCCC_0_GL1), .EN(mem_1__1_sqmuxa), .ALn(un1_mem_0_5_136_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_1_rs[0] ));
    CFG4 #( .INIT(16'h0200) )  \WRITE_GEN.mem_10__2_i_a2[7]  (.A(
        CoreAPB3_0_APBmslave2_PADDR[3]), .B(
        CoreAPB3_0_APBmslave2_PADDR[2]), .C(
        CoreAPB3_0_APBmslave2_PADDR[0]), .D(
        CoreAPB3_0_APBmslave2_PADDR[1]), .Y(N_471));
    CFG3 #( .INIT(8'h02) )  un1_mem_0_5_102 (.A(\mem_10_[5]_net_1 ), 
        .B(N_471), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_102_net_1));
    CFG3 #( .INIT(8'hF8) )  un1_mem_0_5_133_rs_RNIRKPK (.A(
        un1_mem_0_5_86_set_net_1), .B(un1_mem_0_5_133_rs_net_1), .C(
        \mem_0_rs[5] ), .Y(\mem_0_[5]_net_1 ));
    SLE \mem_9_[0]  (.D(CoreAPB3_0_APBmslave2_PWDATA[0]), .CLK(
        FCCC_0_GL1), .EN(mem_9__1_sqmuxa), .ALn(un1_mem_0_5_175_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_9_rs[0] ));
    SLE un1_mem_0_5_38_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_2__1_sqmuxa), .ALn(un1_mem_0_5_38_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_mem_0_5_38_set_net_1));
    CFG3 #( .INIT(8'hF8) )  \mem_3__RNITLDU[5]  (.A(
        un1_mem_0_5_52_set_net_1), .B(un1_mem_0_5_157_rs_net_1), .C(
        \mem_3_rs[5] ), .Y(\mem_3_[5]_net_1 ));
    CFG3 #( .INIT(8'hF8) )  un1_mem_0_5_47_set_RNIO6TL (.A(
        un1_mem_0_5_47_set_net_1), .B(un1_mem_0_5_141_rs_net_1), .C(
        \mem_1_rs[5] ), .Y(\mem_1_[5]_net_1 ));
    SLE un1_mem_0_5_244_rs (.D(VCC_net_1), .CLK(un1_mem_0_5_116_net_1), 
        .EN(VCC_net_1), .ALn(un1_mem_0_5_244_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(VCC_net_1), .Q(
        un1_mem_0_5_244_rs_net_1));
    CFG1 #( .INIT(2'h1) )  un1_mem_0_5_58_set_RNO (.A(
        un1_mem_0_5_58_net_1), .Y(un1_mem_0_5_58_i));
    SLE un1_mem_0_5_156_rs (.D(VCC_net_1), .CLK(un1_mem_0_5_50_net_1), 
        .EN(VCC_net_1), .ALn(un1_mem_0_5_156_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(VCC_net_1), .Q(
        un1_mem_0_5_156_rs_net_1));
    SLE \mem_15_[3]  (.D(CoreAPB3_0_APBmslave2_PWDATA[3]), .CLK(
        FCCC_0_GL1), .EN(mem_15__1_sqmuxa), .ALn(un1_mem_0_5_251_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_15_rs[3] ));
    SLE \mem_14_[4]  (.D(CoreAPB3_0_APBmslave2_PWDATA[4]), .CLK(
        FCCC_0_GL1), .EN(mem_14__1_sqmuxa), .ALn(un1_mem_0_5_244_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_14_rs[4] ));
    CFG3 #( .INIT(8'hF8) )  un1_mem_0_5_182_rs_RNI06B41 (.A(
        un1_mem_0_5_46_set_net_1), .B(un1_mem_0_5_182_rs_net_1), .C(
        \mem_5_rs[5] ), .Y(\mem_5_[5]_net_1 ));
    CFG1 #( .INIT(2'h1) )  un1_mem_0_5_20_set_RNO (.A(
        un1_mem_0_5_20_net_1), .Y(un1_mem_0_5_20_i));
    SLE \mem_10_[2]  (.D(CoreAPB3_0_APBmslave2_PWDATA[2]), .CLK(
        FCCC_0_GL1), .EN(mem_10__1_sqmuxa), .ALn(un1_mem_0_5_195_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_10_rs[2] ));
    SLE un1_mem_0_5_3_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_7__1_sqmuxa), .ALn(un1_mem_0_5_3_i), .ADn(GND_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_mem_0_5_3_set_net_1));
    SLE un1_mem_0_5_218_rs (.D(VCC_net_1), .CLK(un1_mem_0_5_94_net_1), 
        .EN(VCC_net_1), .ALn(un1_mem_0_5_218_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(VCC_net_1), .Q(
        un1_mem_0_5_218_rs_net_1));
    CFG3 #( .INIT(8'h02) )  un1_mem_0_5_33 (.A(\mem_6_[2]_net_1 ), .B(
        N_468), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_33_net_1));
    SLE un1_mem_0_5_138_rs (.D(VCC_net_1), .CLK(un1_mem_0_5_14_net_1), 
        .EN(VCC_net_1), .ALn(un1_mem_0_5_138_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(VCC_net_1), .Q(
        un1_mem_0_5_138_rs_net_1));
    SLE un1_mem_0_5_123_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_6__1_sqmuxa), .ALn(un1_mem_0_5_123_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_mem_0_5_123_set_net_1));
    CFG1 #( .INIT(2'h1) )  un1_mem_0_5_5_set_RNO (.A(
        un1_mem_0_5_5_net_1), .Y(un1_mem_0_5_5_i));
    CFG3 #( .INIT(8'hF2) )  un1_mem_0_5_211 (.A(\mem_11_[2]_net_1 ), 
        .B(N_475), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_211_i));
    SLE un1_mem_0_5_62_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_15__1_sqmuxa), .ALn(un1_mem_0_5_62_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_mem_0_5_62_set_net_1));
    SLE un1_mem_0_5_165_rs (.D(VCC_net_1), .CLK(un1_mem_0_5_65_net_1), 
        .EN(VCC_net_1), .ALn(un1_mem_0_5_165_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(VCC_net_1), .Q(
        un1_mem_0_5_165_rs_net_1));
    SLE un1_mem_0_5_217_rs (.D(VCC_net_1), .CLK(un1_mem_0_5_1_net_1), 
        .EN(VCC_net_1), .ALn(un1_mem_0_5_217_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(VCC_net_1), .Q(
        un1_mem_0_5_217_rs_net_1));
    CFG3 #( .INIT(8'hF8) )  un1_mem_0_5_180_rs_RNIRMOP (.A(
        un1_mem_0_5_44_set_net_1), .B(un1_mem_0_5_180_rs_net_1), .C(
        \mem_5_rs[4] ), .Y(\mem_5_[4]_net_1 ));
    SLE \mem_3_[2]  (.D(CoreAPB3_0_APBmslave2_PWDATA[2]), .CLK(
        FCCC_0_GL1), .EN(mem_3__1_sqmuxa), .ALn(un1_mem_0_5_154_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_3_rs[2] ));
    CFG3 #( .INIT(8'hF2) )  un1_mem_0_5_203 (.A(\mem_10_[6]_net_1 ), 
        .B(N_471), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_203_i));
    SLE un1_mem_0_5_41_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_1__1_sqmuxa), .ALn(un1_mem_0_5_41_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_mem_0_5_41_set_net_1));
    SLE un1_mem_0_5_161_rs (.D(VCC_net_1), .CLK(un1_mem_0_5_net_1), 
        .EN(VCC_net_1), .ALn(un1_mem_0_5_161_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(VCC_net_1), .Q(
        un1_mem_0_5_161_rs_net_1));
    SLE \mem_14_[6]  (.D(CoreAPB3_0_APBmslave2_PWDATA[6]), .CLK(
        FCCC_0_GL1), .EN(mem_14__1_sqmuxa), .ALn(un1_mem_0_5_246_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_14_rs[6] ));
    CFG3 #( .INIT(8'h02) )  un1_mem_0_5_22 (.A(\mem_12_[6]_net_1 ), .B(
        N_469), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_22_net_1));
    CFG3 #( .INIT(8'hF8) )  un1_mem_0_5_206_rs_RNIB7OM (.A(
        un1_mem_0_5_127_set_net_1), .B(un1_mem_0_5_206_rs_net_1), .C(
        \mem_7_rs[1] ), .Y(\mem_7_[1]_net_1 ));
    CFG3 #( .INIT(8'hF8) )  un1_mem_0_5_18_set_RNI9K6V (.A(
        un1_mem_0_5_18_set_net_1), .B(un1_mem_0_5_226_rs_net_1), .C(
        \mem_12_rs[2] ), .Y(\mem_12_[2]_net_1 ));
    CFG3 #( .INIT(8'hF2) )  un1_mem_0_5_217 (.A(\mem_7_[7]_net_1 ), .B(
        N_480), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_217_i));
    CFG3 #( .INIT(8'hF2) )  un1_mem_0_5_180 (.A(\mem_5_[4]_net_1 ), .B(
        N_472), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_180_i));
    SLE un1_mem_0_5_65_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_4__1_sqmuxa), .ALn(un1_mem_0_5_65_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_mem_0_5_65_set_net_1));
    CFG3 #( .INIT(8'h02) )  un1_mem_0_5_90 (.A(\mem_11_[2]_net_1 ), .B(
        N_475), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_90_net_1));
    CFG1 #( .INIT(2'h1) )  un1_mem_0_5_74_set_RNO (.A(
        un1_mem_0_5_74_net_1), .Y(un1_mem_0_5_74_i));
    CFG3 #( .INIT(8'hF2) )  un1_mem_0_5_190 (.A(\mem_6_[1]_net_1 ), .B(
        N_468), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_190_i));
    CFG3 #( .INIT(8'h02) )  un1_mem_0_5_61 (.A(\mem_15_[3]_net_1 ), .B(
        N_474), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_61_net_1));
    SLE \mem_8_[7]  (.D(CoreAPB3_0_APBmslave2_PWDATA[7]), .CLK(
        FCCC_0_GL1), .EN(mem_8__1_sqmuxa), .ALn(un1_mem_0_5_173_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_8_rs[7] ));
    SLE un1_mem_0_5_104_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_13__1_sqmuxa), .ALn(un1_mem_0_5_104_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_mem_0_5_104_set_net_1));
    SLE \mem_5_[4]  (.D(CoreAPB3_0_APBmslave2_PWDATA[4]), .CLK(
        FCCC_0_GL1), .EN(mem_5__1_sqmuxa), .ALn(un1_mem_0_5_180_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_5_rs[4] ));
    CFG3 #( .INIT(8'h02) )  un1_mem_0_5_1 (.A(\mem_7_[7]_net_1 ), .B(
        N_480), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_1_net_1));
    CFG4 #( .INIT(16'h0100) )  \WRITE_GEN.mem_2__2_i_a2[7]  (.A(
        CoreAPB3_0_APBmslave2_PADDR[3]), .B(
        CoreAPB3_0_APBmslave2_PADDR[2]), .C(
        CoreAPB3_0_APBmslave2_PADDR[0]), .D(
        CoreAPB3_0_APBmslave2_PADDR[1]), .Y(N_478));
    CFG1 #( .INIT(2'h1) )  un1_mem_0_5_52_set_RNO (.A(
        un1_mem_0_5_52_net_1), .Y(un1_mem_0_5_52_i));
    SLE un1_mem_0_5_175_rs (.D(VCC_net_1), .CLK(un1_mem_0_5_72_net_1), 
        .EN(VCC_net_1), .ALn(un1_mem_0_5_175_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(VCC_net_1), .Q(
        un1_mem_0_5_175_rs_net_1));
    SLE \data_out[1]  (.D(\temp_data[1]_net_1 ), .CLK(FCCC_0_GL1), .EN(
        VCC_net_1), .ALn(VCC_net_1), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(
        CoreAPB3_0_APBmslave3_PRDATA[1]));
    SLE \mem_8_[5]  (.D(CoreAPB3_0_APBmslave2_PWDATA[5]), .CLK(
        FCCC_0_GL1), .EN(mem_8__1_sqmuxa), .ALn(un1_mem_0_5_169_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_8_rs[5] ));
    CFG3 #( .INIT(8'h02) )  un1_mem_0_5_46 (.A(\mem_5_[5]_net_1 ), .B(
        N_472), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_46_net_1));
    SLE un1_mem_0_5_183_rs (.D(VCC_net_1), .CLK(un1_mem_0_5_76_net_1), 
        .EN(VCC_net_1), .ALn(un1_mem_0_5_183_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(VCC_net_1), .Q(
        un1_mem_0_5_183_rs_net_1));
    CFG3 #( .INIT(8'h02) )  un1_mem_0_5_52 (.A(\mem_3_[5]_net_1 ), .B(
        N_470), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_52_net_1));
    CFG4 #( .INIT(16'h0001) )  \temp_data_RNO[2]  (.A(
        \temp_data_2_15_i_4[2]_net_1 ), .B(
        \temp_data_2_15_i_5[2]_net_1 ), .C(
        \temp_data_2_15_i_11[2]_net_1 ), .D(
        \temp_data_2_15_i_12[2]_net_1 ), .Y(N_10_i_0));
    SLE un1_mem_0_5_59_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_15__1_sqmuxa), .ALn(un1_mem_0_5_59_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_mem_0_5_59_set_net_1));
    SLE un1_mem_0_5_171_rs (.D(VCC_net_1), .CLK(un1_mem_0_5_70_net_1), 
        .EN(VCC_net_1), .ALn(un1_mem_0_5_171_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(VCC_net_1), .Q(
        un1_mem_0_5_171_rs_net_1));
    CFG3 #( .INIT(8'hF8) )  un1_mem_0_5_20_set_RNI616Q (.A(
        un1_mem_0_5_20_set_net_1), .B(un1_mem_0_5_228_rs_net_1), .C(
        \mem_12_rs[4] ), .Y(\mem_12_[4]_net_1 ));
    CFG3 #( .INIT(8'hF8) )  un1_mem_0_5_50_set_RNIP9UK (.A(
        un1_mem_0_5_50_set_net_1), .B(un1_mem_0_5_156_rs_net_1), .C(
        \mem_3_rs[4] ), .Y(\mem_3_[4]_net_1 ));
    SLE un1_mem_0_5_90_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_11__1_sqmuxa), .ALn(un1_mem_0_5_90_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_mem_0_5_90_set_net_1));
    CFG3 #( .INIT(8'h02) )  un1_mem_0_5_30 (.A(\mem_2_[2]_net_1 ), .B(
        N_478), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_30_net_1));
    SLE un1_mem_0_5_20_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_12__1_sqmuxa), .ALn(un1_mem_0_5_20_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_mem_0_5_20_set_net_1));
    CFG3 #( .INIT(8'h02) )  un1_mem_0_5_113 (.A(\mem_14_[1]_net_1 ), 
        .B(N_482), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_113_net_1));
    CFG3 #( .INIT(8'hF2) )  un1_mem_0_5_175 (.A(\mem_9_[0]_net_1 ), .B(
        N_467), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_175_i));
    SLE un1_mem_0_5_196_rs (.D(VCC_net_1), .CLK(un1_mem_0_5_37_net_1), 
        .EN(VCC_net_1), .ALn(un1_mem_0_5_196_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(VCC_net_1), .Q(
        un1_mem_0_5_196_rs_net_1));
    CFG3 #( .INIT(8'hF8) )  \mem_6__RNIRPQL[2]  (.A(
        un1_mem_0_5_33_set_net_1), .B(un1_mem_0_5_192_rs_net_1), .C(
        \mem_6_rs[2] ), .Y(\mem_6_[2]_net_1 ));
    SLE un1_mem_0_5_162_rs (.D(VCC_net_1), .CLK(un1_mem_0_5_2_net_1), 
        .EN(VCC_net_1), .ALn(un1_mem_0_5_162_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(VCC_net_1), .Q(
        un1_mem_0_5_162_rs_net_1));
    CFG4 #( .INIT(16'h7350) )  \temp_data_2_15_i_5[3]  (.A(
        \mem_7_[3]_net_1 ), .B(\mem_5_[3]_net_1 ), .C(N_480), .D(N_472)
        , .Y(\temp_data_2_15_i_5[3]_net_1 ));
    CFG2 #( .INIT(4'h8) )  mem_6__1_sqmuxa_0_a2 (.A(N_468), .B(
        wr_enable), .Y(mem_6__1_sqmuxa));
    SLE un1_mem_0_5_169_rs (.D(VCC_net_1), .CLK(un1_mem_0_5_69_net_1), 
        .EN(VCC_net_1), .ALn(un1_mem_0_5_169_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(VCC_net_1), .Q(
        un1_mem_0_5_169_rs_net_1));
    CFG3 #( .INIT(8'hF8) )  un1_mem_0_5_168_rs_RNIJ8NM (.A(
        un1_mem_0_5_9_set_net_1), .B(un1_mem_0_5_168_rs_net_1), .C(
        \mem_4_rs[6] ), .Y(\mem_4_[6]_net_1 ));
    SLE un1_mem_0_5_234_rs (.D(VCC_net_1), .CLK(un1_mem_0_5_106_net_1), 
        .EN(VCC_net_1), .ALn(un1_mem_0_5_234_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(VCC_net_1), .Q(
        un1_mem_0_5_234_rs_net_1));
    CFG2 #( .INIT(4'h2) )  \temp_data_2_15_i_a2_13[4]  (.A(N_476), .B(
        \mem_4_[4]_net_1 ), .Y(N_393));
    CFG3 #( .INIT(8'hF8) )  \mem_6__RNI8DDT[7]  (.A(
        un1_mem_0_5_123_set_net_1), .B(un1_mem_0_5_202_rs_net_1), .C(
        \mem_6_rs[7] ), .Y(\mem_6_[7]_net_1 ));
    SLE un1_mem_0_5_246_rs (.D(VCC_net_1), .CLK(un1_mem_0_5_118_net_1), 
        .EN(VCC_net_1), .ALn(un1_mem_0_5_246_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(VCC_net_1), .Q(
        un1_mem_0_5_246_rs_net_1));
    CFG3 #( .INIT(8'hF8) )  \mem_2__RNIK0IK[0]  (.A(
        un1_mem_0_5_26_set_net_1), .B(un1_mem_0_5_144_rs_net_1), .C(
        \mem_2_rs[0] ), .Y(\mem_2_[0]_net_1 ));
    SLE un1_mem_0_5_102_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_10__1_sqmuxa), .ALn(un1_mem_0_5_102_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_mem_0_5_102_set_net_1));
    CFG4 #( .INIT(16'h7530) )  \temp_data_2_15_i_0[5]  (.A(
        \mem_9_[5]_net_1 ), .B(\mem_1_[5]_net_1 ), .C(N_481), .D(N_467)
        , .Y(\temp_data_2_15_i_0[5]_net_1 ));
    CFG4 #( .INIT(16'h7530) )  \temp_data_2_15_i_0[1]  (.A(
        \mem_9_[1]_net_1 ), .B(\mem_1_[1]_net_1 ), .C(N_481), .D(N_467)
        , .Y(\temp_data_2_15_i_0[1]_net_1 ));
    CFG3 #( .INIT(8'hF8) )  un1_mem_0_5_171_rs_RNIV2EH (.A(
        un1_mem_0_5_70_set_net_1), .B(un1_mem_0_5_171_rs_net_1), .C(
        \mem_8_rs[6] ), .Y(\mem_8_[6]_net_1 ));
    SLE \mem_5_[0]  (.D(CoreAPB3_0_APBmslave2_PWDATA[0]), .CLK(
        FCCC_0_GL1), .EN(mem_5__1_sqmuxa), .ALn(un1_mem_0_5_172_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_5_rs[0] ));
    CFG4 #( .INIT(16'hEFEE) )  \temp_data_2_15_i_11[4]  (.A(N_393), .B(
        \temp_data_2_15_i_7[4]_net_1 ), .C(\mem_0_[4]_net_1 ), .D(
        N_473), .Y(\temp_data_2_15_i_11[4]_net_1 ));
    SLE \mem_3_[1]  (.D(CoreAPB3_0_APBmslave2_PWDATA[1]), .CLK(
        FCCC_0_GL1), .EN(mem_3__1_sqmuxa), .ALn(un1_mem_0_5_153_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_3_rs[1] ));
    CFG1 #( .INIT(2'h1) )  un1_mem_0_5_33_set_RNO (.A(
        un1_mem_0_5_33_net_1), .Y(un1_mem_0_5_33_i));
    SLE un1_mem_0_5_33_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_6__1_sqmuxa), .ALn(un1_mem_0_5_33_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_mem_0_5_33_set_net_1));
    CFG3 #( .INIT(8'hF8) )  un1_mem_0_5_211_rs_RNI25BI (.A(
        un1_mem_0_5_90_set_net_1), .B(un1_mem_0_5_211_rs_net_1), .C(
        \mem_11_rs[2] ), .Y(\mem_11_[2]_net_1 ));
    CFG1 #( .INIT(2'h1) )  un1_mem_0_5_97_set_RNO (.A(
        un1_mem_0_5_97_net_1), .Y(un1_mem_0_5_97_i));
    CFG3 #( .INIT(8'h02) )  un1_mem_0_5_119 (.A(\mem_14_[7]_net_1 ), 
        .B(N_482), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_119_net_1));
    CFG3 #( .INIT(8'h02) )  un1_mem_0_5_117 (.A(\mem_14_[5]_net_1 ), 
        .B(N_482), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_117_net_1));
    CFG3 #( .INIT(8'hF2) )  un1_mem_0_5_224 (.A(\mem_12_[1]_net_1 ), 
        .B(N_469), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_224_i));
    SLE un1_mem_0_5_172_rs (.D(VCC_net_1), .CLK(un1_mem_0_5_13_net_1), 
        .EN(VCC_net_1), .ALn(un1_mem_0_5_172_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(VCC_net_1), .Q(
        un1_mem_0_5_172_rs_net_1));
    CFG4 #( .INIT(16'h7350) )  \temp_data_2_15_i_3[5]  (.A(
        \mem_14_[5]_net_1 ), .B(\mem_2_[5]_net_1 ), .C(N_482), .D(
        N_478), .Y(\temp_data_2_15_i_3[5]_net_1 ));
    CFG4 #( .INIT(16'h7350) )  \temp_data_2_15_i_5[4]  (.A(
        \mem_7_[4]_net_1 ), .B(\mem_5_[4]_net_1 ), .C(N_480), .D(N_472)
        , .Y(\temp_data_2_15_i_5[4]_net_1 ));
    SLE un1_mem_0_5_179_rs (.D(VCC_net_1), .CLK(un1_mem_0_5_74_net_1), 
        .EN(VCC_net_1), .ALn(un1_mem_0_5_179_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(VCC_net_1), .Q(
        un1_mem_0_5_179_rs_net_1));
    CFG1 #( .INIT(2'h1) )  un1_mem_0_5_95_set_RNO (.A(
        un1_mem_0_5_95_net_1), .Y(un1_mem_0_5_95_i));
    CFG3 #( .INIT(8'hF8) )  un1_mem_0_5_16_set_RNI1UDI (.A(
        un1_mem_0_5_16_set_net_1), .B(un1_mem_0_5_222_rs_net_1), .C(
        \mem_12_rs[0] ), .Y(\mem_12_[0]_net_1 ));
    CFG3 #( .INIT(8'hF2) )  un1_mem_0_5_150 (.A(\mem_2_[6]_net_1 ), .B(
        N_478), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_150_i));
    CFG3 #( .INIT(8'hF2) )  un1_mem_0_5_128 (.A(\mem_0_[1]_net_1 ), .B(
        N_473), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_128_i));
    SLE \mem_10_[7]  (.D(CoreAPB3_0_APBmslave2_PWDATA[7]), .CLK(
        FCCC_0_GL1), .EN(mem_10__1_sqmuxa), .ALn(un1_mem_0_5_205_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_10_rs[7] ));
    CFG1 #( .INIT(2'h1) )  un1_mem_0_5_43_set_RNO (.A(
        un1_mem_0_5_43_net_1), .Y(un1_mem_0_5_43_i));
    SLE un1_mem_0_5_69_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_8__1_sqmuxa), .ALn(un1_mem_0_5_69_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_mem_0_5_69_set_net_1));
    CFG1 #( .INIT(2'h1) )  un1_mem_0_5_61_set_RNO (.A(
        un1_mem_0_5_61_net_1), .Y(un1_mem_0_5_61_i));
    SLE \mem_15_[0]  (.D(CoreAPB3_0_APBmslave2_PWDATA[0]), .CLK(
        FCCC_0_GL1), .EN(mem_15__1_sqmuxa), .ALn(un1_mem_0_5_248_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_15_rs[0] ));
    CFG3 #( .INIT(8'hF2) )  un1_mem_0_5_185 (.A(\mem_9_[5]_net_1 ), .B(
        N_467), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_185_i));
    SLE un1_mem_0_5_2_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_4__1_sqmuxa), .ALn(un1_mem_0_5_2_i), .ADn(GND_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_mem_0_5_2_set_net_1));
    CFG3 #( .INIT(8'hF8) )  un1_mem_0_5_81_set_RNIM74H (.A(
        un1_mem_0_5_81_set_net_1), .B(un1_mem_0_5_128_rs_net_1), .C(
        \mem_0_rs[1] ), .Y(\mem_0_[1]_net_1 ));
    CFG3 #( .INIT(8'h02) )  un1_mem_0_5_7 (.A(\mem_8_[0]_net_1 ), .B(
        N_479), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_7_net_1));
    SLE un1_mem_0_5_44_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_5__1_sqmuxa), .ALn(un1_mem_0_5_44_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_mem_0_5_44_set_net_1));
    CFG3 #( .INIT(8'h02) )  un1_mem_0_5_67 (.A(\mem_4_[5]_net_1 ), .B(
        N_476), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_67_net_1));
    CFG3 #( .INIT(8'hF2) )  un1_mem_0_5_195 (.A(\mem_10_[2]_net_1 ), 
        .B(N_471), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_195_i));
    CFG3 #( .INIT(8'hF8) )  un1_mem_0_5_165_rs_RNI08GR (.A(
        un1_mem_0_5_65_set_net_1), .B(un1_mem_0_5_165_rs_net_1), .C(
        \mem_4_rs[4] ), .Y(\mem_4_[4]_net_1 ));
    CFG1 #( .INIT(2'h1) )  un1_mem_0_5_3_set_RNO (.A(
        un1_mem_0_5_3_net_1), .Y(un1_mem_0_5_3_i));
    SLE un1_mem_0_5_37_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_6__1_sqmuxa), .ALn(un1_mem_0_5_37_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_mem_0_5_37_set_net_1));
    CFG3 #( .INIT(8'hF2) )  un1_mem_0_5_140 (.A(\mem_1_[4]_net_1 ), .B(
        N_481), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_140_i));
    CFG3 #( .INIT(8'hF8) )  \mem_10__RNIDDPI[5]  (.A(
        un1_mem_0_5_102_set_net_1), .B(un1_mem_0_5_201_rs_net_1), .C(
        \mem_10_rs[5] ), .Y(\mem_10_[5]_net_1 ));
    SLE un1_mem_0_5_242_rs (.D(VCC_net_1), .CLK(un1_mem_0_5_114_net_1), 
        .EN(VCC_net_1), .ALn(un1_mem_0_5_242_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(VCC_net_1), .Q(
        un1_mem_0_5_242_rs_net_1));
    CFG1 #( .INIT(2'h1) )  un1_mem_0_5_113_set_RNO (.A(
        un1_mem_0_5_113_net_1), .Y(un1_mem_0_5_113_i));
    CFG4 #( .INIT(16'h7350) )  \temp_data_2_15_i_5[6]  (.A(
        \mem_7_[6]_net_1 ), .B(\mem_5_[6]_net_1 ), .C(N_480), .D(N_472)
        , .Y(\temp_data_2_15_i_5[6]_net_1 ));
    CFG3 #( .INIT(8'hF2) )  un1_mem_0_5_216 (.A(\mem_11_[5]_net_1 ), 
        .B(N_475), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_216_i));
    CFG2 #( .INIT(4'h8) )  mem_1__1_sqmuxa_0_a2 (.A(N_481), .B(
        wr_enable), .Y(mem_1__1_sqmuxa));
    SLE un1_mem_0_5_92_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_11__1_sqmuxa), .ALn(un1_mem_0_5_92_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_mem_0_5_92_set_net_1));
    CFG4 #( .INIT(16'hEFEE) )  \temp_data_2_15_i_11[2]  (.A(N_361), .B(
        \temp_data_2_15_i_7[2]_net_1 ), .C(\mem_0_[2]_net_1 ), .D(
        N_473), .Y(\temp_data_2_15_i_11[2]_net_1 ));
    SLE \temp_data[1]  (.D(N_8_i_0), .CLK(FCCC_0_GL1), .EN(rd_enable), 
        .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\temp_data[1]_net_1 ));
    SLE un1_mem_0_5_140_rs (.D(VCC_net_1), .CLK(un1_mem_0_5_41_net_1), 
        .EN(VCC_net_1), .ALn(un1_mem_0_5_140_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(VCC_net_1), .Q(
        un1_mem_0_5_140_rs_net_1));
    SLE un1_mem_0_5_164_rs (.D(VCC_net_1), .CLK(un1_mem_0_5_6_net_1), 
        .EN(VCC_net_1), .ALn(un1_mem_0_5_164_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(VCC_net_1), .Q(
        un1_mem_0_5_164_rs_net_1));
    SLE \temp_data[0]  (.D(N_4_i_0), .CLK(FCCC_0_GL1), .EN(rd_enable), 
        .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\temp_data[0]_net_1 ));
    SLE un1_mem_0_5_36_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_2__1_sqmuxa), .ALn(un1_mem_0_5_36_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_mem_0_5_36_set_net_1));
    CFG4 #( .INIT(16'h7350) )  \temp_data_2_15_i_4[6]  (.A(
        \mem_10_[6]_net_1 ), .B(\mem_6_[6]_net_1 ), .C(N_471), .D(
        N_468), .Y(\temp_data_2_15_i_4[6]_net_1 ));
    CFG1 #( .INIT(2'h1) )  un1_mem_0_5_87_set_RNO (.A(
        un1_mem_0_5_87_net_1), .Y(un1_mem_0_5_87_i));
    SLE un1_mem_0_5_22_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_12__1_sqmuxa), .ALn(un1_mem_0_5_22_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_mem_0_5_22_set_net_1));
    CFG1 #( .INIT(2'h1) )  un1_mem_0_5_26_set_RNO (.A(
        un1_mem_0_5_26_net_1), .Y(un1_mem_0_5_26_i));
    CFG4 #( .INIT(16'h7530) )  \temp_data_2_15_i_7[1]  (.A(
        \mem_12_[1]_net_1 ), .B(\mem_8_[1]_net_1 ), .C(N_479), .D(
        N_469), .Y(\temp_data_2_15_i_7[1]_net_1 ));
    CFG3 #( .INIT(8'hF8) )  \mem_14__RNISAMI[4]  (.A(
        un1_mem_0_5_116_set_net_1), .B(un1_mem_0_5_244_rs_net_1), .C(
        \mem_14_rs[4] ), .Y(\mem_14_[4]_net_1 ));
    CFG3 #( .INIT(8'hF2) )  un1_mem_0_5_173 (.A(\mem_8_[7]_net_1 ), .B(
        N_479), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_173_i));
    CFG3 #( .INIT(8'hF2) )  un1_mem_0_5_225 (.A(\mem_8_[3]_net_1 ), .B(
        N_479), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_225_i));
    CFG1 #( .INIT(2'h1) )  un1_mem_0_5_99_set_RNO (.A(
        un1_mem_0_5_99_net_1), .Y(un1_mem_0_5_99_i));
    SLE un1_mem_0_5_236_rs (.D(VCC_net_1), .CLK(un1_mem_0_5_108_net_1), 
        .EN(VCC_net_1), .ALn(un1_mem_0_5_236_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(VCC_net_1), .Q(
        un1_mem_0_5_236_rs_net_1));
    SLE un1_mem_0_5_153_rs (.D(VCC_net_1), .CLK(un1_mem_0_5_124_net_1), 
        .EN(VCC_net_1), .ALn(un1_mem_0_5_153_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(VCC_net_1), .Q(
        un1_mem_0_5_153_rs_net_1));
    CFG4 #( .INIT(16'h7530) )  \temp_data_2_15_i_7[2]  (.A(
        \mem_12_[2]_net_1 ), .B(\mem_8_[2]_net_1 ), .C(N_479), .D(
        N_469), .Y(\temp_data_2_15_i_7[2]_net_1 ));
    CFG1 #( .INIT(2'h1) )  un1_mem_0_5_85_set_RNO (.A(
        un1_mem_0_5_85_net_1), .Y(un1_mem_0_5_85_i));
    CFG3 #( .INIT(8'hF2) )  un1_mem_0_5_130 (.A(\mem_0_[3]_net_1 ), .B(
        N_473), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_130_i));
    CFG1 #( .INIT(2'h1) )  un1_mem_0_5_28_set_RNO (.A(
        un1_mem_0_5_28_net_1), .Y(un1_mem_0_5_28_i));
    CFG4 #( .INIT(16'h0020) )  \WRITE_GEN.mem_9__2_i_a2[7]  (.A(
        CoreAPB3_0_APBmslave2_PADDR[3]), .B(
        CoreAPB3_0_APBmslave2_PADDR[2]), .C(
        CoreAPB3_0_APBmslave2_PADDR[0]), .D(
        CoreAPB3_0_APBmslave2_PADDR[1]), .Y(N_467));
    SLE un1_mem_0_5_95_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_11__1_sqmuxa), .ALn(un1_mem_0_5_95_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_mem_0_5_95_set_net_1));
    CFG2 #( .INIT(4'h8) )  mem_11__1_sqmuxa_0_a2 (.A(N_475), .B(
        wr_enable), .Y(mem_11__1_sqmuxa));
    CFG3 #( .INIT(8'hF8) )  un1_mem_0_5_54_set_RNISMNC (.A(
        un1_mem_0_5_54_set_net_1), .B(un1_mem_0_5_213_rs_net_1), .C(
        \mem_7_rs[5] ), .Y(\mem_7_[5]_net_1 ));
    SLE un1_mem_0_5_25_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_5__1_sqmuxa), .ALn(un1_mem_0_5_25_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_mem_0_5_25_set_net_1));
    CFG3 #( .INIT(8'hF8) )  un1_mem_0_5_210_rs_RNIKVRC (.A(
        un1_mem_0_5_51_set_net_1), .B(un1_mem_0_5_210_rs_net_1), .C(
        \mem_7_rs[3] ), .Y(\mem_7_[3]_net_1 ));
    CFG3 #( .INIT(8'hF8) )  un1_mem_0_5_129_rs_RNIPFDM (.A(
        un1_mem_0_5_82_set_net_1), .B(un1_mem_0_5_129_rs_net_1), .C(
        \mem_0_rs[2] ), .Y(\mem_0_[2]_net_1 ));
    CFG3 #( .INIT(8'h02) )  un1_mem_0_5_114 (.A(\mem_14_[2]_net_1 ), 
        .B(N_482), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_114_net_1));
    CFG1 #( .INIT(2'h1) )  un1_mem_0_5_103_set_RNO (.A(
        un1_mem_0_5_103_net_1), .Y(un1_mem_0_5_103_i));
    CFG3 #( .INIT(8'hF8) )  un1_mem_0_5_89_set_RNIGNAI (.A(
        un1_mem_0_5_89_set_net_1), .B(un1_mem_0_5_209_rs_net_1), .C(
        \mem_11_rs[1] ), .Y(\mem_11_[1]_net_1 ));
    CFG1 #( .INIT(2'h1) )  un1_mem_0_5_34_set_RNO (.A(
        un1_mem_0_5_34_net_1), .Y(un1_mem_0_5_34_i));
    SLE \mem_6_[2]  (.D(CoreAPB3_0_APBmslave2_PWDATA[2]), .CLK(
        FCCC_0_GL1), .EN(mem_6__1_sqmuxa), .ALn(un1_mem_0_5_192_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_6_rs[2] ));
    CFG3 #( .INIT(8'h02) )  un1_mem_0_5_68 (.A(\mem_8_[4]_net_1 ), .B(
        N_479), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_68_net_1));
    SLE un1_mem_0_5_174_rs (.D(VCC_net_1), .CLK(un1_mem_0_5_15_net_1), 
        .EN(VCC_net_1), .ALn(un1_mem_0_5_174_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(VCC_net_1), .Q(
        un1_mem_0_5_174_rs_net_1));
    CFG3 #( .INIT(8'h02) )  un1_mem_0_5_26 (.A(\mem_2_[0]_net_1 ), .B(
        N_478), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_26_net_1));
    SLE un1_mem_0_5_101_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_10__1_sqmuxa), .ALn(un1_mem_0_5_101_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_mem_0_5_101_set_net_1));
    CFG4 #( .INIT(16'h7530) )  \temp_data_2_15_i_7[7]  (.A(
        \mem_12_[7]_net_1 ), .B(\mem_8_[7]_net_1 ), .C(N_479), .D(
        N_469), .Y(\temp_data_2_15_i_7[7]_net_1 ));
    CFG3 #( .INIT(8'h02) )  un1_mem_0_5_69 (.A(\mem_8_[5]_net_1 ), .B(
        N_479), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_69_net_1));
    CFG1 #( .INIT(2'h1) )  un1_mem_0_5_126_set_RNO (.A(
        un1_mem_0_5_126_net_1), .Y(un1_mem_0_5_126_i));
    CFG3 #( .INIT(8'hF2) )  un1_mem_0_5_179 (.A(\mem_9_[2]_net_1 ), .B(
        N_467), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_179_i));
    SLE \temp_data[2]  (.D(N_10_i_0), .CLK(FCCC_0_GL1), .EN(rd_enable), 
        .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\temp_data[2]_net_1 ));
    CFG3 #( .INIT(8'hF2) )  un1_mem_0_5_177 (.A(\mem_9_[1]_net_1 ), .B(
        N_467), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_177_i));
    SLE \mem_7_[7]  (.D(CoreAPB3_0_APBmslave2_PWDATA[7]), .CLK(
        FCCC_0_GL1), .EN(mem_7__1_sqmuxa), .ALn(un1_mem_0_5_217_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_7_rs[7] ));
    CFG3 #( .INIT(8'hF8) )  un1_mem_0_5_8_set_RNI90TH (.A(
        un1_mem_0_5_8_set_net_1), .B(un1_mem_0_5_135_rs_net_1), .C(
        \mem_0_rs[7] ), .Y(\mem_0_[7]_net_1 ));
    CFG3 #( .INIT(8'hF8) )  un1_mem_0_5_104_set_RNIHBD51 (.A(
        un1_mem_0_5_104_set_net_1), .B(un1_mem_0_5_232_rs_net_1), .C(
        \mem_13_rs[0] ), .Y(\mem_13_[0]_net_1 ));
    CFG1 #( .INIT(2'h1) )  un1_mem_0_5_44_set_RNO (.A(
        un1_mem_0_5_44_net_1), .Y(un1_mem_0_5_44_i));
    SLE \mem_0_[2]  (.D(CoreAPB3_0_APBmslave2_PWDATA[2]), .CLK(
        FCCC_0_GL1), .EN(mem_0__1_sqmuxa), .ALn(un1_mem_0_5_129_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_0_rs[2] ));
    CFG3 #( .INIT(8'hF2) )  un1_mem_0_5_155 (.A(\mem_3_[3]_net_1 ), .B(
        N_470), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_155_i));
    SLE \mem_3_[6]  (.D(CoreAPB3_0_APBmslave2_PWDATA[6]), .CLK(
        FCCC_0_GL1), .EN(mem_3__1_sqmuxa), .ALn(un1_mem_0_5_159_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_3_rs[6] ));
    SLE \mem_2_[7]  (.D(CoreAPB3_0_APBmslave2_PWDATA[7]), .CLK(
        FCCC_0_GL1), .EN(mem_2__1_sqmuxa), .ALn(un1_mem_0_5_151_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_2_rs[7] ));
    SLE un1_mem_0_5_100_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_10__1_sqmuxa), .ALn(un1_mem_0_5_100_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_mem_0_5_100_set_net_1));
    SLE \mem_7_[5]  (.D(CoreAPB3_0_APBmslave2_PWDATA[5]), .CLK(
        FCCC_0_GL1), .EN(mem_7__1_sqmuxa), .ALn(un1_mem_0_5_213_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_7_rs[5] ));
    SLE un1_mem_0_5_200_rs (.D(VCC_net_1), .CLK(un1_mem_0_5_121_net_1), 
        .EN(VCC_net_1), .ALn(un1_mem_0_5_200_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(VCC_net_1), .Q(
        un1_mem_0_5_200_rs_net_1));
    CFG3 #( .INIT(8'h02) )  un1_mem_0_5_56 (.A(\mem_15_[2]_net_1 ), .B(
        N_474), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_56_net_1));
    CFG3 #( .INIT(8'hF2) )  un1_mem_0_5_183 (.A(\mem_9_[4]_net_1 ), .B(
        N_467), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_183_i));
    CFG1 #( .INIT(2'h1) )  un1_mem_0_5_22_set_RNO (.A(
        un1_mem_0_5_22_net_1), .Y(un1_mem_0_5_22_i));
    SLE \mem_2_[5]  (.D(CoreAPB3_0_APBmslave2_PWDATA[5]), .CLK(
        FCCC_0_GL1), .EN(mem_2__1_sqmuxa), .ALn(un1_mem_0_5_149_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_2_rs[5] ));
    CFG1 #( .INIT(2'h1) )  un1_mem_0_5_90_set_RNO (.A(
        un1_mem_0_5_90_net_1), .Y(un1_mem_0_5_90_i));
    SLE un1_mem_0_5_211_rs (.D(VCC_net_1), .CLK(un1_mem_0_5_90_net_1), 
        .EN(VCC_net_1), .ALn(un1_mem_0_5_211_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(VCC_net_1), .Q(
        un1_mem_0_5_211_rs_net_1));
    SLE \mem_4_[7]  (.D(CoreAPB3_0_APBmslave2_PWDATA[7]), .CLK(
        FCCC_0_GL1), .EN(mem_4__1_sqmuxa), .ALn(un1_mem_0_5_170_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_4_rs[7] ));
    CFG1 #( .INIT(2'h1) )  un1_mem_0_5_89_set_RNO (.A(
        un1_mem_0_5_89_net_1), .Y(un1_mem_0_5_89_i));
    CFG3 #( .INIT(8'h02) )  un1_mem_0_5_100 (.A(\mem_10_[7]_net_1 ), 
        .B(N_471), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_100_net_1));
    SLE un1_mem_0_5_232_rs (.D(VCC_net_1), .CLK(un1_mem_0_5_104_net_1), 
        .EN(VCC_net_1), .ALn(un1_mem_0_5_232_i), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(VCC_net_1), .Q(
        un1_mem_0_5_232_rs_net_1));
    CFG3 #( .INIT(8'hF2) )  un1_mem_0_5_193 (.A(\mem_10_[1]_net_1 ), 
        .B(N_471), .C(MSS_RESET_N_F2M_c), .Y(un1_mem_0_5_193_i));
    SLE \mem_14_[3]  (.D(CoreAPB3_0_APBmslave2_PWDATA[3]), .CLK(
        FCCC_0_GL1), .EN(mem_14__1_sqmuxa), .ALn(un1_mem_0_5_243_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_14_rs[3] ));
    
endmodule


module reg_apb_wrp(
       CoreAPB3_0_APBmslave3_PRDATA,
       CoreAPB3_0_APBmslave2_PWDATA,
       CoreAPB3_0_APBmslave2_PADDR,
       CoreAPB3_0_APBmslave3_PREADY,
       MSS_RESET_N_F2M_c,
       FCCC_0_GL1,
       CoreAPB3_0_APBmslave2_PWRITE,
       CoreAPB3_0_APBmslave3_PSELx
    );
output [7:0] CoreAPB3_0_APBmslave3_PRDATA;
input  [7:0] CoreAPB3_0_APBmslave2_PWDATA;
input  [3:0] CoreAPB3_0_APBmslave2_PADDR;
output CoreAPB3_0_APBmslave3_PREADY;
input  MSS_RESET_N_F2M_c;
input  FCCC_0_GL1;
input  CoreAPB3_0_APBmslave2_PWRITE;
input  CoreAPB3_0_APBmslave3_PSELx;

    wire GND_net_1, N_64_i_0, N_44_i_0, VCC_net_1, wr_enable_net_1, 
        N_70, N_45_i_0, rd_enable_net_1, N_76, \fsm[0]_net_1 , 
        \fsm_ns[0] , \fsm[1]_net_1 , \fsm_ns[1] ;
    
    CFG2 #( .INIT(4'h1) )  rd_enable_RNO (.A(
        CoreAPB3_0_APBmslave2_PWRITE), .B(\fsm[0]_net_1 ), .Y(N_76));
    CFG3 #( .INIT(8'h54) )  \fsm_RNIENS51[1]  (.A(\fsm[1]_net_1 ), .B(
        \fsm[0]_net_1 ), .C(CoreAPB3_0_APBmslave3_PSELx), .Y(N_45_i_0));
    SLE rd_enable (.D(N_76), .CLK(FCCC_0_GL1), .EN(N_45_i_0), .ALn(
        MSS_RESET_N_F2M_c), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(rd_enable_net_1));
    CFG2 #( .INIT(4'hE) )  PREADY_RNO (.A(CoreAPB3_0_APBmslave2_PWRITE)
        , .B(\fsm[1]_net_1 ), .Y(N_64_i_0));
    SLE PREADY (.D(N_64_i_0), .CLK(FCCC_0_GL1), .EN(N_44_i_0), .ALn(
        MSS_RESET_N_F2M_c), .ADn(GND_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(CoreAPB3_0_APBmslave3_PREADY));
    GND GND (.Y(GND_net_1));
    CFG3 #( .INIT(8'h32) )  \fsm_ns_1_0_.m2  (.A(\fsm[1]_net_1 ), .B(
        \fsm[0]_net_1 ), .C(CoreAPB3_0_APBmslave3_PSELx), .Y(
        \fsm_ns[0] ));
    CFG3 #( .INIT(8'h26) )  \fsm_ns_1_0_.m4  (.A(\fsm[1]_net_1 ), .B(
        \fsm[0]_net_1 ), .C(CoreAPB3_0_APBmslave2_PWRITE), .Y(
        \fsm_ns[1] ));
    VCC VCC (.Y(VCC_net_1));
    reg16x8 reg16x8_0 (.CoreAPB3_0_APBmslave3_PRDATA({
        CoreAPB3_0_APBmslave3_PRDATA[7], 
        CoreAPB3_0_APBmslave3_PRDATA[6], 
        CoreAPB3_0_APBmslave3_PRDATA[5], 
        CoreAPB3_0_APBmslave3_PRDATA[4], 
        CoreAPB3_0_APBmslave3_PRDATA[3], 
        CoreAPB3_0_APBmslave3_PRDATA[2], 
        CoreAPB3_0_APBmslave3_PRDATA[1], 
        CoreAPB3_0_APBmslave3_PRDATA[0]}), 
        .CoreAPB3_0_APBmslave2_PWDATA({CoreAPB3_0_APBmslave2_PWDATA[7], 
        CoreAPB3_0_APBmslave2_PWDATA[6], 
        CoreAPB3_0_APBmslave2_PWDATA[5], 
        CoreAPB3_0_APBmslave2_PWDATA[4], 
        CoreAPB3_0_APBmslave2_PWDATA[3], 
        CoreAPB3_0_APBmslave2_PWDATA[2], 
        CoreAPB3_0_APBmslave2_PWDATA[1], 
        CoreAPB3_0_APBmslave2_PWDATA[0]}), 
        .CoreAPB3_0_APBmslave2_PADDR({CoreAPB3_0_APBmslave2_PADDR[3], 
        CoreAPB3_0_APBmslave2_PADDR[2], CoreAPB3_0_APBmslave2_PADDR[1], 
        CoreAPB3_0_APBmslave2_PADDR[0]}), .MSS_RESET_N_F2M_c(
        MSS_RESET_N_F2M_c), .FCCC_0_GL1(FCCC_0_GL1), .rd_enable(
        rd_enable_net_1), .wr_enable(wr_enable_net_1));
    CFG3 #( .INIT(8'h76) )  PREADY_RNO_0 (.A(\fsm[1]_net_1 ), .B(
        \fsm[0]_net_1 ), .C(CoreAPB3_0_APBmslave3_PSELx), .Y(N_44_i_0));
    CFG2 #( .INIT(4'h2) )  wr_enable_RNO (.A(
        CoreAPB3_0_APBmslave2_PWRITE), .B(\fsm[0]_net_1 ), .Y(N_70));
    SLE \fsm[0]  (.D(\fsm_ns[0] ), .CLK(FCCC_0_GL1), .EN(VCC_net_1), 
        .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\fsm[0]_net_1 ));
    SLE wr_enable (.D(N_70), .CLK(FCCC_0_GL1), .EN(N_45_i_0), .ALn(
        MSS_RESET_N_F2M_c), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(wr_enable_net_1));
    SLE \fsm[1]  (.D(\fsm_ns[1] ), .CLK(FCCC_0_GL1), .EN(VCC_net_1), 
        .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\fsm[1]_net_1 ));
    
endmodule


module FIC_MSS(
       CoreAPB3_0_APBmslave2_PADDR,
       FIC_MSS_0_FIC_0_APB_MASTER_PADDR,
       CoreAPB3_0_APBmslave2_PWDATA,
       FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_0,
       FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_1,
       FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_4,
       FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_5,
       FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_6,
       FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_7,
       FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_8,
       FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_9,
       FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_10,
       FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_11,
       FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_12,
       FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_13,
       FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_14,
       FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_15,
       FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_16,
       FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_17,
       FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_18,
       FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_19,
       FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_20,
       FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_21,
       FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_22,
       FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_23,
       FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_24,
       FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_25,
       FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_26,
       FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_27,
       FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_28,
       MMUART_0_TXD,
       MMUART_0_RXD,
       CoreAPB3_0_APBmslave2_PENABLE,
       FIC_MSS_0_FIC_0_APB_MASTER_PSELx,
       CoreAPB3_0_APBmslave2_PWRITE,
       CoreAPB3_N_8_i_0,
       CoreAPB3_N_8_2_i_0,
       CoreAPB3_N_8_3_i_0,
       CoreAPB3_N_8_1_i_0,
       CoreAPB3_N_8_0_i_0,
       PREADY_0_iv_i_0,
       FCCC_0_LOCK,
       MSS_RESET_N_F2M_c,
       FCCC_0_GL1
    );
output [8:0] CoreAPB3_0_APBmslave2_PADDR;
output [31:28] FIC_MSS_0_FIC_0_APB_MASTER_PADDR;
output [31:0] CoreAPB3_0_APBmslave2_PWDATA;
input  FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_0;
input  FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_1;
input  FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_4;
input  FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_5;
input  FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_6;
input  FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_7;
input  FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_8;
input  FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_9;
input  FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_10;
input  FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_11;
input  FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_12;
input  FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_13;
input  FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_14;
input  FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_15;
input  FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_16;
input  FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_17;
input  FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_18;
input  FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_19;
input  FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_20;
input  FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_21;
input  FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_22;
input  FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_23;
input  FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_24;
input  FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_25;
input  FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_26;
input  FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_27;
input  FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_28;
output MMUART_0_TXD;
input  MMUART_0_RXD;
output CoreAPB3_0_APBmslave2_PENABLE;
output FIC_MSS_0_FIC_0_APB_MASTER_PSELx;
output CoreAPB3_0_APBmslave2_PWRITE;
input  CoreAPB3_N_8_i_0;
input  CoreAPB3_N_8_2_i_0;
input  CoreAPB3_N_8_3_i_0;
input  CoreAPB3_N_8_1_i_0;
input  CoreAPB3_N_8_0_i_0;
input  PREADY_0_iv_i_0;
input  FCCC_0_LOCK;
input  MSS_RESET_N_F2M_c;
input  FCCC_0_GL1;

    wire MSS_ADLIB_INST_MMUART0_TXD_USBC_DIR_MGPIO27B_OUT, 
        MSS_ADLIB_INST_MMUART0_TXD_USBC_DIR_MGPIO27B_OE, 
        MMUART_0_RXD_PAD_Y, VCC_net_1, GND_net_1;
    
    INBUF MMUART_0_RXD_PAD (.PAD(MMUART_0_RXD), .Y(MMUART_0_RXD_PAD_Y));
    VCC VCC (.Y(VCC_net_1));
    MSS_010 #( .INIT(1438'h00000000003612000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000F00000000F000000000000000000000000000000007FFFFFFFB000001007C33C000000006092C0104003FFFFE400000000000010000000000001C000001FEDFDC010842108421000001FE34001FF8000000400000000020091007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF)
        , .ACT_UBITS(56'hFFFFFFFFFFFFFF), .MEMORYFILE("ENVM_init.mem")
        , .RTC_MAIN_XTL_FREQ(0.0), .RTC_MAIN_XTL_MODE("") )  
        MSS_ADLIB_INST (.CAN_RXBUS_MGPIO3A_H2F_A(), 
        .CAN_RXBUS_MGPIO3A_H2F_B(), .CAN_TX_EBL_MGPIO4A_H2F_A(), 
        .CAN_TX_EBL_MGPIO4A_H2F_B(), .CAN_TXBUS_MGPIO2A_H2F_A(), 
        .CAN_TXBUS_MGPIO2A_H2F_B(), .CLK_CONFIG_APB(), .COMMS_INT(), 
        .CONFIG_PRESET_N(), .EDAC_ERROR({nc0, nc1, nc2, nc3, nc4, nc5, 
        nc6, nc7}), .F_FM0_RDATA({nc8, nc9, nc10, nc11, nc12, nc13, 
        nc14, nc15, nc16, nc17, nc18, nc19, nc20, nc21, nc22, nc23, 
        nc24, nc25, nc26, nc27, nc28, nc29, nc30, nc31, nc32, nc33, 
        nc34, nc35, nc36, nc37, nc38, nc39}), .F_FM0_READYOUT(), 
        .F_FM0_RESP(), .F_HM0_ADDR({
        FIC_MSS_0_FIC_0_APB_MASTER_PADDR[31], 
        FIC_MSS_0_FIC_0_APB_MASTER_PADDR[30], 
        FIC_MSS_0_FIC_0_APB_MASTER_PADDR[29], 
        FIC_MSS_0_FIC_0_APB_MASTER_PADDR[28], nc40, nc41, nc42, nc43, 
        nc44, nc45, nc46, nc47, nc48, nc49, nc50, nc51, nc52, nc53, 
        nc54, nc55, nc56, nc57, nc58, CoreAPB3_0_APBmslave2_PADDR[8], 
        CoreAPB3_0_APBmslave2_PADDR[7], CoreAPB3_0_APBmslave2_PADDR[6], 
        CoreAPB3_0_APBmslave2_PADDR[5], CoreAPB3_0_APBmslave2_PADDR[4], 
        CoreAPB3_0_APBmslave2_PADDR[3], CoreAPB3_0_APBmslave2_PADDR[2], 
        CoreAPB3_0_APBmslave2_PADDR[1], CoreAPB3_0_APBmslave2_PADDR[0]})
        , .F_HM0_ENABLE(CoreAPB3_0_APBmslave2_PENABLE), .F_HM0_SEL(
        FIC_MSS_0_FIC_0_APB_MASTER_PSELx), .F_HM0_SIZE({nc59, nc60}), 
        .F_HM0_TRANS1(), .F_HM0_WDATA({
        CoreAPB3_0_APBmslave2_PWDATA[31], 
        CoreAPB3_0_APBmslave2_PWDATA[30], 
        CoreAPB3_0_APBmslave2_PWDATA[29], 
        CoreAPB3_0_APBmslave2_PWDATA[28], 
        CoreAPB3_0_APBmslave2_PWDATA[27], 
        CoreAPB3_0_APBmslave2_PWDATA[26], 
        CoreAPB3_0_APBmslave2_PWDATA[25], 
        CoreAPB3_0_APBmslave2_PWDATA[24], 
        CoreAPB3_0_APBmslave2_PWDATA[23], 
        CoreAPB3_0_APBmslave2_PWDATA[22], 
        CoreAPB3_0_APBmslave2_PWDATA[21], 
        CoreAPB3_0_APBmslave2_PWDATA[20], 
        CoreAPB3_0_APBmslave2_PWDATA[19], 
        CoreAPB3_0_APBmslave2_PWDATA[18], 
        CoreAPB3_0_APBmslave2_PWDATA[17], 
        CoreAPB3_0_APBmslave2_PWDATA[16], 
        CoreAPB3_0_APBmslave2_PWDATA[15], 
        CoreAPB3_0_APBmslave2_PWDATA[14], 
        CoreAPB3_0_APBmslave2_PWDATA[13], 
        CoreAPB3_0_APBmslave2_PWDATA[12], 
        CoreAPB3_0_APBmslave2_PWDATA[11], 
        CoreAPB3_0_APBmslave2_PWDATA[10], 
        CoreAPB3_0_APBmslave2_PWDATA[9], 
        CoreAPB3_0_APBmslave2_PWDATA[8], 
        CoreAPB3_0_APBmslave2_PWDATA[7], 
        CoreAPB3_0_APBmslave2_PWDATA[6], 
        CoreAPB3_0_APBmslave2_PWDATA[5], 
        CoreAPB3_0_APBmslave2_PWDATA[4], 
        CoreAPB3_0_APBmslave2_PWDATA[3], 
        CoreAPB3_0_APBmslave2_PWDATA[2], 
        CoreAPB3_0_APBmslave2_PWDATA[1], 
        CoreAPB3_0_APBmslave2_PWDATA[0]}), .F_HM0_WRITE(
        CoreAPB3_0_APBmslave2_PWRITE), .FAB_CHRGVBUS(), 
        .FAB_DISCHRGVBUS(), .FAB_DMPULLDOWN(), .FAB_DPPULLDOWN(), 
        .FAB_DRVVBUS(), .FAB_IDPULLUP(), .FAB_OPMODE({nc61, nc62}), 
        .FAB_SUSPENDM(), .FAB_TERMSEL(), .FAB_TXVALID(), .FAB_VCONTROL({
        nc63, nc64, nc65, nc66}), .FAB_VCONTROLLOADM(), .FAB_XCVRSEL({
        nc67, nc68}), .FAB_XDATAOUT({nc69, nc70, nc71, nc72, nc73, 
        nc74, nc75, nc76}), .FACC_GLMUX_SEL(), .FIC32_0_MASTER({nc77, 
        nc78}), .FIC32_1_MASTER({nc79, nc80}), .FPGA_RESET_N(), 
        .GTX_CLK(), .H2F_INTERRUPT({nc81, nc82, nc83, nc84, nc85, nc86, 
        nc87, nc88, nc89, nc90, nc91, nc92, nc93, nc94, nc95, nc96}), 
        .H2F_NMI(), .H2FCALIB(), .I2C0_SCL_MGPIO31B_H2F_A(), 
        .I2C0_SCL_MGPIO31B_H2F_B(), .I2C0_SDA_MGPIO30B_H2F_A(), 
        .I2C0_SDA_MGPIO30B_H2F_B(), .I2C1_SCL_MGPIO1A_H2F_A(), 
        .I2C1_SCL_MGPIO1A_H2F_B(), .I2C1_SDA_MGPIO0A_H2F_A(), 
        .I2C1_SDA_MGPIO0A_H2F_B(), .MDCF(), .MDOENF(), .MDOF(), 
        .MMUART0_CTS_MGPIO19B_H2F_A(), .MMUART0_CTS_MGPIO19B_H2F_B(), 
        .MMUART0_DCD_MGPIO22B_H2F_A(), .MMUART0_DCD_MGPIO22B_H2F_B(), 
        .MMUART0_DSR_MGPIO20B_H2F_A(), .MMUART0_DSR_MGPIO20B_H2F_B(), 
        .MMUART0_DTR_MGPIO18B_H2F_A(), .MMUART0_DTR_MGPIO18B_H2F_B(), 
        .MMUART0_RI_MGPIO21B_H2F_A(), .MMUART0_RI_MGPIO21B_H2F_B(), 
        .MMUART0_RTS_MGPIO17B_H2F_A(), .MMUART0_RTS_MGPIO17B_H2F_B(), 
        .MMUART0_RXD_MGPIO28B_H2F_A(), .MMUART0_RXD_MGPIO28B_H2F_B(), 
        .MMUART0_SCK_MGPIO29B_H2F_A(), .MMUART0_SCK_MGPIO29B_H2F_B(), 
        .MMUART0_TXD_MGPIO27B_H2F_A(), .MMUART0_TXD_MGPIO27B_H2F_B(), 
        .MMUART1_DTR_MGPIO12B_H2F_A(), .MMUART1_RTS_MGPIO11B_H2F_A(), 
        .MMUART1_RTS_MGPIO11B_H2F_B(), .MMUART1_RXD_MGPIO26B_H2F_A(), 
        .MMUART1_RXD_MGPIO26B_H2F_B(), .MMUART1_SCK_MGPIO25B_H2F_A(), 
        .MMUART1_SCK_MGPIO25B_H2F_B(), .MMUART1_TXD_MGPIO24B_H2F_A(), 
        .MMUART1_TXD_MGPIO24B_H2F_B(), .MPLL_LOCK(), 
        .PER2_FABRIC_PADDR({nc97, nc98, nc99, nc100, nc101, nc102, 
        nc103, nc104, nc105, nc106, nc107, nc108, nc109, nc110}), 
        .PER2_FABRIC_PENABLE(), .PER2_FABRIC_PSEL(), 
        .PER2_FABRIC_PWDATA({nc111, nc112, nc113, nc114, nc115, nc116, 
        nc117, nc118, nc119, nc120, nc121, nc122, nc123, nc124, nc125, 
        nc126, nc127, nc128, nc129, nc130, nc131, nc132, nc133, nc134, 
        nc135, nc136, nc137, nc138, nc139, nc140, nc141, nc142}), 
        .PER2_FABRIC_PWRITE(), .RTC_MATCH(), .SLEEPDEEP(), 
        .SLEEPHOLDACK(), .SLEEPING(), .SMBALERT_NO0(), .SMBALERT_NO1(), 
        .SMBSUS_NO0(), .SMBSUS_NO1(), .SPI0_CLK_OUT(), 
        .SPI0_SDI_MGPIO5A_H2F_A(), .SPI0_SDI_MGPIO5A_H2F_B(), 
        .SPI0_SDO_MGPIO6A_H2F_A(), .SPI0_SDO_MGPIO6A_H2F_B(), 
        .SPI0_SS0_MGPIO7A_H2F_A(), .SPI0_SS0_MGPIO7A_H2F_B(), 
        .SPI0_SS1_MGPIO8A_H2F_A(), .SPI0_SS1_MGPIO8A_H2F_B(), 
        .SPI0_SS2_MGPIO9A_H2F_A(), .SPI0_SS2_MGPIO9A_H2F_B(), 
        .SPI0_SS3_MGPIO10A_H2F_A(), .SPI0_SS3_MGPIO10A_H2F_B(), 
        .SPI0_SS4_MGPIO19A_H2F_A(), .SPI0_SS5_MGPIO20A_H2F_A(), 
        .SPI0_SS6_MGPIO21A_H2F_A(), .SPI0_SS7_MGPIO22A_H2F_A(), 
        .SPI1_CLK_OUT(), .SPI1_SDI_MGPIO11A_H2F_A(), 
        .SPI1_SDI_MGPIO11A_H2F_B(), .SPI1_SDO_MGPIO12A_H2F_A(), 
        .SPI1_SDO_MGPIO12A_H2F_B(), .SPI1_SS0_MGPIO13A_H2F_A(), 
        .SPI1_SS0_MGPIO13A_H2F_B(), .SPI1_SS1_MGPIO14A_H2F_A(), 
        .SPI1_SS1_MGPIO14A_H2F_B(), .SPI1_SS2_MGPIO15A_H2F_A(), 
        .SPI1_SS2_MGPIO15A_H2F_B(), .SPI1_SS3_MGPIO16A_H2F_A(), 
        .SPI1_SS3_MGPIO16A_H2F_B(), .SPI1_SS4_MGPIO17A_H2F_A(), 
        .SPI1_SS5_MGPIO18A_H2F_A(), .SPI1_SS6_MGPIO23A_H2F_A(), 
        .SPI1_SS7_MGPIO24A_H2F_A(), .TCGF({nc143, nc144, nc145, nc146, 
        nc147, nc148, nc149, nc150, nc151, nc152}), .TRACECLK(), 
        .TRACEDATA({nc153, nc154, nc155, nc156}), .TX_CLK(), .TX_ENF(), 
        .TX_ERRF(), .TXCTL_EN_RIF(), .TXD_RIF({nc157, nc158, nc159, 
        nc160}), .TXDF({nc161, nc162, nc163, nc164, nc165, nc166, 
        nc167, nc168}), .TXEV(), .WDOGTIMEOUT(), .F_ARREADY_HREADYOUT1(
        ), .F_AWREADY_HREADYOUT0(), .F_BID({nc169, nc170, nc171, nc172})
        , .F_BRESP_HRESP0({nc173, nc174}), .F_BVALID(), 
        .F_RDATA_HRDATA01({nc175, nc176, nc177, nc178, nc179, nc180, 
        nc181, nc182, nc183, nc184, nc185, nc186, nc187, nc188, nc189, 
        nc190, nc191, nc192, nc193, nc194, nc195, nc196, nc197, nc198, 
        nc199, nc200, nc201, nc202, nc203, nc204, nc205, nc206, nc207, 
        nc208, nc209, nc210, nc211, nc212, nc213, nc214, nc215, nc216, 
        nc217, nc218, nc219, nc220, nc221, nc222, nc223, nc224, nc225, 
        nc226, nc227, nc228, nc229, nc230, nc231, nc232, nc233, nc234, 
        nc235, nc236, nc237, nc238}), .F_RID({nc239, nc240, nc241, 
        nc242}), .F_RLAST(), .F_RRESP_HRESP1({nc243, nc244}), 
        .F_RVALID(), .F_WREADY(), .MDDR_FABRIC_PRDATA({nc245, nc246, 
        nc247, nc248, nc249, nc250, nc251, nc252, nc253, nc254, nc255, 
        nc256, nc257, nc258, nc259, nc260}), .MDDR_FABRIC_PREADY(), 
        .MDDR_FABRIC_PSLVERR(), .CAN_RXBUS_F2H_SCP(VCC_net_1), 
        .CAN_TX_EBL_F2H_SCP(VCC_net_1), .CAN_TXBUS_F2H_SCP(VCC_net_1), 
        .COLF(VCC_net_1), .CRSF(VCC_net_1), .F2_DMAREADY({VCC_net_1, 
        VCC_net_1}), .F2H_INTERRUPT({GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1}), .F2HCALIB(VCC_net_1), 
        .F_DMAREADY({VCC_net_1, VCC_net_1}), .F_FM0_ADDR({GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1}), .F_FM0_ENABLE(GND_net_1), .F_FM0_MASTLOCK(
        GND_net_1), .F_FM0_READY(VCC_net_1), .F_FM0_SEL(GND_net_1), 
        .F_FM0_SIZE({GND_net_1, GND_net_1}), .F_FM0_TRANS1(GND_net_1), 
        .F_FM0_WDATA({GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1}), .F_FM0_WRITE(GND_net_1), 
        .F_HM0_RDATA({FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_28, 
        FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_27, 
        FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_26, 
        FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_25, 
        FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_24, 
        FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_23, 
        FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_22, 
        FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_21, 
        FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_20, 
        FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_19, 
        FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_18, 
        FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_17, 
        FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_16, 
        FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_15, 
        FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_14, 
        FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_13, 
        FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_12, 
        FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_11, 
        FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_10, 
        FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_9, 
        FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_8, 
        FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_7, 
        FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_6, 
        FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_5, 
        FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_4, CoreAPB3_N_8_0_i_0, 
        CoreAPB3_N_8_1_i_0, FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_1, 
        FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_0, CoreAPB3_N_8_3_i_0, 
        CoreAPB3_N_8_2_i_0, CoreAPB3_N_8_i_0}), .F_HM0_READY(
        PREADY_0_iv_i_0), .F_HM0_RESP(GND_net_1), .FAB_AVALID(
        VCC_net_1), .FAB_HOSTDISCON(VCC_net_1), .FAB_IDDIG(VCC_net_1), 
        .FAB_LINESTATE({VCC_net_1, VCC_net_1}), .FAB_M3_RESET_N(
        VCC_net_1), .FAB_PLL_LOCK(FCCC_0_LOCK), .FAB_RXACTIVE(
        VCC_net_1), .FAB_RXERROR(VCC_net_1), .FAB_RXVALID(VCC_net_1), 
        .FAB_RXVALIDH(GND_net_1), .FAB_SESSEND(VCC_net_1), 
        .FAB_TXREADY(VCC_net_1), .FAB_VBUSVALID(VCC_net_1), 
        .FAB_VSTATUS({VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1}), .FAB_XDATAIN({
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1}), .GTX_CLKPF(VCC_net_1), 
        .I2C0_BCLK(VCC_net_1), .I2C0_SCL_F2H_SCP(VCC_net_1), 
        .I2C0_SDA_F2H_SCP(VCC_net_1), .I2C1_BCLK(VCC_net_1), 
        .I2C1_SCL_F2H_SCP(VCC_net_1), .I2C1_SDA_F2H_SCP(VCC_net_1), 
        .MDIF(VCC_net_1), .MGPIO0A_F2H_GPIN(VCC_net_1), 
        .MGPIO10A_F2H_GPIN(VCC_net_1), .MGPIO11A_F2H_GPIN(VCC_net_1), 
        .MGPIO11B_F2H_GPIN(VCC_net_1), .MGPIO12A_F2H_GPIN(VCC_net_1), 
        .MGPIO13A_F2H_GPIN(VCC_net_1), .MGPIO14A_F2H_GPIN(VCC_net_1), 
        .MGPIO15A_F2H_GPIN(VCC_net_1), .MGPIO16A_F2H_GPIN(VCC_net_1), 
        .MGPIO17B_F2H_GPIN(VCC_net_1), .MGPIO18B_F2H_GPIN(VCC_net_1), 
        .MGPIO19B_F2H_GPIN(VCC_net_1), .MGPIO1A_F2H_GPIN(VCC_net_1), 
        .MGPIO20B_F2H_GPIN(VCC_net_1), .MGPIO21B_F2H_GPIN(VCC_net_1), 
        .MGPIO22B_F2H_GPIN(VCC_net_1), .MGPIO24B_F2H_GPIN(VCC_net_1), 
        .MGPIO25B_F2H_GPIN(VCC_net_1), .MGPIO26B_F2H_GPIN(VCC_net_1), 
        .MGPIO27B_F2H_GPIN(VCC_net_1), .MGPIO28B_F2H_GPIN(VCC_net_1), 
        .MGPIO29B_F2H_GPIN(VCC_net_1), .MGPIO2A_F2H_GPIN(VCC_net_1), 
        .MGPIO30B_F2H_GPIN(VCC_net_1), .MGPIO31B_F2H_GPIN(VCC_net_1), 
        .MGPIO3A_F2H_GPIN(VCC_net_1), .MGPIO4A_F2H_GPIN(VCC_net_1), 
        .MGPIO5A_F2H_GPIN(VCC_net_1), .MGPIO6A_F2H_GPIN(VCC_net_1), 
        .MGPIO7A_F2H_GPIN(VCC_net_1), .MGPIO8A_F2H_GPIN(VCC_net_1), 
        .MGPIO9A_F2H_GPIN(VCC_net_1), .MMUART0_CTS_F2H_SCP(VCC_net_1), 
        .MMUART0_DCD_F2H_SCP(VCC_net_1), .MMUART0_DSR_F2H_SCP(
        VCC_net_1), .MMUART0_DTR_F2H_SCP(VCC_net_1), 
        .MMUART0_RI_F2H_SCP(VCC_net_1), .MMUART0_RTS_F2H_SCP(VCC_net_1)
        , .MMUART0_RXD_F2H_SCP(VCC_net_1), .MMUART0_SCK_F2H_SCP(
        VCC_net_1), .MMUART0_TXD_F2H_SCP(VCC_net_1), 
        .MMUART1_CTS_F2H_SCP(VCC_net_1), .MMUART1_DCD_F2H_SCP(
        VCC_net_1), .MMUART1_DSR_F2H_SCP(VCC_net_1), 
        .MMUART1_RI_F2H_SCP(VCC_net_1), .MMUART1_RTS_F2H_SCP(VCC_net_1)
        , .MMUART1_RXD_F2H_SCP(VCC_net_1), .MMUART1_SCK_F2H_SCP(
        VCC_net_1), .MMUART1_TXD_F2H_SCP(VCC_net_1), 
        .PER2_FABRIC_PRDATA({VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1}), 
        .PER2_FABRIC_PREADY(VCC_net_1), .PER2_FABRIC_PSLVERR(VCC_net_1)
        , .RCGF({VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1}), 
        .RX_CLKPF(VCC_net_1), .RX_DVF(VCC_net_1), .RX_ERRF(VCC_net_1), 
        .RX_EV(VCC_net_1), .RXDF({VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1}), 
        .SLEEPHOLDREQ(GND_net_1), .SMBALERT_NI0(VCC_net_1), 
        .SMBALERT_NI1(VCC_net_1), .SMBSUS_NI0(VCC_net_1), .SMBSUS_NI1(
        VCC_net_1), .SPI0_CLK_IN(VCC_net_1), .SPI0_SDI_F2H_SCP(
        VCC_net_1), .SPI0_SDO_F2H_SCP(VCC_net_1), .SPI0_SS0_F2H_SCP(
        VCC_net_1), .SPI0_SS1_F2H_SCP(VCC_net_1), .SPI0_SS2_F2H_SCP(
        VCC_net_1), .SPI0_SS3_F2H_SCP(VCC_net_1), .SPI1_CLK_IN(
        VCC_net_1), .SPI1_SDI_F2H_SCP(VCC_net_1), .SPI1_SDO_F2H_SCP(
        VCC_net_1), .SPI1_SS0_F2H_SCP(VCC_net_1), .SPI1_SS1_F2H_SCP(
        VCC_net_1), .SPI1_SS2_F2H_SCP(VCC_net_1), .SPI1_SS3_F2H_SCP(
        VCC_net_1), .TX_CLKPF(VCC_net_1), .USER_MSS_GPIO_RESET_N(
        VCC_net_1), .USER_MSS_RESET_N(MSS_RESET_N_F2M_c), .XCLK_FAB(
        VCC_net_1), .CLK_BASE(FCCC_0_GL1), .CLK_MDDR_APB(VCC_net_1), 
        .F_ARADDR_HADDR1({VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1}), .F_ARBURST_HTRANS1({
        GND_net_1, GND_net_1}), .F_ARID_HSEL1({GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1}), .F_ARLEN_HBURST1({GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1}), .F_ARLOCK_HMASTLOCK1({GND_net_1, 
        GND_net_1}), .F_ARSIZE_HSIZE1({GND_net_1, GND_net_1}), 
        .F_ARVALID_HWRITE1(GND_net_1), .F_AWADDR_HADDR0({VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1}), .F_AWBURST_HTRANS0({GND_net_1, GND_net_1}), 
        .F_AWID_HSEL0({GND_net_1, GND_net_1, GND_net_1, GND_net_1}), 
        .F_AWLEN_HBURST0({GND_net_1, GND_net_1, GND_net_1, GND_net_1}), 
        .F_AWLOCK_HMASTLOCK0({GND_net_1, GND_net_1}), .F_AWSIZE_HSIZE0({
        GND_net_1, GND_net_1}), .F_AWVALID_HWRITE0(GND_net_1), 
        .F_BREADY(GND_net_1), .F_RMW_AXI(GND_net_1), .F_RREADY(
        GND_net_1), .F_WDATA_HWDATA01({VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1}), .F_WID_HREADY01({GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1}), .F_WLAST(GND_net_1), .F_WSTRB({GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1}), .F_WVALID(GND_net_1), 
        .FPGA_MDDR_ARESET_N(VCC_net_1), .MDDR_FABRIC_PADDR({VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1}), .MDDR_FABRIC_PENABLE(
        VCC_net_1), .MDDR_FABRIC_PSEL(VCC_net_1), .MDDR_FABRIC_PWDATA({
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1}), .MDDR_FABRIC_PWRITE(VCC_net_1), .PRESET_N(
        GND_net_1), .CAN_RXBUS_USBA_DATA1_MGPIO3A_IN(GND_net_1), 
        .CAN_TX_EBL_USBA_DATA2_MGPIO4A_IN(GND_net_1), 
        .CAN_TXBUS_USBA_DATA0_MGPIO2A_IN(GND_net_1), .DM_IN({GND_net_1, 
        GND_net_1, GND_net_1}), .DRAM_DQ_IN({GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1}), .DRAM_DQS_IN({GND_net_1, GND_net_1, GND_net_1}), 
        .DRAM_FIFO_WE_IN({GND_net_1, GND_net_1}), 
        .I2C0_SCL_USBC_DATA1_MGPIO31B_IN(GND_net_1), 
        .I2C0_SDA_USBC_DATA0_MGPIO30B_IN(GND_net_1), 
        .I2C1_SCL_USBA_DATA4_MGPIO1A_IN(GND_net_1), 
        .I2C1_SDA_USBA_DATA3_MGPIO0A_IN(GND_net_1), 
        .MMUART0_CTS_USBC_DATA7_MGPIO19B_IN(GND_net_1), 
        .MMUART0_DCD_MGPIO22B_IN(GND_net_1), .MMUART0_DSR_MGPIO20B_IN(
        GND_net_1), .MMUART0_DTR_USBC_DATA6_MGPIO18B_IN(GND_net_1), 
        .MMUART0_RI_MGPIO21B_IN(GND_net_1), 
        .MMUART0_RTS_USBC_DATA5_MGPIO17B_IN(GND_net_1), 
        .MMUART0_RXD_USBC_STP_MGPIO28B_IN(MMUART_0_RXD_PAD_Y), 
        .MMUART0_SCK_USBC_NXT_MGPIO29B_IN(GND_net_1), 
        .MMUART0_TXD_USBC_DIR_MGPIO27B_IN(GND_net_1), 
        .MMUART1_RXD_USBC_DATA3_MGPIO26B_IN(GND_net_1), 
        .MMUART1_SCK_USBC_DATA4_MGPIO25B_IN(GND_net_1), 
        .MMUART1_TXD_USBC_DATA2_MGPIO24B_IN(GND_net_1), 
        .RGMII_GTX_CLK_RMII_CLK_USBB_XCLK_IN(GND_net_1), 
        .RGMII_MDC_RMII_MDC_IN(GND_net_1), 
        .RGMII_MDIO_RMII_MDIO_USBB_DATA7_IN(GND_net_1), 
        .RGMII_RX_CLK_IN(GND_net_1), 
        .RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_IN(GND_net_1), 
        .RGMII_RXD0_RMII_RXD0_USBB_DATA0_IN(GND_net_1), 
        .RGMII_RXD1_RMII_RXD1_USBB_DATA1_IN(GND_net_1), 
        .RGMII_RXD2_RMII_RX_ER_USBB_DATA3_IN(GND_net_1), 
        .RGMII_RXD3_USBB_DATA4_IN(GND_net_1), .RGMII_TX_CLK_IN(
        GND_net_1), .RGMII_TX_CTL_RMII_TX_EN_USBB_NXT_IN(GND_net_1), 
        .RGMII_TXD0_RMII_TXD0_USBB_DIR_IN(GND_net_1), 
        .RGMII_TXD1_RMII_TXD1_USBB_STP_IN(GND_net_1), 
        .RGMII_TXD2_USBB_DATA5_IN(GND_net_1), 
        .RGMII_TXD3_USBB_DATA6_IN(GND_net_1), .SPI0_SCK_USBA_XCLK_IN(
        GND_net_1), .SPI0_SDI_USBA_DIR_MGPIO5A_IN(GND_net_1), 
        .SPI0_SDO_USBA_STP_MGPIO6A_IN(GND_net_1), 
        .SPI0_SS0_USBA_NXT_MGPIO7A_IN(GND_net_1), 
        .SPI0_SS1_USBA_DATA5_MGPIO8A_IN(GND_net_1), 
        .SPI0_SS2_USBA_DATA6_MGPIO9A_IN(GND_net_1), 
        .SPI0_SS3_USBA_DATA7_MGPIO10A_IN(GND_net_1), .SPI1_SCK_IN(
        GND_net_1), .SPI1_SDI_MGPIO11A_IN(GND_net_1), 
        .SPI1_SDO_MGPIO12A_IN(GND_net_1), .SPI1_SS0_MGPIO13A_IN(
        GND_net_1), .SPI1_SS1_MGPIO14A_IN(GND_net_1), 
        .SPI1_SS2_MGPIO15A_IN(GND_net_1), .SPI1_SS3_MGPIO16A_IN(
        GND_net_1), .SPI1_SS4_MGPIO17A_IN(GND_net_1), 
        .SPI1_SS5_MGPIO18A_IN(GND_net_1), .SPI1_SS6_MGPIO23A_IN(
        GND_net_1), .SPI1_SS7_MGPIO24A_IN(GND_net_1), .USBC_XCLK_IN(
        GND_net_1), .CAN_RXBUS_USBA_DATA1_MGPIO3A_OUT(), 
        .CAN_TX_EBL_USBA_DATA2_MGPIO4A_OUT(), 
        .CAN_TXBUS_USBA_DATA0_MGPIO2A_OUT(), .DRAM_ADDR({nc261, nc262, 
        nc263, nc264, nc265, nc266, nc267, nc268, nc269, nc270, nc271, 
        nc272, nc273, nc274, nc275, nc276}), .DRAM_BA({nc277, nc278, 
        nc279}), .DRAM_CASN(), .DRAM_CKE(), .DRAM_CLK(), .DRAM_CSN(), 
        .DRAM_DM_RDQS_OUT({nc280, nc281, nc282}), .DRAM_DQ_OUT({nc283, 
        nc284, nc285, nc286, nc287, nc288, nc289, nc290, nc291, nc292, 
        nc293, nc294, nc295, nc296, nc297, nc298, nc299, nc300}), 
        .DRAM_DQS_OUT({nc301, nc302, nc303}), .DRAM_FIFO_WE_OUT({nc304, 
        nc305}), .DRAM_ODT(), .DRAM_RASN(), .DRAM_RSTN(), .DRAM_WEN(), 
        .I2C0_SCL_USBC_DATA1_MGPIO31B_OUT(), 
        .I2C0_SDA_USBC_DATA0_MGPIO30B_OUT(), 
        .I2C1_SCL_USBA_DATA4_MGPIO1A_OUT(), 
        .I2C1_SDA_USBA_DATA3_MGPIO0A_OUT(), 
        .MMUART0_CTS_USBC_DATA7_MGPIO19B_OUT(), 
        .MMUART0_DCD_MGPIO22B_OUT(), .MMUART0_DSR_MGPIO20B_OUT(), 
        .MMUART0_DTR_USBC_DATA6_MGPIO18B_OUT(), 
        .MMUART0_RI_MGPIO21B_OUT(), 
        .MMUART0_RTS_USBC_DATA5_MGPIO17B_OUT(), 
        .MMUART0_RXD_USBC_STP_MGPIO28B_OUT(), 
        .MMUART0_SCK_USBC_NXT_MGPIO29B_OUT(), 
        .MMUART0_TXD_USBC_DIR_MGPIO27B_OUT(
        MSS_ADLIB_INST_MMUART0_TXD_USBC_DIR_MGPIO27B_OUT), 
        .MMUART1_RXD_USBC_DATA3_MGPIO26B_OUT(), 
        .MMUART1_SCK_USBC_DATA4_MGPIO25B_OUT(), 
        .MMUART1_TXD_USBC_DATA2_MGPIO24B_OUT(), 
        .RGMII_GTX_CLK_RMII_CLK_USBB_XCLK_OUT(), 
        .RGMII_MDC_RMII_MDC_OUT(), 
        .RGMII_MDIO_RMII_MDIO_USBB_DATA7_OUT(), .RGMII_RX_CLK_OUT(), 
        .RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_OUT(), 
        .RGMII_RXD0_RMII_RXD0_USBB_DATA0_OUT(), 
        .RGMII_RXD1_RMII_RXD1_USBB_DATA1_OUT(), 
        .RGMII_RXD2_RMII_RX_ER_USBB_DATA3_OUT(), 
        .RGMII_RXD3_USBB_DATA4_OUT(), .RGMII_TX_CLK_OUT(), 
        .RGMII_TX_CTL_RMII_TX_EN_USBB_NXT_OUT(), 
        .RGMII_TXD0_RMII_TXD0_USBB_DIR_OUT(), 
        .RGMII_TXD1_RMII_TXD1_USBB_STP_OUT(), 
        .RGMII_TXD2_USBB_DATA5_OUT(), .RGMII_TXD3_USBB_DATA6_OUT(), 
        .SPI0_SCK_USBA_XCLK_OUT(), .SPI0_SDI_USBA_DIR_MGPIO5A_OUT(), 
        .SPI0_SDO_USBA_STP_MGPIO6A_OUT(), 
        .SPI0_SS0_USBA_NXT_MGPIO7A_OUT(), 
        .SPI0_SS1_USBA_DATA5_MGPIO8A_OUT(), 
        .SPI0_SS2_USBA_DATA6_MGPIO9A_OUT(), 
        .SPI0_SS3_USBA_DATA7_MGPIO10A_OUT(), .SPI1_SCK_OUT(), 
        .SPI1_SDI_MGPIO11A_OUT(), .SPI1_SDO_MGPIO12A_OUT(), 
        .SPI1_SS0_MGPIO13A_OUT(), .SPI1_SS1_MGPIO14A_OUT(), 
        .SPI1_SS2_MGPIO15A_OUT(), .SPI1_SS3_MGPIO16A_OUT(), 
        .SPI1_SS4_MGPIO17A_OUT(), .SPI1_SS5_MGPIO18A_OUT(), 
        .SPI1_SS6_MGPIO23A_OUT(), .SPI1_SS7_MGPIO24A_OUT(), 
        .USBC_XCLK_OUT(), .CAN_RXBUS_USBA_DATA1_MGPIO3A_OE(), 
        .CAN_TX_EBL_USBA_DATA2_MGPIO4A_OE(), 
        .CAN_TXBUS_USBA_DATA0_MGPIO2A_OE(), .DM_OE({nc306, nc307, 
        nc308}), .DRAM_DQ_OE({nc309, nc310, nc311, nc312, nc313, nc314, 
        nc315, nc316, nc317, nc318, nc319, nc320, nc321, nc322, nc323, 
        nc324, nc325, nc326}), .DRAM_DQS_OE({nc327, nc328, nc329}), 
        .I2C0_SCL_USBC_DATA1_MGPIO31B_OE(), 
        .I2C0_SDA_USBC_DATA0_MGPIO30B_OE(), 
        .I2C1_SCL_USBA_DATA4_MGPIO1A_OE(), 
        .I2C1_SDA_USBA_DATA3_MGPIO0A_OE(), 
        .MMUART0_CTS_USBC_DATA7_MGPIO19B_OE(), 
        .MMUART0_DCD_MGPIO22B_OE(), .MMUART0_DSR_MGPIO20B_OE(), 
        .MMUART0_DTR_USBC_DATA6_MGPIO18B_OE(), .MMUART0_RI_MGPIO21B_OE(
        ), .MMUART0_RTS_USBC_DATA5_MGPIO17B_OE(), 
        .MMUART0_RXD_USBC_STP_MGPIO28B_OE(), 
        .MMUART0_SCK_USBC_NXT_MGPIO29B_OE(), 
        .MMUART0_TXD_USBC_DIR_MGPIO27B_OE(
        MSS_ADLIB_INST_MMUART0_TXD_USBC_DIR_MGPIO27B_OE), 
        .MMUART1_RXD_USBC_DATA3_MGPIO26B_OE(), 
        .MMUART1_SCK_USBC_DATA4_MGPIO25B_OE(), 
        .MMUART1_TXD_USBC_DATA2_MGPIO24B_OE(), 
        .RGMII_GTX_CLK_RMII_CLK_USBB_XCLK_OE(), .RGMII_MDC_RMII_MDC_OE(
        ), .RGMII_MDIO_RMII_MDIO_USBB_DATA7_OE(), .RGMII_RX_CLK_OE(), 
        .RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_OE(), 
        .RGMII_RXD0_RMII_RXD0_USBB_DATA0_OE(), 
        .RGMII_RXD1_RMII_RXD1_USBB_DATA1_OE(), 
        .RGMII_RXD2_RMII_RX_ER_USBB_DATA3_OE(), 
        .RGMII_RXD3_USBB_DATA4_OE(), .RGMII_TX_CLK_OE(), 
        .RGMII_TX_CTL_RMII_TX_EN_USBB_NXT_OE(), 
        .RGMII_TXD0_RMII_TXD0_USBB_DIR_OE(), 
        .RGMII_TXD1_RMII_TXD1_USBB_STP_OE(), .RGMII_TXD2_USBB_DATA5_OE(
        ), .RGMII_TXD3_USBB_DATA6_OE(), .SPI0_SCK_USBA_XCLK_OE(), 
        .SPI0_SDI_USBA_DIR_MGPIO5A_OE(), .SPI0_SDO_USBA_STP_MGPIO6A_OE(
        ), .SPI0_SS0_USBA_NXT_MGPIO7A_OE(), 
        .SPI0_SS1_USBA_DATA5_MGPIO8A_OE(), 
        .SPI0_SS2_USBA_DATA6_MGPIO9A_OE(), 
        .SPI0_SS3_USBA_DATA7_MGPIO10A_OE(), .SPI1_SCK_OE(), 
        .SPI1_SDI_MGPIO11A_OE(), .SPI1_SDO_MGPIO12A_OE(), 
        .SPI1_SS0_MGPIO13A_OE(), .SPI1_SS1_MGPIO14A_OE(), 
        .SPI1_SS2_MGPIO15A_OE(), .SPI1_SS3_MGPIO16A_OE(), 
        .SPI1_SS4_MGPIO17A_OE(), .SPI1_SS5_MGPIO18A_OE(), 
        .SPI1_SS6_MGPIO23A_OE(), .SPI1_SS7_MGPIO24A_OE(), 
        .USBC_XCLK_OE());
    GND GND (.Y(GND_net_1));
    TRIBUFF MMUART_0_TXD_PAD (.D(
        MSS_ADLIB_INST_MMUART0_TXD_USBC_DIR_MGPIO27B_OUT), .E(
        MSS_ADLIB_INST_MMUART0_TXD_USBC_DIR_MGPIO27B_OE), .PAD(
        MMUART_0_TXD));
    
endmodule


module CoreGPIO_Z3(
       CoreAPB3_0_APBmslave2_PWDATA,
       GPIO_IN_c,
       GPIO_OUT_net_2,
       CoreAPB3_0_APBmslave2_PADDR,
       iPSELS_2,
       GPOUT_reg_31,
       GPOUT_reg_30,
       GPOUT_reg_29,
       GPOUT_reg_28,
       GPOUT_reg_27,
       GPOUT_reg_26,
       GPOUT_reg_25,
       GPOUT_reg_24,
       GPOUT_reg_23,
       GPOUT_reg_22,
       GPOUT_reg_21,
       GPOUT_reg_20,
       GPOUT_reg_19,
       GPOUT_reg_18,
       GPOUT_reg_17,
       GPOUT_reg_16,
       GPOUT_reg_15,
       GPOUT_reg_14,
       GPOUT_reg_13,
       GPOUT_reg_12,
       GPOUT_reg_11,
       GPOUT_reg_10,
       GPOUT_reg_9,
       GPOUT_reg_8,
       GPOUT_reg_6,
       GPOUT_reg_5,
       GPOUT_reg_4,
       GPOUT_reg_2,
       GPOUT_reg_1,
       GPOUT_reg_0,
       \CONFIG_reg[6]_1 ,
       \CONFIG_reg[5]_1 ,
       \CONFIG_reg[3]_1 ,
       \CONFIG_reg[2]_1 ,
       \CONFIG_reg[1]_1 ,
       \CONFIG_reg[0]_1 ,
       INTR_reg_23,
       INTR_reg_24,
       INTR_reg_25,
       INTR_reg_26,
       INTR_reg_27,
       INTR_reg_28,
       INTR_reg_29,
       INTR_reg_30,
       INTR_reg_31,
       INTR_reg_8,
       INTR_reg_9,
       INTR_reg_10,
       INTR_reg_11,
       INTR_reg_12,
       INTR_reg_13,
       INTR_reg_14,
       INTR_reg_15,
       INTR_reg_16,
       INTR_reg_17,
       INTR_reg_18,
       INTR_reg_19,
       INTR_reg_20,
       INTR_reg_21,
       INTR_reg_22,
       INTR_reg_0,
       INTR_reg_1,
       INTR_reg_2,
       INTR_reg_4,
       INTR_reg_5,
       INTR_reg_6,
       INTR_reg_7,
       gpin3_5,
       gpin3_6,
       gpin3_0,
       gpin3_1,
       gpin3_2,
       gpin3_3,
       FIC_MSS_0_FIC_0_APB_MASTER_PADDR_2,
       FIC_MSS_0_FIC_0_APB_MASTER_PADDR_0,
       MSS_RESET_N_F2M_c,
       FCCC_0_GL1,
       PRDATA_N_3_0,
       N_4801,
       N_4762,
       N_4706,
       N_4682,
       N_4852,
       N_4857,
       N_4825,
       N_4736,
       N_4705,
       N_4858,
       N_4819,
       N_4851,
       N_4761,
       N_4802,
       N_4738,
       N_4880,
       N_4879,
       N_4877,
       N_4735,
       N_4881,
       N_4798,
       N_4797,
       N_4796,
       N_4758,
       N_4757,
       N_4756,
       N_4878,
       N_4823,
       N_4876,
       N_4734,
       N_4733,
       N_4732,
       N_4731,
       N_4676,
       N_4675,
       N_4795,
       N_4826,
       N_4701,
       N_4882,
       N_4755,
       N_4702,
       N_4853,
       N_4677,
       N_4820,
       N_4854,
       N_4759,
       N_4678,
       N_4760,
       N_4681,
       N_4824,
       N_4703,
       N_4737,
       N_4704,
       N_4679,
       N_4699,
       N_4799,
       N_4855,
       N_4680,
       N_4875,
       N_4800,
       N_4822,
       N_4821,
       N_4700,
       N_4856,
       N_610,
       N_603,
       PRDATA_m1_e_1,
       N_245,
       N_452,
       N_247,
       CoreAPB3_0_APBmslave5_PSELx,
       wen_0,
       \CONFIG_reg[4]2_0_a4_0_a2_0_RNIBB9M2 
    );
input  [31:0] CoreAPB3_0_APBmslave2_PWDATA;
input  [6:0] GPIO_IN_c;
output [6:0] GPIO_OUT_net_2;
input  [7:0] CoreAPB3_0_APBmslave2_PADDR;
input  [5:5] iPSELS_2;
output GPOUT_reg_31;
output GPOUT_reg_30;
output GPOUT_reg_29;
output GPOUT_reg_28;
output GPOUT_reg_27;
output GPOUT_reg_26;
output GPOUT_reg_25;
output GPOUT_reg_24;
output GPOUT_reg_23;
output GPOUT_reg_22;
output GPOUT_reg_21;
output GPOUT_reg_20;
output GPOUT_reg_19;
output GPOUT_reg_18;
output GPOUT_reg_17;
output GPOUT_reg_16;
output GPOUT_reg_15;
output GPOUT_reg_14;
output GPOUT_reg_13;
output GPOUT_reg_12;
output GPOUT_reg_11;
output GPOUT_reg_10;
output GPOUT_reg_9;
output GPOUT_reg_8;
output GPOUT_reg_6;
output GPOUT_reg_5;
output GPOUT_reg_4;
output GPOUT_reg_2;
output GPOUT_reg_1;
output GPOUT_reg_0;
output \CONFIG_reg[6]_1 ;
output \CONFIG_reg[5]_1 ;
output \CONFIG_reg[3]_1 ;
output \CONFIG_reg[2]_1 ;
output \CONFIG_reg[1]_1 ;
output \CONFIG_reg[0]_1 ;
output INTR_reg_23;
output INTR_reg_24;
output INTR_reg_25;
output INTR_reg_26;
output INTR_reg_27;
output INTR_reg_28;
output INTR_reg_29;
output INTR_reg_30;
output INTR_reg_31;
output INTR_reg_8;
output INTR_reg_9;
output INTR_reg_10;
output INTR_reg_11;
output INTR_reg_12;
output INTR_reg_13;
output INTR_reg_14;
output INTR_reg_15;
output INTR_reg_16;
output INTR_reg_17;
output INTR_reg_18;
output INTR_reg_19;
output INTR_reg_20;
output INTR_reg_21;
output INTR_reg_22;
output INTR_reg_0;
output INTR_reg_1;
output INTR_reg_2;
output INTR_reg_4;
output INTR_reg_5;
output INTR_reg_6;
output INTR_reg_7;
output gpin3_5;
output gpin3_6;
output gpin3_0;
output gpin3_1;
output gpin3_2;
output gpin3_3;
input  FIC_MSS_0_FIC_0_APB_MASTER_PADDR_2;
input  FIC_MSS_0_FIC_0_APB_MASTER_PADDR_0;
input  MSS_RESET_N_F2M_c;
input  FCCC_0_GL1;
output PRDATA_N_3_0;
output N_4801;
output N_4762;
output N_4706;
output N_4682;
output N_4852;
output N_4857;
output N_4825;
output N_4736;
output N_4705;
output N_4858;
output N_4819;
output N_4851;
output N_4761;
output N_4802;
output N_4738;
output N_4880;
output N_4879;
output N_4877;
output N_4735;
output N_4881;
output N_4798;
output N_4797;
output N_4796;
output N_4758;
output N_4757;
output N_4756;
output N_4878;
output N_4823;
output N_4876;
output N_4734;
output N_4733;
output N_4732;
output N_4731;
output N_4676;
output N_4675;
output N_4795;
output N_4826;
output N_4701;
output N_4882;
output N_4755;
output N_4702;
output N_4853;
output N_4677;
output N_4820;
output N_4854;
output N_4759;
output N_4678;
output N_4760;
output N_4681;
output N_4824;
output N_4703;
output N_4737;
output N_4704;
output N_4679;
output N_4699;
output N_4799;
output N_4855;
output N_4680;
output N_4875;
output N_4800;
output N_4822;
output N_4821;
output N_4700;
output N_4856;
output N_610;
output N_603;
output PRDATA_m1_e_1;
output N_245;
output N_452;
output N_247;
input  CoreAPB3_0_APBmslave5_PSELx;
input  wen_0;
output \CONFIG_reg[4]2_0_a4_0_a2_0_RNIBB9M2 ;

    wire \edge_pos[31] , VCC_net_1, \edge_neg_443[31] , 
        edge_pos_2_sqmuxa_19_i_1, GND_net_1, \edge_pos[30] , 
        \edge_neg_429[30] , edge_neg_2_sqmuxa_6_i_1, \edge_pos[29] , 
        \edge_neg_415[29] , N_190, \edge_pos[28] , N_87_i_0, N_163, 
        \edge_neg[27] , N_5912_i_0, N_161, \edge_pos[26] , N_106_i_0, 
        N_159, \edge_neg[25] , N_5911_i_0, N_157, \edge_pos[24] , 
        N_100_i_0, N_155, \edge_neg[23] , N_96_i_0, 
        edge_pos_2_sqmuxa_26_i_1, \edge_neg[22] , \edge_neg_317[22] , 
        N_200, \edge_neg[21] , \edge_neg_303[21] , N_198, 
        \edge_neg[20] , \edge_neg_289[20] , N_196, \edge_neg[19] , 
        \edge_neg_275[19] , N_194, \edge_neg[18] , \edge_neg_261[18] , 
        N_192, \edge_neg[17] , \edge_neg_247[17] , 
        edge_pos_2_sqmuxa_30_i_1, \edge_neg[16] , \edge_neg_233[16] , 
        edge_pos_2_sqmuxa_29_i_1, \edge_neg[14] , \edge_neg_205[14] , 
        edge_pos_2_sqmuxa_8_i_1, \edge_neg[13] , \edge_neg_191[13] , 
        edge_pos_2_sqmuxa_9_i_1, \edge_neg[12] , \edge_neg_177[12] , 
        N_188, \edge_neg[11] , \edge_neg_163[11] , N_186, 
        \edge_pos[10] , \edge_neg_149[10] , N_184, \edge_neg[9] , 
        \edge_neg_135[9] , N_182, \edge_pos[8] , \edge_neg_121[8] , 
        edge_neg_2_sqmuxa_4_i_1, \edge_pos[7] , N_83_i_0, 
        edge_pos_2_sqmuxa_1_i_1, \edge_both[6] , N_22_i_0, N_78, 
        \edge_both[5] , N_89, N_76, \edge_both[4] , N_91, N_84, 
        \edge_both[3] , \edge_both_51_iv_i_0[3] , 
        edge_both_2_sqmuxa_12_i_1, \edge_both[2] , N_93, N_86, 
        \edge_both[1] , N_95, N_82, \edge_both[0] , N_97, N_80, 
        \edge_neg[6] , N_113, N_62, \edge_neg[5] , N_115, N_60, 
        \edge_neg[4] , N_117, N_58, \edge_neg[3] , 
        \edge_neg_51_iv_i_1[3] , N_81, \edge_neg[2] , N_119, N_56, 
        \edge_neg[1] , N_121, N_54, \edge_neg[0] , N_123, N_52, 
        \edge_neg[15] , \edge_pos_219[15] , edge_pos_2_sqmuxa_7_i_1, 
        \edge_pos[6] , N_99, N_72, \edge_pos[5] , N_101, N_70, 
        \edge_pos[4] , N_103, N_68, \edge_pos[3] , N_73, N_79, 
        \edge_pos[2] , N_105, N_64, \edge_pos[1] , N_107, N_66, 
        \edge_pos[0] , N_109, N_74, GPOUT_reg_0_sqmuxa, \GPOUT_reg[7] , 
        \GPOUT_reg[3] , \CONFIG_reg[31][0] , \CONFIG_reg[31]2 , 
        \CONFIG_reg[31][1] , \CONFIG_reg[31][2] , \CONFIG_reg[31][3] , 
        \CONFIG_reg[31][4] , \CONFIG_reg[31][5] , \CONFIG_reg[31][6] , 
        \CONFIG_reg[31][7] , \CONFIG_reg[30][0] , \CONFIG_reg[30]2 , 
        \CONFIG_reg[30][1] , \CONFIG_reg[30][2] , \CONFIG_reg[30][3] , 
        \CONFIG_reg[30][4] , \CONFIG_reg[30][5] , \CONFIG_reg[30][6] , 
        \CONFIG_reg[30][7] , \CONFIG_reg[29][0] , \CONFIG_reg[29]2 , 
        \CONFIG_reg[29][1] , \CONFIG_reg[29][2] , \CONFIG_reg[29][3] , 
        \CONFIG_reg[29][4] , \CONFIG_reg[29][5] , \CONFIG_reg[29][6] , 
        \CONFIG_reg[29][7] , \CONFIG_reg[28][0] , \CONFIG_reg[28]2 , 
        \CONFIG_reg[28][1] , \CONFIG_reg[28][2] , \CONFIG_reg[28][3] , 
        \CONFIG_reg[28][4] , \CONFIG_reg[28][5] , \CONFIG_reg[28][6] , 
        \CONFIG_reg[28][7] , \CONFIG_reg[27][0] , \CONFIG_reg[27]2 , 
        \CONFIG_reg[27][1] , \CONFIG_reg[27][2] , \CONFIG_reg[27][3] , 
        \CONFIG_reg[27][4] , \CONFIG_reg[27][5] , \CONFIG_reg[27][6] , 
        \CONFIG_reg[27][7] , \CONFIG_reg[26][0] , \CONFIG_reg[26]2 , 
        \CONFIG_reg[26][1] , \CONFIG_reg[26][2] , \CONFIG_reg[26][3] , 
        \CONFIG_reg[26][4] , \CONFIG_reg[26][5] , \CONFIG_reg[26][6] , 
        \CONFIG_reg[26][7] , \CONFIG_reg[25][0] , \CONFIG_reg[25]2 , 
        \CONFIG_reg[25][1] , \CONFIG_reg[25][2] , \CONFIG_reg[25][3] , 
        \CONFIG_reg[25][4] , \CONFIG_reg[25][5] , \CONFIG_reg[25][6] , 
        \CONFIG_reg[25][7] , \CONFIG_reg[24][0] , \CONFIG_reg[24]2 , 
        \CONFIG_reg[24][1] , \CONFIG_reg[24][2] , \CONFIG_reg[24][3] , 
        \CONFIG_reg[24][4] , \CONFIG_reg[24][5] , \CONFIG_reg[24][6] , 
        \CONFIG_reg[24][7] , \CONFIG_reg[23][0] , \CONFIG_reg[23]2 , 
        \CONFIG_reg[23][1] , \CONFIG_reg[23][2] , \CONFIG_reg[23][3] , 
        \CONFIG_reg[23][4] , \CONFIG_reg[23][5] , \CONFIG_reg[23][6] , 
        \CONFIG_reg[23][7] , \CONFIG_reg[22][0] , \CONFIG_reg[22]2 , 
        \CONFIG_reg[22][1] , \CONFIG_reg[22][2] , \CONFIG_reg[22][3] , 
        \CONFIG_reg[22][4] , \CONFIG_reg[22][5] , \CONFIG_reg[22][6] , 
        \CONFIG_reg[22][7] , \CONFIG_reg[21][0] , \CONFIG_reg[21]2 , 
        \CONFIG_reg[21][1] , \CONFIG_reg[21][2] , \CONFIG_reg[21][3] , 
        \CONFIG_reg[21][4] , \CONFIG_reg[21][5] , \CONFIG_reg[21][6] , 
        \CONFIG_reg[21][7] , \CONFIG_reg[20][0] , \CONFIG_reg[20]2 , 
        \CONFIG_reg[20][1] , \CONFIG_reg[20][2] , \CONFIG_reg[20][3] , 
        \CONFIG_reg[20][4] , \CONFIG_reg[20][5] , \CONFIG_reg[20][6] , 
        \CONFIG_reg[20][7] , \CONFIG_reg[19][0] , \CONFIG_reg[19]2 , 
        \CONFIG_reg[19][1] , \CONFIG_reg[19][2] , \CONFIG_reg[19][3] , 
        \CONFIG_reg[19][4] , \CONFIG_reg[19][5] , \CONFIG_reg[19][6] , 
        \CONFIG_reg[19][7] , \CONFIG_reg[18][0] , \CONFIG_reg[18]2 , 
        \CONFIG_reg[18][1] , \CONFIG_reg[18][2] , \CONFIG_reg[18][3] , 
        \CONFIG_reg[18][4] , \CONFIG_reg[18][5] , \CONFIG_reg[18][6] , 
        \CONFIG_reg[18][7] , \CONFIG_reg[17][0] , \CONFIG_reg[17]2 , 
        \CONFIG_reg[17][1] , \CONFIG_reg[17][2] , \CONFIG_reg[17][3] , 
        \CONFIG_reg[17][4] , \CONFIG_reg[17][5] , \CONFIG_reg[17][6] , 
        \CONFIG_reg[17][7] , \CONFIG_reg[16][0] , \CONFIG_reg[16]2 , 
        \CONFIG_reg[16][1] , \CONFIG_reg[16][2] , \CONFIG_reg[16][3] , 
        \CONFIG_reg[16][4] , \CONFIG_reg[16][5] , \CONFIG_reg[16][6] , 
        \CONFIG_reg[16][7] , \CONFIG_reg[15][0] , \CONFIG_reg[15]2 , 
        \CONFIG_reg[15][1] , \CONFIG_reg[15][2] , \CONFIG_reg[15][3] , 
        \CONFIG_reg[15][4] , \CONFIG_reg[15][5] , \CONFIG_reg[15][6] , 
        \CONFIG_reg[15][7] , \CONFIG_reg[14][0] , \CONFIG_reg[14]2 , 
        \CONFIG_reg[14][1] , \CONFIG_reg[14][2] , \CONFIG_reg[14][3] , 
        \CONFIG_reg[14][4] , \CONFIG_reg[14][5] , \CONFIG_reg[14][6] , 
        \CONFIG_reg[14][7] , \CONFIG_reg[13][0] , \CONFIG_reg[13]2 , 
        \CONFIG_reg[13][1] , \CONFIG_reg[13][2] , \CONFIG_reg[13][3] , 
        \CONFIG_reg[13][4] , \CONFIG_reg[13][5] , \CONFIG_reg[13][6] , 
        \CONFIG_reg[13][7] , \CONFIG_reg[12][0] , \CONFIG_reg[12]2 , 
        \CONFIG_reg[12][1] , \CONFIG_reg[12][2] , \CONFIG_reg[12][3] , 
        \CONFIG_reg[12][4] , \CONFIG_reg[12][5] , \CONFIG_reg[12][6] , 
        \CONFIG_reg[12][7] , \CONFIG_reg[11][0] , \CONFIG_reg[11]2 , 
        \CONFIG_reg[11][1] , \CONFIG_reg[11][2] , \CONFIG_reg[11][3] , 
        \CONFIG_reg[11][4] , \CONFIG_reg[11][5] , \CONFIG_reg[11][6] , 
        \CONFIG_reg[11][7] , \CONFIG_reg[10][0] , \CONFIG_reg[10]2 , 
        \CONFIG_reg[10][1] , \CONFIG_reg[10][2] , \CONFIG_reg[10][3] , 
        \CONFIG_reg[10][4] , \CONFIG_reg[10][5] , \CONFIG_reg[10][6] , 
        \CONFIG_reg[10][7] , \CONFIG_reg[9][0] , \CONFIG_reg[9]2 , 
        \CONFIG_reg[9][1] , \CONFIG_reg[9][2] , \CONFIG_reg[9][3] , 
        \CONFIG_reg[9][4] , \CONFIG_reg[9][5] , \CONFIG_reg[9][6] , 
        \CONFIG_reg[9][7] , \CONFIG_reg[8][0] , \CONFIG_reg[8]2 , 
        \CONFIG_reg[8][1] , \CONFIG_reg[8][2] , \CONFIG_reg[8][3] , 
        \CONFIG_reg[8][4] , \CONFIG_reg[8][5] , \CONFIG_reg[8][6] , 
        \CONFIG_reg[8][7] , \CONFIG_reg[7][0] , \CONFIG_reg[7]2 , 
        \CONFIG_reg[7][1] , \CONFIG_reg[7][2] , \CONFIG_reg[7][3] , 
        \CONFIG_reg[7][4] , \CONFIG_reg[7][5] , \CONFIG_reg[7][6] , 
        \CONFIG_reg[7][7] , \CONFIG_reg[6][0] , \CONFIG_reg[6]2 , 
        \CONFIG_reg[6][2] , \CONFIG_reg[6][3] , \CONFIG_reg[6][4] , 
        \CONFIG_reg[6][5] , \CONFIG_reg[6][6] , \CONFIG_reg[6][7] , 
        \CONFIG_reg[5][0] , \CONFIG_reg[5]2 , \CONFIG_reg[5][2] , 
        \CONFIG_reg[5][3] , \CONFIG_reg[5][4] , \CONFIG_reg[5][5] , 
        \CONFIG_reg[5][6] , \CONFIG_reg[5][7] , \CONFIG_reg[4][0] , 
        \CONFIG_reg[4]2 , \CONFIG_reg[4][1] , \CONFIG_reg[4][2] , 
        \CONFIG_reg[4][3] , \CONFIG_reg[4][4] , \CONFIG_reg[4][5] , 
        \CONFIG_reg[4][6] , \CONFIG_reg[4][7] , \CONFIG_reg[3][0] , 
        \CONFIG_reg[3]2 , \CONFIG_reg[3][2] , \CONFIG_reg[3][3] , 
        \CONFIG_reg[3][4] , \CONFIG_reg[3][5] , \CONFIG_reg[3][6] , 
        \CONFIG_reg[3][7] , \CONFIG_reg[2][0] , \CONFIG_reg[2]2 , 
        \CONFIG_reg[2][2] , \CONFIG_reg[2][3] , \CONFIG_reg[2][4] , 
        \CONFIG_reg[2][5] , \CONFIG_reg[2][6] , \CONFIG_reg[2][7] , 
        \CONFIG_reg[1][0] , \CONFIG_reg[1]2 , \CONFIG_reg[1][2] , 
        \CONFIG_reg[1][3] , \CONFIG_reg[1][4] , \CONFIG_reg[1][5] , 
        \CONFIG_reg[1][6] , \CONFIG_reg[1][7] , \CONFIG_reg[0][0] , 
        \CONFIG_reg[0]2 , \CONFIG_reg[0][2] , \CONFIG_reg[0][3] , 
        \CONFIG_reg[0][4] , \CONFIG_reg[0][5] , \CONFIG_reg[0][6] , 
        \CONFIG_reg[0][7] , \INTR_reg_308[23] , \INTR_reg_321[24] , 
        \INTR_reg_334[25] , \INTR_reg_347[26] , \INTR_reg_360[27] , 
        \INTR_reg_373[28] , \INTR_reg_386[29] , \INTR_reg_399[30] , 
        \INTR_reg_412[31] , \INTR_reg_113[8] , \INTR_reg_126[9] , 
        \INTR_reg_139[10] , \INTR_reg_152[11] , \INTR_reg_165[12] , 
        \INTR_reg_178[13] , \INTR_reg_191[14] , \INTR_reg_204[15] , 
        \INTR_reg_217[16] , \INTR_reg_230[17] , \INTR_reg_243[18] , 
        \INTR_reg_256[19] , \INTR_reg_269[20] , \INTR_reg_282[21] , 
        \INTR_reg_295[22] , \INTR_reg_9[0] , \INTR_reg_22[1] , 
        \INTR_reg_35[2] , \INTR_reg[3] , \INTR_reg_48[3] , 
        \INTR_reg_61[4] , \INTR_reg_74[5] , \INTR_reg_87[6] , 
        \INTR_reg_100[7] , \gpin3[4] , \gpin2[4] , \gpin2[5] , 
        \gpin2[6] , \gpin2[0] , \gpin2[1] , \gpin2[2] , \gpin2[3] , 
        \gpin1[4] , \gpin1[5] , \gpin1[6] , \gpin1[0] , \gpin1[1] , 
        \gpin1[2] , \gpin1[3] , un34_intr_u_ns_1, 
        \INTR_reg_87_0_0_0_tz_1[6] , N_5939, \INTR_reg_87_0_0_0_tz[6] , 
        \INTR_reg_74_0_0_0_tz_1[5] , N_5940, \INTR_reg_74_0_0_0_tz[5] , 
        \INTR_reg_61_0_0_0_tz_1[4] , N_179, \INTR_reg_61_0_0_0_tz[4] , 
        \INTR_reg_35_0_0_0_tz_1[2] , N_178, \INTR_reg_35_0_0_0_tz[2] , 
        \INTR_reg_22_0_0_0_tz_1[1] , N_177, \INTR_reg_22_0_0_0_tz[1] , 
        \INTR_reg_9_0_0_0_tz_1[0] , N_5941, \INTR_reg_9_0_0_0_tz[0] , 
        \CONFIG_reg_o_2_18_1_1[6] , \CONFIG_reg_o_2_13_1_1[7] , 
        \CONFIG_reg_o_2_6_1_1[7] , \CONFIG_reg_o_2_3_1_1[7] , 
        \CONFIG_reg_o_2_25_1_1[1] , \CONFIG_reg_o_2_25_1_1[6] , 
        \CONFIG_reg_o_2_21_1_1[6] , \CONFIG_reg_o_2_10_1_1[5] , 
        \CONFIG_reg_o_2_6_1_1[6] , \CONFIG_reg_o_2_25_1_1[7] , 
        \CONFIG_reg_o_2_21_1[0] , \CONFIG_reg_o_2_25_1_1[0] , 
        \CONFIG_reg_o_2_13_1_1[6] , \CONFIG_reg_o_2_18_1_1[7] , 
        \CONFIG_reg_o_2_10_1_1[7] , \CONFIG_reg_o_2_28_1_1[5] , 
        \CONFIG_reg_o_2_28_1_1[4] , \CONFIG_reg_o_2_28_1_1[2] , 
        \CONFIG_reg_o_2_10_1_1[4] , \CONFIG_reg_o_2_28_1_1[6] , 
        \CONFIG_reg_o_2_18_1[3] , \CONFIG_reg_o_2_18_1_1[2] , 
        \CONFIG_reg_o_2_18_1_1[1] , \CONFIG_reg_o_2_13_1_1[3] , 
        \CONFIG_reg_o_2_13_1_1[2] , \CONFIG_reg_o_2_13_1_1[1] , 
        \CONFIG_reg_o_2_28_1_1[3] , \CONFIG_reg_o_2_21_1[4] , 
        \CONFIG_reg_o_2_28_1_1[1] , \CONFIG_reg_o_2_10_1_1[3] , 
        \CONFIG_reg_o_2_10_1_1[2] , \CONFIG_reg_o_2_10_1_1[1] , 
        \CONFIG_reg_o_2_10_1_1[0] , \CONFIG_reg_o_2_3_1_1[1] , 
        \CONFIG_reg_o_2_3_1[0] , \CONFIG_reg_o_2_18_1[0] , 
        \CONFIG_reg_o_2_21_1_1[7] , \CONFIG_reg_o_2_6_1_1[2] , 
        \CONFIG_reg_o_2_28_1_1[7] , \CONFIG_reg_o_2_13_1_1[0] , 
        \CONFIG_reg_o_2_6_1[3] , \CONFIG_reg_o_2_25_1_1[2] , 
        \CONFIG_reg_o_2_3_1_1[2] , \CONFIG_reg_o_2_21_1_1[1] , 
        \CONFIG_reg_o_2_25_1_1[3] , \CONFIG_reg_o_2_13_1_1[4] , 
        \CONFIG_reg_o_2_3_1[3] , \CONFIG_reg_o_2_13_1_1[5] , 
        \CONFIG_reg_o_2_3_1_1[6] , \CONFIG_reg_o_2_21_1_1[5] , 
        \CONFIG_reg_o_2_6_1[4] , \CONFIG_reg_o_2_10_1_1[6] , 
        \CONFIG_reg_o_2_6_1_1[5] , \CONFIG_reg_o_2_3_1[4] , 
        \CONFIG_reg_o_2_6_1[0] , \CONFIG_reg_o_2_18_1[4] , 
        \CONFIG_reg_o_2_25_1_1[4] , \CONFIG_reg_o_2_3_1_1[5] , 
        \CONFIG_reg_o_2_28_1_1[0] , \CONFIG_reg_o_2_18_1_1[5] , 
        \CONFIG_reg_o_2_21_1[3] , \CONFIG_reg_o_2_21_1_1[2] , 
        \CONFIG_reg_o_2_6_1_1[1] , \CONFIG_reg_o_2_25_1_1[5] , 
        un34_intr_u_bm, un34_intr, r_m1_e_1_0, 
        un5_PRDATA_o_0_a2_0_o2_out, N_395, N_396, N_397, N_398, N_399, 
        N_400, N_401, N_402, N_405, N_406, N_139_i, N_141_i, N_142_i, 
        N_143_i, N_144_i, N_605, N_606, N_686, N_687, N_688, N_689, 
        N_252_i, N_253_i, N_4549, N_172, N_173, N_174, N_175, N_5938, 
        N_171, GEN_m3_e_1, N_243, \INTR_reg_217_0_o2_0[16] , 
        \INTR_reg_139_0_o2_0[10] , \INTR_reg_152_0_o2_0[11] , 
        \INTR_reg_113_0_o2_0[8] , \INTR_reg_191_0_o2_0[14] , 
        \INTR_reg_334_0_o2_0[25] , \INTR_reg_373_0_o2_0[28] , 
        \INTR_reg_412_0_o2_0[31] , \INTR_reg_282_0_o2_0[21] , 
        \INTR_reg_256_0_o2_0[19] , \INTR_reg_321_0_o2_0[24] , 
        \INTR_reg_347_0_o2_0[26] , \INTR_reg_399_0_o2_0[30] , 
        \INTR_reg_269_0_o2_0[20] , \INTR_reg_295_0_o2_0[22] , 
        \INTR_reg_165_0_o2_0[12] , \INTR_reg_178_0_o2_0[13] , 
        \INTR_reg_204_0_o2_0[15] , \INTR_reg_386_0_o2_0[29] , 
        \INTR_reg_308_0_o2_0[23] , \INTR_reg_126_0_o2_0[9] , 
        \INTR_reg_360_0_o2_0[27] , \INTR_reg_230_0_o2_0[17] , 
        \INTR_reg_100_0_o2_0[7] , \INTR_reg_243_0_o2_0[18] , 
        \INTR_reg_217_0_o2_1[16] , \INTR_reg_139_0_o2_1[10] , 
        \INTR_reg_152_0_o2_1[11] , \INTR_reg_113_0_o2_1[8] , 
        \INTR_reg_191_0_o2_1[14] , \INTR_reg_334_0_o2_1[25] , 
        \INTR_reg_373_0_o2_1[28] , \INTR_reg_412_0_o2_1[31] , 
        \INTR_reg_282_0_o2_1[21] , \INTR_reg_256_0_o2_1[19] , 
        \INTR_reg_321_0_o2_1[24] , \INTR_reg_347_0_o2_1[26] , 
        \INTR_reg_399_0_o2_1[30] , \INTR_reg_269_0_o2_1[20] , 
        \INTR_reg_295_0_o2_1[22] , \INTR_reg_165_0_o2_1[12] , 
        \INTR_reg_178_0_o2_1[13] , \INTR_reg_204_0_o2_1[15] , 
        \INTR_reg_386_0_o2_1[29] , \INTR_reg_308_0_o2_1[23] , 
        \INTR_reg_126_0_o2_1[9] , \INTR_reg_360_0_o2_1[27] , 
        \INTR_reg_230_0_o2_1[17] , \INTR_reg_100_0_o2_1[7] , 
        \INTR_reg_243_0_o2_1[18] , edge_N_5_mux, N_598, N_604, N_678;
    
    SLE \xhdl1.GEN_BITS[18].APB_32.INTR_reg[18]  (.D(
        \INTR_reg_243[18] ), .CLK(FCCC_0_GL1), .EN(VCC_net_1), .ALn(
        MSS_RESET_N_F2M_c), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(INTR_reg_18));
    SLE \xhdl1.GEN_BITS[2].gpin1[2]  (.D(GPIO_IN_c[2]), .CLK(
        FCCC_0_GL1), .EN(VCC_net_1), .ALn(MSS_RESET_N_F2M_c), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\gpin1[2] ));
    SLE \xhdl1.GEN_BITS[16].APB_32.edge_both[16]  (.D(
        \edge_neg_233[16] ), .CLK(FCCC_0_GL1), .EN(
        edge_pos_2_sqmuxa_29_i_1), .ALn(MSS_RESET_N_F2M_c), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\edge_neg[16] ));
    CFG3 #( .INIT(8'hFB) )  edge_neg_2_sqmuxa_9_i_0 (.A(edge_N_5_mux), 
        .B(\CONFIG_reg[3][3] ), .C(N_686), .Y(N_81));
    CFG4 #( .INIT(16'h4000) )  
        \xhdl1.GEN_BITS[13].REG_GEN.CONFIG_reg[13]2_0_a4_0_a2  (.A(
        CoreAPB3_0_APBmslave2_PADDR[3]), .B(
        CoreAPB3_0_APBmslave2_PADDR[2]), .C(N_604), .D(N_605), .Y(
        \CONFIG_reg[13]2 ));
    SLE \xhdl1.GEN_BITS[26].REG_GEN.CONFIG_reg[26][4]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[4]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[26]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[26][4] ));
    CFG2 #( .INIT(4'h4) )  edge_neg_2_sqmuxa_8_i_a2 (.A(\gpin2[4] ), 
        .B(\gpin3[4] ), .Y(N_397));
    CFG4 #( .INIT(16'h0ACC) )  
        \xhdl1.GEN_BITS[3].APB_32.INTR_reg_48_0[3]  (.A(\INTR_reg[3] ), 
        .B(un34_intr), .C(CoreAPB3_0_APBmslave2_PWDATA[3]), .D(
        edge_N_5_mux), .Y(\INTR_reg_48[3] ));
    CFG4 #( .INIT(16'h0F35) )  
        \xhdl1.GEN_BITS[19].REG_GEN.CONFIG_reg[19]_RNIGR391[2]  (.A(
        \CONFIG_reg[3][2] ), .B(\CONFIG_reg[19][2] ), .C(
        CoreAPB3_0_APBmslave2_PADDR[6]), .D(
        CoreAPB3_0_APBmslave2_PADDR[5]), .Y(\CONFIG_reg_o_2_25_1_1[2] )
        );
    SLE \xhdl1.GEN_BITS[11].REG_GEN.CONFIG_reg[11][1]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[1]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[11]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[11][1] ));
    SLE \xhdl1.GEN_BITS[13].APB_32.GPOUT_reg[13]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[13]), .CLK(FCCC_0_GL1), .EN(
        GPOUT_reg_0_sqmuxa), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        GPOUT_reg_13));
    CFG4 #( .INIT(16'h0F35) )  
        \xhdl1.GEN_BITS[20].REG_GEN.CONFIG_reg[20]_RNI89V31[5]  (.A(
        \CONFIG_reg[4][5] ), .B(\CONFIG_reg[20][5] ), .C(
        CoreAPB3_0_APBmslave2_PADDR[6]), .D(
        CoreAPB3_0_APBmslave2_PADDR[5]), .Y(\CONFIG_reg_o_2_6_1_1[5] ));
    SLE \xhdl1.GEN_BITS[20].REG_GEN.CONFIG_reg[20][4]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[4]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[20]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[20][4] ));
    SLE \xhdl1.GEN_BITS[2].APB_32.edge_neg[2]  (.D(N_119), .CLK(
        FCCC_0_GL1), .EN(N_56), .ALn(MSS_RESET_N_F2M_c), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\edge_neg[2] ));
    CFG2 #( .INIT(4'hB) )  edge_both_2_sqmuxa_7_i (.A(edge_N_5_mux), 
        .B(\CONFIG_reg[21][3] ), .Y(N_198));
    CFG4 #( .INIT(16'hAC0F) )  
        \xhdl1.GEN_BITS[28].REG_GEN.CONFIG_reg[28]_RNIUIKA2[0]  (.A(
        \CONFIG_reg[12][0] ), .B(\CONFIG_reg[28][0] ), .C(
        \CONFIG_reg_o_2_6_1[0] ), .D(CoreAPB3_0_APBmslave2_PADDR[5]), 
        .Y(N_4699));
    SLE \xhdl1.GEN_BITS[31].REG_GEN.CONFIG_reg[31][4]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[4]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[31]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[31][4] ));
    SLE \xhdl1.GEN_BITS[0].APB_32.edge_pos[0]  (.D(N_109), .CLK(
        FCCC_0_GL1), .EN(N_74), .ALn(MSS_RESET_N_F2M_c), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\edge_pos[0] ));
    SLE \xhdl1.GEN_BITS[2].APB_32.GPOUT_reg[2]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[2]), .CLK(FCCC_0_GL1), .EN(
        GPOUT_reg_0_sqmuxa), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        GPOUT_reg_2));
    SLE \xhdl1.GEN_BITS[1].gpin1[1]  (.D(GPIO_IN_c[1]), .CLK(
        FCCC_0_GL1), .EN(VCC_net_1), .ALn(MSS_RESET_N_F2M_c), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\gpin1[1] ));
    SLE \xhdl1.GEN_BITS[0].APB_32.INTR_reg[0]  (.D(\INTR_reg_9[0] ), 
        .CLK(FCCC_0_GL1), .EN(VCC_net_1), .ALn(MSS_RESET_N_F2M_c), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(INTR_reg_0));
    CFG4 #( .INIT(16'hC5CA) )  
        \xhdl1.GEN_BITS[3].REG_INT.un34_intr_u_bm  (.A(gpin3_3), .B(
        N_4549), .C(\CONFIG_reg[3][6] ), .D(\CONFIG_reg[3][5] ), .Y(
        un34_intr_u_bm));
    SLE \xhdl1.GEN_BITS[2].REG_GEN.CONFIG_reg[2][5]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[5]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[2]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[2][5] ));
    CFG4 #( .INIT(16'h1000) )  
        \xhdl1.GEN_BITS[24].REG_GEN.CONFIG_reg[24]2_0_a4_0_a2  (.A(
        CoreAPB3_0_APBmslave2_PADDR[3]), .B(
        CoreAPB3_0_APBmslave2_PADDR[2]), .C(N_598), .D(N_610), .Y(
        \CONFIG_reg[24]2 ));
    CFG3 #( .INIT(8'hFB) )  edge_both_2_sqmuxa_14_i_0 (.A(edge_N_5_mux)
        , .B(\CONFIG_reg[1][3] ), .C(N_142_i), .Y(N_82));
    CFG4 #( .INIT(16'hC5CA) )  
        \xhdl1.GEN_BITS[4].APB_32.INTR_reg_61_0_m2[4]  (.A(\gpin3[4] ), 
        .B(N_172), .C(\CONFIG_reg[4][6] ), .D(\CONFIG_reg[4][5] ), .Y(
        N_179));
    CFG4 #( .INIT(16'hC480) )  
        \xhdl1.GEN_BITS[6].APB_32.INTR_reg_87_0_0_0_tz[6]  (.A(
        \CONFIG_reg[6][7] ), .B(\CONFIG_reg[6][3] ), .C(
        \INTR_reg_87_0_0_0_tz_1[6] ), .D(N_5939), .Y(
        \INTR_reg_87_0_0_0_tz[6] ));
    SLE \xhdl1.GEN_BITS[28].REG_GEN.CONFIG_reg[28][5]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[5]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[28]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[28][5] ));
    SLE \xhdl1.GEN_BITS[22].REG_GEN.CONFIG_reg[22][4]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[4]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[22]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[22][4] ));
    CFG4 #( .INIT(16'hAA08) )  
        \xhdl1.GEN_BITS[1].APB_32.edge_pos_23_iv_i_0[1]  (.A(
        \CONFIG_reg[1][3] ), .B(\edge_pos[1] ), .C(
        CoreAPB3_0_APBmslave2_PWDATA[1]), .D(N_400), .Y(N_107));
    CFG4 #( .INIT(16'hA9FF) )  
        \xhdl1.GEN_BITS[14].APB_32.INTR_reg_191_0_o2_0_0[14]  (.A(
        \CONFIG_reg[14][7] ), .B(\CONFIG_reg[14][6] ), .C(
        \CONFIG_reg[14][5] ), .D(\CONFIG_reg[14][3] ), .Y(
        \INTR_reg_191_0_o2_0[14] ));
    CFG4 #( .INIT(16'h0F35) )  
        \xhdl1.GEN_BITS[16].REG_GEN.CONFIG_reg[16]_RNI44E11[2]  (.A(
        \CONFIG_reg[0][2] ), .B(\CONFIG_reg[16][2] ), .C(
        CoreAPB3_0_APBmslave2_PADDR[6]), .D(
        CoreAPB3_0_APBmslave2_PADDR[5]), .Y(\CONFIG_reg_o_2_3_1_1[2] ));
    CFG4 #( .INIT(16'h0A33) )  
        \xhdl1.GEN_BITS[14].APB_32.INTR_reg_191_0[14]  (.A(INTR_reg_14)
        , .B(\INTR_reg_191_0_o2_1[14] ), .C(
        CoreAPB3_0_APBmslave2_PWDATA[14]), .D(edge_N_5_mux), .Y(
        \INTR_reg_191[14] ));
    SLE \xhdl1.GEN_BITS[6].APB_32.edge_both[6]  (.D(N_22_i_0), .CLK(
        FCCC_0_GL1), .EN(N_78), .ALn(MSS_RESET_N_F2M_c), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\edge_both[6] ));
    SLE \xhdl1.GEN_BITS[5].REG_GEN.CONFIG_reg[5][4]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[4]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[5]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[5][4] ));
    CFG4 #( .INIT(16'hAC0F) )  
        \xhdl1.GEN_BITS[14].REG_GEN.CONFIG_reg[14]_RNIC4Q82[4]  (.A(
        \CONFIG_reg[14][4] ), .B(\CONFIG_reg[30][4] ), .C(
        \CONFIG_reg_o_2_13_1_1[4] ), .D(CoreAPB3_0_APBmslave2_PADDR[5])
        , .Y(N_4759));
    CFG2 #( .INIT(4'h2) )  edge_pos_2_sqmuxa_4_i_a2 (.A(\gpin2[4] ), 
        .B(\gpin3[4] ), .Y(N_398));
    CFG4 #( .INIT(16'hAA08) )  
        \xhdl1.GEN_BITS[2].APB_32.edge_both_37_iv_i_0[2]  (.A(
        \CONFIG_reg[2][3] ), .B(\edge_both[2] ), .C(
        CoreAPB3_0_APBmslave2_PWDATA[2]), .D(N_144_i), .Y(N_93));
    CFG3 #( .INIT(8'hFB) )  edge_neg_2_sqmuxa_10_i_0 (.A(edge_N_5_mux), 
        .B(\CONFIG_reg[2][3] ), .C(N_395), .Y(N_56));
    SLE \xhdl1.GEN_BITS[13].APB_32.INTR_reg[13]  (.D(
        \INTR_reg_178[13] ), .CLK(FCCC_0_GL1), .EN(VCC_net_1), .ALn(
        MSS_RESET_N_F2M_c), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(INTR_reg_13));
    SLE \xhdl1.GEN_BITS[0].APB_32.edge_neg[0]  (.D(N_123), .CLK(
        FCCC_0_GL1), .EN(N_52), .ALn(MSS_RESET_N_F2M_c), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\edge_neg[0] ));
    SLE \xhdl1.GEN_BITS[13].REG_GEN.CONFIG_reg[13][2]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[2]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[13]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[13][2] ));
    CFG4 #( .INIT(16'h8000) )  
        \xhdl1.GEN_BITS[15].REG_GEN.CONFIG_reg[15]2_0_a4_0_a2  (.A(
        CoreAPB3_0_APBmslave2_PADDR[3]), .B(
        CoreAPB3_0_APBmslave2_PADDR[2]), .C(N_604), .D(N_605), .Y(
        \CONFIG_reg[15]2 ));
    SLE \xhdl1.GEN_BITS[16].REG_GEN.CONFIG_reg[16][5]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[5]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[16]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[16][5] ));
    SLE \xhdl1.GEN_BITS[25].REG_GEN.CONFIG_reg[25][7]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[7]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[25]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[25][7] ));
    CFG4 #( .INIT(16'hA9FF) )  
        \xhdl1.GEN_BITS[10].APB_32.INTR_reg_139_0_o2_0_0[10]  (.A(
        \CONFIG_reg[10][7] ), .B(\CONFIG_reg[10][6] ), .C(
        \CONFIG_reg[10][5] ), .D(\CONFIG_reg[10][3] ), .Y(
        \INTR_reg_139_0_o2_0[10] ));
    SLE \xhdl1.GEN_BITS[4].REG_GEN.CONFIG_reg[4][4]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[4]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[4]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[4][4] ));
    CFG4 #( .INIT(16'hAC0F) )  
        \xhdl1.GEN_BITS[24].REG_GEN.CONFIG_reg[24]_RNI2KQ22[0]  (.A(
        \CONFIG_reg[8][0] ), .B(\CONFIG_reg[24][0] ), .C(
        \CONFIG_reg_o_2_3_1[0] ), .D(CoreAPB3_0_APBmslave2_PADDR[5]), 
        .Y(N_4675));
    CFG4 #( .INIT(16'h4000) )  
        \xhdl1.GEN_BITS[29].REG_GEN.CONFIG_reg[29]2_0_a4_0_a2  (.A(
        CoreAPB3_0_APBmslave2_PADDR[3]), .B(
        CoreAPB3_0_APBmslave2_PADDR[2]), .C(N_598), .D(N_605), .Y(
        \CONFIG_reg[29]2 ));
    SLE \xhdl1.GEN_BITS[5].APB_32.GPOUT_reg[5]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[5]), .CLK(FCCC_0_GL1), .EN(
        GPOUT_reg_0_sqmuxa), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        GPOUT_reg_5));
    CFG2 #( .INIT(4'hB) )  edge_both_2_sqmuxa_6_i (.A(edge_N_5_mux), 
        .B(\CONFIG_reg[22][3] ), .Y(N_200));
    SLE \xhdl1.GEN_BITS[1].REG_GEN.CONFIG_reg[1][5]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[5]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[1]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[1][5] ));
    SLE \xhdl1.GEN_BITS[18].APB_32.GPOUT_reg[18]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[18]), .CLK(FCCC_0_GL1), .EN(
        GPOUT_reg_0_sqmuxa), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        GPOUT_reg_18));
    CFG4 #( .INIT(16'h0F35) )  
        \xhdl1.GEN_BITS[21].REG_GEN.CONFIG_reg[21]_RNIC6H61[5]  (.A(
        \CONFIG_reg[5][5] ), .B(\CONFIG_reg[21][5] ), .C(
        CoreAPB3_0_APBmslave2_PADDR[6]), .D(
        CoreAPB3_0_APBmslave2_PADDR[5]), .Y(\CONFIG_reg_o_2_21_1_1[5] )
        );
    CFG4 #( .INIT(16'h0F35) )  
        \xhdl1.GEN_BITS[7].REG_GEN.CONFIG_reg[7]_RNIIUKB1[4]  (.A(
        \CONFIG_reg[7][4] ), .B(\CONFIG_reg[23][4] ), .C(
        CoreAPB3_0_APBmslave2_PADDR[6]), .D(
        CoreAPB3_0_APBmslave2_PADDR[5]), .Y(\CONFIG_reg_o_2_28_1_1[4] )
        );
    SLE \xhdl1.GEN_BITS[14].REG_GEN.CONFIG_reg[14][3]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[3]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[14]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[14][3] ));
    SLE \xhdl1.GEN_BITS[0].REG_GEN.CONFIG_reg[0][1]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[1]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[0]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[0]_1 ));
    SLE \xhdl1.GEN_BITS[30].REG_GEN.CONFIG_reg[30][0]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[0]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[30]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[30][0] ));
    SLE \xhdl1.GEN_BITS[25].APB_32.GPOUT_reg[25]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[25]), .CLK(FCCC_0_GL1), .EN(
        GPOUT_reg_0_sqmuxa), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        GPOUT_reg_25));
    SLE \xhdl1.GEN_BITS[22].REG_GEN.CONFIG_reg[22][5]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[5]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[22]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[22][5] ));
    CFG4 #( .INIT(16'hF2F3) )  
        \xhdl1.GEN_BITS[28].APB_32.INTR_reg_373_0_o2_1_0[28]  (.A(
        \CONFIG_reg[28][6] ), .B(\edge_pos[28] ), .C(
        \INTR_reg_373_0_o2_0[28] ), .D(\CONFIG_reg[28][5] ), .Y(
        \INTR_reg_373_0_o2_1[28] ));
    CFG4 #( .INIT(16'h0A33) )  
        \xhdl1.GEN_BITS[10].APB_32.INTR_reg_139_0[10]  (.A(INTR_reg_10)
        , .B(\INTR_reg_139_0_o2_1[10] ), .C(
        CoreAPB3_0_APBmslave2_PWDATA[10]), .D(edge_N_5_mux), .Y(
        \INTR_reg_139[10] ));
    SLE \xhdl1.GEN_BITS[31].REG_GEN.CONFIG_reg[31][5]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[5]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[31]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[31][5] ));
    CFG4 #( .INIT(16'hC5CA) )  
        \xhdl1.GEN_BITS[5].APB_32.INTR_reg_74_0_0_m2[5]  (.A(gpin3_5), 
        .B(N_171), .C(\CONFIG_reg[5][6] ), .D(\CONFIG_reg[5][5] ), .Y(
        N_5940));
    CFG4 #( .INIT(16'hAC0F) )  
        \xhdl1.GEN_BITS[9].REG_GEN.CONFIG_reg[9]_RNI27V72[6]  (.A(
        \CONFIG_reg[9][6] ), .B(\CONFIG_reg[25][6] ), .C(
        \CONFIG_reg_o_2_18_1_1[6] ), .D(CoreAPB3_0_APBmslave2_PADDR[5])
        , .Y(N_4801));
    SLE \xhdl1.GEN_BITS[5].REG_GEN.CONFIG_reg[5][6]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[6]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[5]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[5][6] ));
    CFG4 #( .INIT(16'hAC0F) )  
        \xhdl1.GEN_BITS[28].REG_GEN.CONFIG_reg[28]_RNI6RKA2[2]  (.A(
        \CONFIG_reg[12][2] ), .B(\CONFIG_reg[28][2] ), .C(
        \CONFIG_reg_o_2_6_1_1[2] ), .D(CoreAPB3_0_APBmslave2_PADDR[5]), 
        .Y(N_4701));
    SLE \xhdl1.GEN_BITS[7].REG_GEN.CONFIG_reg[7][4]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[4]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[7]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[7][4] ));
    CFG4 #( .INIT(16'h0F35) )  
        \xhdl1.GEN_BITS[4].REG_GEN.CONFIG_reg[4]_RNICDV31[7]  (.A(
        \CONFIG_reg[4][7] ), .B(\CONFIG_reg[20][7] ), .C(
        CoreAPB3_0_APBmslave2_PADDR[6]), .D(
        CoreAPB3_0_APBmslave2_PADDR[5]), .Y(\CONFIG_reg_o_2_6_1_1[7] ));
    SLE \xhdl1.GEN_BITS[25].REG_GEN.CONFIG_reg[25][1]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[1]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[25]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[25][1] ));
    CFG4 #( .INIT(16'hA9FF) )  
        \xhdl1.GEN_BITS[24].APB_32.INTR_reg_321_0_o2_0_0[24]  (.A(
        \CONFIG_reg[24][7] ), .B(\CONFIG_reg[24][6] ), .C(
        \CONFIG_reg[24][5] ), .D(\CONFIG_reg[24][3] ), .Y(
        \INTR_reg_321_0_o2_0[24] ));
    SLE \xhdl1.GEN_BITS[10].REG_GEN.CONFIG_reg[10][5]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[5]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[10]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[10][5] ));
    SLE \xhdl1.GEN_BITS[17].REG_GEN.CONFIG_reg[17][2]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[2]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[17]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[17][2] ));
    SLE \xhdl1.GEN_BITS[23].REG_GEN.CONFIG_reg[23][4]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[4]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[23]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[23][4] ));
    SLE \xhdl1.GEN_BITS[18].REG_GEN.CONFIG_reg[18][3]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[3]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[18]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[18][3] ));
    CFG4 #( .INIT(16'hAC0F) )  
        \xhdl1.GEN_BITS[15].REG_GEN.CONFIG_reg[15]_RNI4FN32[0]  (.A(
        \CONFIG_reg[15][0] ), .B(\CONFIG_reg[31][0] ), .C(
        \CONFIG_reg_o_2_28_1_1[0] ), .D(CoreAPB3_0_APBmslave2_PADDR[5])
        , .Y(N_4875));
    CFG3 #( .INIT(8'h20) )  
        \xhdl1.GEN_BITS[23].APB_32.edge_both_RNO[23]  (.A(
        \CONFIG_reg[23][3] ), .B(CoreAPB3_0_APBmslave2_PWDATA[23]), .C(
        \edge_neg[23] ), .Y(N_96_i_0));
    SLE \xhdl1.GEN_BITS[4].REG_GEN.CONFIG_reg[4][6]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[6]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[4]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[4][6] ));
    SLE \xhdl1.GEN_BITS[26].REG_GEN.CONFIG_reg[26][6]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[6]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[26]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[26][6] ));
    SLE \xhdl1.GEN_BITS[29].APB_32.INTR_reg[29]  (.D(
        \INTR_reg_386[29] ), .CLK(FCCC_0_GL1), .EN(VCC_net_1), .ALn(
        MSS_RESET_N_F2M_c), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(INTR_reg_29));
    SLE \xhdl1.GEN_BITS[10].REG_GEN.CONFIG_reg[10][2]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[2]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[10]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[10][2] ));
    SLE \xhdl1.GEN_BITS[25].APB_32.INTR_reg[25]  (.D(
        \INTR_reg_334[25] ), .CLK(FCCC_0_GL1), .EN(VCC_net_1), .ALn(
        MSS_RESET_N_F2M_c), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(INTR_reg_25));
    CFG4 #( .INIT(16'hA9FF) )  
        \xhdl1.GEN_BITS[13].APB_32.INTR_reg_178_0_o2_0_0[13]  (.A(
        \CONFIG_reg[13][7] ), .B(\CONFIG_reg[13][6] ), .C(
        \CONFIG_reg[13][5] ), .D(\CONFIG_reg[13][3] ), .Y(
        \INTR_reg_178_0_o2_0[13] ));
    SLE \xhdl1.GEN_BITS[28].REG_GEN.CONFIG_reg[28][1]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[1]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[28]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[28][1] ));
    SLE \xhdl1.GEN_BITS[6].APB_32.edge_neg[6]  (.D(N_113), .CLK(
        FCCC_0_GL1), .EN(N_62), .ALn(MSS_RESET_N_F2M_c), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\edge_neg[6] ));
    SLE \xhdl1.GEN_BITS[20].REG_GEN.CONFIG_reg[20][7]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[7]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[20]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[20][7] ));
    CFG4 #( .INIT(16'h4000) )  
        \xhdl1.GEN_BITS[17].REG_GEN.CONFIG_reg[17]2_0_a4_0_a2  (.A(
        CoreAPB3_0_APBmslave2_PADDR[3]), .B(
        CoreAPB3_0_APBmslave2_PADDR[2]), .C(N_598), .D(N_606), .Y(
        \CONFIG_reg[17]2 ));
    SLE \xhdl1.GEN_BITS[30].REG_GEN.CONFIG_reg[30][2]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[2]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[30]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[30][2] ));
    SLE \xhdl1.GEN_BITS[26].APB_32.INTR_reg[26]  (.D(
        \INTR_reg_347[26] ), .CLK(FCCC_0_GL1), .EN(VCC_net_1), .ALn(
        MSS_RESET_N_F2M_c), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(INTR_reg_26));
    SLE \xhdl1.GEN_BITS[27].APB_32.edge_both[27]  (.D(N_5912_i_0), 
        .CLK(FCCC_0_GL1), .EN(N_161), .ALn(MSS_RESET_N_F2M_c), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\edge_neg[27] ));
    CFG2 #( .INIT(4'h6) )  edge_both_2_sqmuxa_11_i_x2 (.A(\gpin2[4] ), 
        .B(\gpin3[4] ), .Y(N_143_i));
    SLE \xhdl1.GEN_BITS[27].REG_GEN.CONFIG_reg[27][7]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[7]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[27]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[27][7] ));
    SLE \xhdl1.GEN_BITS[22].REG_GEN.CONFIG_reg[22][3]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[3]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[22]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[22][3] ));
    SLE \xhdl1.GEN_BITS[25].APB_32.edge_both[25]  (.D(N_5911_i_0), 
        .CLK(FCCC_0_GL1), .EN(N_157), .ALn(MSS_RESET_N_F2M_c), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\edge_neg[25] ));
    SLE \xhdl1.GEN_BITS[25].REG_GEN.CONFIG_reg[25][6]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[6]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[25]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[25][6] ));
    CFG4 #( .INIT(16'hC480) )  
        \xhdl1.GEN_BITS[0].APB_32.INTR_reg_9_0_0_0_tz[0]  (.A(
        \CONFIG_reg[0][7] ), .B(\CONFIG_reg[0][3] ), .C(
        \INTR_reg_9_0_0_0_tz_1[0] ), .D(N_5941), .Y(
        \INTR_reg_9_0_0_0_tz[0] ));
    CFG2 #( .INIT(4'h2) )  edge_pos_2_sqmuxa_i_a2 (.A(\gpin2[0] ), .B(
        gpin3_0), .Y(N_402));
    SLE \xhdl1.GEN_BITS[7].REG_GEN.CONFIG_reg[7][6]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[6]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[7]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[7][6] ));
    CFG4 #( .INIT(16'h4000) )  
        \xhdl1.GEN_BITS[1].REG_GEN.CONFIG_reg[1]2_0_a4_0_a2  (.A(
        CoreAPB3_0_APBmslave2_PADDR[3]), .B(
        CoreAPB3_0_APBmslave2_PADDR[2]), .C(N_604), .D(N_606), .Y(
        \CONFIG_reg[1]2 ));
    CFG4 #( .INIT(16'hA9FF) )  
        \xhdl1.GEN_BITS[28].APB_32.INTR_reg_373_0_o2_0_0[28]  (.A(
        \CONFIG_reg[28][7] ), .B(\CONFIG_reg[28][6] ), .C(
        \CONFIG_reg[28][5] ), .D(\CONFIG_reg[28][3] ), .Y(
        \INTR_reg_373_0_o2_0[28] ));
    CFG4 #( .INIT(16'hAC0F) )  
        \xhdl1.GEN_BITS[11].REG_GEN.CONFIG_reg[11]_RNIKPD72[3]  (.A(
        \CONFIG_reg[11][3] ), .B(\CONFIG_reg[27][3] ), .C(
        \CONFIG_reg_o_2_25_1_1[3] ), .D(CoreAPB3_0_APBmslave2_PADDR[5])
        , .Y(N_4854));
    SLE \xhdl1.GEN_BITS[4].APB_32.GPOUT_reg[4]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[4]), .CLK(FCCC_0_GL1), .EN(
        GPOUT_reg_0_sqmuxa), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        GPOUT_reg_4));
    CFG3 #( .INIT(8'h01) )  \xhdl1.GEN_m3_e_1  (.A(
        CoreAPB3_0_APBmslave2_PADDR[7]), .B(
        FIC_MSS_0_FIC_0_APB_MASTER_PADDR_2), .C(
        FIC_MSS_0_FIC_0_APB_MASTER_PADDR_0), .Y(GEN_m3_e_1));
    SLE \xhdl1.GEN_BITS[19].REG_GEN.CONFIG_reg[19][7]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[7]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[19]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[19][7] ));
    SLE \xhdl1.GEN_BITS[18].REG_GEN.CONFIG_reg[18][6]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[6]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[18]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[18][6] ));
    CFG2 #( .INIT(4'hE) )  
        \xhdl1.GEN_BITS[0].APB_32.un5_PRDATA_o_0_a2_0_o2  (.A(N_245), 
        .B(un5_PRDATA_o_0_a2_0_o2_out), .Y(N_247));
    CFG4 #( .INIT(16'hAC0F) )  
        \xhdl1.GEN_BITS[29].REG_GEN.CONFIG_reg[29]_RNIAII52[1]  (.A(
        \CONFIG_reg[13][1] ), .B(\CONFIG_reg[29][1] ), .C(
        \CONFIG_reg_o_2_21_1_1[1] ), .D(CoreAPB3_0_APBmslave2_PADDR[5])
        , .Y(N_4820));
    SLE \xhdl1.GEN_BITS[12].APB_32.INTR_reg[12]  (.D(
        \INTR_reg_165[12] ), .CLK(FCCC_0_GL1), .EN(VCC_net_1), .ALn(
        MSS_RESET_N_F2M_c), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(INTR_reg_12));
    CFG3 #( .INIT(8'hB8) )  
        \xhdl1.GEN_BITS[5].APB_32.INTR_reg_74_0_m2_0_i_m2[5]  (.A(
        \edge_neg[5] ), .B(\CONFIG_reg[5][5] ), .C(\edge_pos[5] ), .Y(
        N_171));
    SLE \xhdl1.GEN_BITS[13].REG_GEN.CONFIG_reg[13][1]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[1]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[13]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[13][1] ));
    CFG3 #( .INIT(8'hFB) )  edge_both_2_sqmuxa_23_i_0 (.A(edge_N_5_mux)
        , .B(\CONFIG_reg[5][3] ), .C(N_139_i), .Y(N_76));
    SLE \xhdl1.GEN_BITS[28].REG_GEN.CONFIG_reg[28][7]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[7]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[28]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[28][7] ));
    CFG2 #( .INIT(4'h6) )  edge_both_2_sqmuxa_23_i_x2 (.A(\gpin2[5] ), 
        .B(gpin3_5), .Y(N_139_i));
    CFG4 #( .INIT(16'h0F35) )  
        \xhdl1.GEN_BITS[16].REG_GEN.CONFIG_reg[16]_RNIEEE11[7]  (.A(
        \CONFIG_reg[0][7] ), .B(\CONFIG_reg[16][7] ), .C(
        CoreAPB3_0_APBmslave2_PADDR[6]), .D(
        CoreAPB3_0_APBmslave2_PADDR[5]), .Y(\CONFIG_reg_o_2_3_1_1[7] ));
    SLE \xhdl1.GEN_BITS[5].REG_GEN.CONFIG_reg[5][0]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[0]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[5]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[5][0] ));
    CFG4 #( .INIT(16'h0A33) )  
        \xhdl1.GEN_BITS[21].APB_32.INTR_reg_282_0[21]  (.A(INTR_reg_21)
        , .B(\INTR_reg_282_0_o2_1[21] ), .C(
        CoreAPB3_0_APBmslave2_PWDATA[21]), .D(edge_N_5_mux), .Y(
        \INTR_reg_282[21] ));
    CFG2 #( .INIT(4'h8) )  
        \xhdl1.GEN_BITS[0].REG_GPOUT.un5_GPIO_OUT_i  (.A(GPOUT_reg_0), 
        .B(\CONFIG_reg[0][0] ), .Y(GPIO_OUT_net_2[0]));
    CFG4 #( .INIT(16'h2000) )  
        \xhdl1.GEN_BITS[30].REG_GEN.CONFIG_reg[30]2_0_a4_0_a2  (.A(
        CoreAPB3_0_APBmslave2_PADDR[3]), .B(
        CoreAPB3_0_APBmslave2_PADDR[2]), .C(N_598), .D(N_605), .Y(
        \CONFIG_reg[30]2 ));
    SLE \xhdl1.GEN_BITS[31].APB_32.INTR_reg[31]  (.D(
        \INTR_reg_412[31] ), .CLK(FCCC_0_GL1), .EN(VCC_net_1), .ALn(
        MSS_RESET_N_F2M_c), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(INTR_reg_31));
    SLE \xhdl1.GEN_BITS[13].REG_GEN.CONFIG_reg[13][7]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[7]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[13]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[13][7] ));
    GND GND (.Y(GND_net_1));
    SLE \xhdl1.GEN_BITS[31].APB_32.GPOUT_reg[31]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[31]), .CLK(FCCC_0_GL1), .EN(
        GPOUT_reg_0_sqmuxa), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        GPOUT_reg_31));
    SLE \xhdl1.GEN_BITS[20].REG_GEN.CONFIG_reg[20][6]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[6]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[20]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[20][6] ));
    CFG3 #( .INIT(8'hB8) )  
        \xhdl1.GEN_BITS[1].APB_32.INTR_reg_22_0_m2_0[1]  (.A(
        \edge_neg[1] ), .B(\CONFIG_reg[1][5] ), .C(\edge_pos[1] ), .Y(
        N_174));
    CFG4 #( .INIT(16'hAC0F) )  
        \xhdl1.GEN_BITS[24].REG_GEN.CONFIG_reg[24]_RNIQCR22[6]  (.A(
        \CONFIG_reg[8][6] ), .B(\CONFIG_reg[24][6] ), .C(
        \CONFIG_reg_o_2_3_1_1[6] ), .D(CoreAPB3_0_APBmslave2_PADDR[5]), 
        .Y(N_4681));
    CFG4 #( .INIT(16'h8000) )  
        \xhdl1.GEN_BITS[16].REG_GEN.CONFIG_reg[16]2_0_a4_0_a2_1  (.A(
        CoreAPB3_0_APBmslave2_PADDR[6]), .B(wen_0), .C(GEN_m3_e_1), .D(
        iPSELS_2[5]), .Y(N_598));
    SLE \xhdl1.GEN_BITS[22].REG_GEN.CONFIG_reg[22][1]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[1]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[22]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[22][1] ));
    CFG4 #( .INIT(16'h0F35) )  
        \xhdl1.GEN_BITS[17].REG_GEN.CONFIG_reg[17]_RNIC50K1[4]  (.A(
        \CONFIG_reg[1][4] ), .B(\CONFIG_reg[17][4] ), .C(
        CoreAPB3_0_APBmslave2_PADDR[6]), .D(
        CoreAPB3_0_APBmslave2_PADDR[5]), .Y(\CONFIG_reg_o_2_18_1[4] ));
    SLE \xhdl1.GEN_BITS[26].APB_32.GPOUT_reg[26]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[26]), .CLK(FCCC_0_GL1), .EN(
        GPOUT_reg_0_sqmuxa), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        GPOUT_reg_26));
    SLE \xhdl1.GEN_BITS[4].REG_GEN.CONFIG_reg[4][0]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[0]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[4]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[4][0] ));
    CFG4 #( .INIT(16'hA9FF) )  
        \xhdl1.GEN_BITS[21].APB_32.INTR_reg_282_0_o2_0_0[21]  (.A(
        \CONFIG_reg[21][7] ), .B(\CONFIG_reg[21][6] ), .C(
        \CONFIG_reg[21][5] ), .D(\CONFIG_reg[21][3] ), .Y(
        \INTR_reg_282_0_o2_0[21] ));
    CFG4 #( .INIT(16'hA9FF) )  
        \xhdl1.GEN_BITS[19].APB_32.INTR_reg_256_0_o2_0_0[19]  (.A(
        \CONFIG_reg[19][7] ), .B(\CONFIG_reg[19][6] ), .C(
        \CONFIG_reg[19][5] ), .D(\CONFIG_reg[19][3] ), .Y(
        \INTR_reg_256_0_o2_0[19] ));
    SLE \xhdl1.GEN_BITS[11].APB_32.edge_both[11]  (.D(
        \edge_neg_163[11] ), .CLK(FCCC_0_GL1), .EN(N_186), .ALn(
        MSS_RESET_N_F2M_c), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\edge_neg[11] ));
    CFG4 #( .INIT(16'hAC0F) )  
        \xhdl1.GEN_BITS[14].REG_GEN.CONFIG_reg[14]_RNI80Q82[3]  (.A(
        \CONFIG_reg[14][3] ), .B(\CONFIG_reg[30][3] ), .C(
        \CONFIG_reg_o_2_13_1_1[3] ), .D(CoreAPB3_0_APBmslave2_PADDR[5])
        , .Y(N_4758));
    CFG4 #( .INIT(16'h0F35) )  
        \xhdl1.GEN_BITS[21].REG_GEN.CONFIG_reg[21]_RNIGAH61[7]  (.A(
        \CONFIG_reg[5][7] ), .B(\CONFIG_reg[21][7] ), .C(
        CoreAPB3_0_APBmslave2_PADDR[6]), .D(
        CoreAPB3_0_APBmslave2_PADDR[5]), .Y(\CONFIG_reg_o_2_21_1_1[7] )
        );
    SLE \xhdl1.GEN_BITS[22].REG_GEN.CONFIG_reg[22][6]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[6]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[22]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[22][6] ));
    SLE \xhdl1.GEN_BITS[2].REG_GEN.CONFIG_reg[2][3]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[3]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[2]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[2][3] ));
    SLE \xhdl1.GEN_BITS[13].REG_GEN.CONFIG_reg[13][4]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[4]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[13]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[13][4] ));
    CFG4 #( .INIT(16'h1000) )  
        \xhdl1.GEN_BITS[20].REG_GEN.CONFIG_reg[20]2_0_a4_0_a2  (.A(
        CoreAPB3_0_APBmslave2_PADDR[3]), .B(
        CoreAPB3_0_APBmslave2_PADDR[2]), .C(N_598), .D(N_603), .Y(
        \CONFIG_reg[20]2 ));
    SLE \xhdl1.GEN_BITS[12].REG_GEN.CONFIG_reg[12][6]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[6]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[12]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[12][6] ));
    SLE \xhdl1.GEN_BITS[31].REG_GEN.CONFIG_reg[31][1]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[1]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[31]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[31][1] ));
    CFG4 #( .INIT(16'h0A33) )  
        \xhdl1.GEN_BITS[28].APB_32.INTR_reg_373_0[28]  (.A(INTR_reg_28)
        , .B(\INTR_reg_373_0_o2_1[28] ), .C(
        CoreAPB3_0_APBmslave2_PWDATA[28]), .D(edge_N_5_mux), .Y(
        \INTR_reg_373[28] ));
    CFG4 #( .INIT(16'h0F35) )  
        \xhdl1.GEN_BITS[16].REG_GEN.CONFIG_reg[16]_RNI88E11[4]  (.A(
        \CONFIG_reg[0][4] ), .B(\CONFIG_reg[16][4] ), .C(
        CoreAPB3_0_APBmslave2_PADDR[6]), .D(
        CoreAPB3_0_APBmslave2_PADDR[5]), .Y(\CONFIG_reg_o_2_3_1[4] ));
    CFG4 #( .INIT(16'hAC0F) )  
        \xhdl1.GEN_BITS[14].REG_GEN.CONFIG_reg[14]_RNI4SP82[2]  (.A(
        \CONFIG_reg[14][2] ), .B(\CONFIG_reg[30][2] ), .C(
        \CONFIG_reg_o_2_13_1_1[2] ), .D(CoreAPB3_0_APBmslave2_PADDR[5])
        , .Y(N_4757));
    SLE \xhdl1.GEN_BITS[2].REG_GEN.CONFIG_reg[2][7]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[7]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[2]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[2][7] ));
    SLE \xhdl1.GEN_BITS[7].REG_GEN.CONFIG_reg[7][0]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[0]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[7]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[7][0] ));
    CFG4 #( .INIT(16'hF2F3) )  
        \xhdl1.GEN_BITS[11].APB_32.INTR_reg_152_0_o2_1_0[11]  (.A(
        \CONFIG_reg[11][6] ), .B(\edge_neg[11] ), .C(
        \INTR_reg_152_0_o2_0[11] ), .D(\CONFIG_reg[11][5] ), .Y(
        \INTR_reg_152_0_o2_1[11] ));
    CFG4 #( .INIT(16'h0F35) )  
        \xhdl1.GEN_BITS[17].REG_GEN.CONFIG_reg[17]_RNIIB0K1[7]  (.A(
        \CONFIG_reg[1][7] ), .B(\CONFIG_reg[17][7] ), .C(
        CoreAPB3_0_APBmslave2_PADDR[6]), .D(
        CoreAPB3_0_APBmslave2_PADDR[5]), .Y(\CONFIG_reg_o_2_18_1_1[7] )
        );
    SLE \xhdl1.GEN_BITS[22].REG_GEN.CONFIG_reg[22][2]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[2]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[22]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[22][2] ));
    SLE \xhdl1.GEN_BITS[28].REG_GEN.CONFIG_reg[28][2]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[2]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[28]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[28][2] ));
    SLE \xhdl1.GEN_BITS[27].REG_GEN.CONFIG_reg[27][0]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[0]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[27]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[27][0] ));
    CFG4 #( .INIT(16'h0A33) )  
        \xhdl1.GEN_BITS[17].APB_32.INTR_reg_230_0[17]  (.A(INTR_reg_17)
        , .B(\INTR_reg_230_0_o2_1[17] ), .C(
        CoreAPB3_0_APBmslave2_PWDATA[17]), .D(edge_N_5_mux), .Y(
        \INTR_reg_230[17] ));
    CFG4 #( .INIT(16'hF2F3) )  
        \xhdl1.GEN_BITS[24].APB_32.INTR_reg_321_0_o2_1_0[24]  (.A(
        \CONFIG_reg[24][6] ), .B(\edge_pos[24] ), .C(
        \INTR_reg_321_0_o2_0[24] ), .D(\CONFIG_reg[24][5] ), .Y(
        \INTR_reg_321_0_o2_1[24] ));
    CFG4 #( .INIT(16'h1000) )  
        \xhdl1.GEN_BITS[28].REG_GEN.CONFIG_reg[28]2_0_a4_0_a2  (.A(
        CoreAPB3_0_APBmslave2_PADDR[3]), .B(
        CoreAPB3_0_APBmslave2_PADDR[2]), .C(N_598), .D(N_605), .Y(
        \CONFIG_reg[28]2 ));
    CFG4 #( .INIT(16'h0A33) )  
        \xhdl1.GEN_BITS[16].APB_32.INTR_reg_217_0[16]  (.A(INTR_reg_16)
        , .B(\INTR_reg_217_0_o2_1[16] ), .C(
        CoreAPB3_0_APBmslave2_PWDATA[16]), .D(edge_N_5_mux), .Y(
        \INTR_reg_217[16] ));
    CFG4 #( .INIT(16'hA9FF) )  
        \xhdl1.GEN_BITS[15].APB_32.INTR_reg_204_0_o2_0_0[15]  (.A(
        \CONFIG_reg[15][7] ), .B(\CONFIG_reg[15][6] ), .C(
        \CONFIG_reg[15][5] ), .D(\CONFIG_reg[15][3] ), .Y(
        \INTR_reg_204_0_o2_0[15] ));
    SLE \xhdl1.GEN_BITS[26].REG_GEN.CONFIG_reg[26][5]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[5]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[26]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[26][5] ));
    SLE \xhdl1.GEN_BITS[28].REG_GEN.CONFIG_reg[28][4]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[4]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[28]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[28][4] ));
    SLE \xhdl1.GEN_BITS[28].APB_32.GPOUT_reg[28]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[28]), .CLK(FCCC_0_GL1), .EN(
        GPOUT_reg_0_sqmuxa), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        GPOUT_reg_28));
    CFG4 #( .INIT(16'hAA08) )  
        \xhdl1.GEN_BITS[0].APB_32.edge_pos_9_iv_i_0[0]  (.A(
        \CONFIG_reg[0][3] ), .B(\edge_pos[0] ), .C(
        CoreAPB3_0_APBmslave2_PWDATA[0]), .D(N_402), .Y(N_109));
    SLE \xhdl1.GEN_BITS[3].gpin1[3]  (.D(GPIO_IN_c[3]), .CLK(
        FCCC_0_GL1), .EN(VCC_net_1), .ALn(MSS_RESET_N_F2M_c), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\gpin1[3] ));
    SLE \xhdl1.GEN_BITS[19].REG_GEN.CONFIG_reg[19][2]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[2]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[19]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[19][2] ));
    CFG4 #( .INIT(16'h1000) )  
        \xhdl1.GEN_BITS[3].REG_INT.un34_intr_u_ns_1  (.A(
        \CONFIG_reg[3][6] ), .B(\CONFIG_reg[3][5] ), .C(\edge_both[3] )
        , .D(\CONFIG_reg[3][7] ), .Y(un34_intr_u_ns_1));
    SLE \xhdl1.GEN_BITS[0].REG_GEN.CONFIG_reg[0][2]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[2]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[0]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[0][2] ));
    SLE \xhdl1.GEN_BITS[9].REG_GEN.CONFIG_reg[9][4]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[4]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[9]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[9][4] ));
    CFG4 #( .INIT(16'h8000) )  
        \xhdl1.GEN_BITS[7].REG_GEN.CONFIG_reg[7]2_0_a4_0_a2  (.A(
        CoreAPB3_0_APBmslave2_PADDR[2]), .B(
        CoreAPB3_0_APBmslave2_PADDR[3]), .C(N_603), .D(N_604), .Y(
        \CONFIG_reg[7]2 ));
    SLE \xhdl1.GEN_BITS[2].gpin2[2]  (.D(\gpin1[2] ), .CLK(FCCC_0_GL1), 
        .EN(VCC_net_1), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(\gpin2[2] ));
    CFG2 #( .INIT(4'h8) )  
        \xhdl1.GEN_BITS[1].REG_GPOUT.un14_GPIO_OUT_i  (.A(GPOUT_reg_1), 
        .B(\CONFIG_reg[1][0] ), .Y(GPIO_OUT_net_2[1]));
    CFG2 #( .INIT(4'hB) )  edge_both_2_sqmuxa_9_i (.A(edge_N_5_mux), 
        .B(\CONFIG_reg[19][3] ), .Y(N_194));
    SLE \xhdl1.GEN_BITS[1].REG_GEN.CONFIG_reg[1][3]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[3]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[1]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[1][3] ));
    CFG4 #( .INIT(16'h0F35) )  
        \xhdl1.GEN_BITS[17].REG_GEN.CONFIG_reg[17]_RNI6VVJ1[1]  (.A(
        \CONFIG_reg[1]_1 ), .B(\CONFIG_reg[17][1] ), .C(
        CoreAPB3_0_APBmslave2_PADDR[6]), .D(
        CoreAPB3_0_APBmslave2_PADDR[5]), .Y(\CONFIG_reg_o_2_18_1_1[1] )
        );
    CFG2 #( .INIT(4'h4) )  edge_neg_2_sqmuxa_i_0_0_a2 (.A(\gpin2[6] ), 
        .B(gpin3_6), .Y(N_688));
    SLE \xhdl1.GEN_BITS[27].REG_GEN.CONFIG_reg[27][2]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[2]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[27]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[27][2] ));
    SLE \xhdl1.GEN_BITS[8].REG_GEN.CONFIG_reg[8][4]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[4]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[8]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[8][4] ));
    CFG4 #( .INIT(16'h0F35) )  
        \xhdl1.GEN_BITS[22].REG_GEN.CONFIG_reg[22]_RNIE1391[4]  (.A(
        \CONFIG_reg[6][4] ), .B(\CONFIG_reg[22][4] ), .C(
        CoreAPB3_0_APBmslave2_PADDR[6]), .D(
        CoreAPB3_0_APBmslave2_PADDR[5]), .Y(\CONFIG_reg_o_2_13_1_1[4] )
        );
    CFG4 #( .INIT(16'hF2F3) )  
        \xhdl1.GEN_BITS[23].APB_32.INTR_reg_308_0_o2_1_0[23]  (.A(
        \CONFIG_reg[23][6] ), .B(\edge_neg[23] ), .C(
        \INTR_reg_308_0_o2_0[23] ), .D(\CONFIG_reg[23][5] ), .Y(
        \INTR_reg_308_0_o2_1[23] ));
    SLE \xhdl1.GEN_BITS[1].REG_GEN.CONFIG_reg[1][7]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[7]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[1]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[1][7] ));
    CFG2 #( .INIT(4'h2) )  edge_pos_2_sqmuxa_2_i_0_0_a2 (.A(\gpin2[6] )
        , .B(gpin3_6), .Y(N_689));
    SLE \xhdl1.GEN_BITS[17].REG_GEN.CONFIG_reg[17][0]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[0]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[17]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[17][0] ));
    CFG4 #( .INIT(16'hF2F3) )  
        \xhdl1.GEN_BITS[10].APB_32.INTR_reg_139_0_o2_1_0[10]  (.A(
        \CONFIG_reg[10][6] ), .B(\edge_pos[10] ), .C(
        \INTR_reg_139_0_o2_0[10] ), .D(\CONFIG_reg[10][5] ), .Y(
        \INTR_reg_139_0_o2_1[10] ));
    SLE \xhdl1.GEN_BITS[30].REG_GEN.CONFIG_reg[30][1]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[1]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[30]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[30][1] ));
    CFG2 #( .INIT(4'h6) )  edge_both_2_sqmuxa_i_x2 (.A(\gpin2[2] ), .B(
        gpin3_2), .Y(N_144_i));
    SLE \xhdl1.GEN_BITS[1].APB_32.edge_neg[1]  (.D(N_121), .CLK(
        FCCC_0_GL1), .EN(N_54), .ALn(MSS_RESET_N_F2M_c), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\edge_neg[1] ));
    SLE \xhdl1.GEN_BITS[10].REG_GEN.CONFIG_reg[10][6]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[6]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[10]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[10][6] ));
    SLE \xhdl1.GEN_BITS[6].gpin2[6]  (.D(\gpin1[6] ), .CLK(FCCC_0_GL1), 
        .EN(VCC_net_1), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(\gpin2[6] ));
    SLE \xhdl1.GEN_BITS[12].REG_GEN.CONFIG_reg[12][1]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[1]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[12]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[12][1] ));
    CFG4 #( .INIT(16'h0F35) )  
        \xhdl1.GEN_BITS[20].REG_GEN.CONFIG_reg[20]_RNIUUU31[0]  (.A(
        \CONFIG_reg[4][0] ), .B(\CONFIG_reg[20][0] ), .C(
        CoreAPB3_0_APBmslave2_PADDR[6]), .D(
        CoreAPB3_0_APBmslave2_PADDR[5]), .Y(\CONFIG_reg_o_2_6_1[0] ));
    CFG4 #( .INIT(16'hAC0F) )  
        \xhdl1.GEN_BITS[24].REG_GEN.CONFIG_reg[24]_RNIUGR22[7]  (.A(
        \CONFIG_reg[8][7] ), .B(\CONFIG_reg[24][7] ), .C(
        \CONFIG_reg_o_2_3_1_1[7] ), .D(CoreAPB3_0_APBmslave2_PADDR[5]), 
        .Y(N_4682));
    CFG3 #( .INIT(8'hB8) )  
        \xhdl1.GEN_BITS[0].APB_32.INTR_reg_9_0_m2_0[0]  (.A(
        \edge_neg[0] ), .B(\CONFIG_reg[0][5] ), .C(\edge_pos[0] ), .Y(
        N_175));
    CFG3 #( .INIT(8'hFB) )  edge_pos_2_sqmuxa_4_i_0 (.A(edge_N_5_mux), 
        .B(\CONFIG_reg[4][3] ), .C(N_398), .Y(N_68));
    CFG3 #( .INIT(8'hB8) )  
        \xhdl1.GEN_BITS[4].APB_32.INTR_reg_61_0_m2_0[4]  (.A(
        \edge_neg[4] ), .B(\CONFIG_reg[4][5] ), .C(\edge_pos[4] ), .Y(
        N_172));
    CFG3 #( .INIT(8'h20) )  
        \xhdl1.GEN_BITS[7].APB_32.edge_both_RNO[7]  (.A(
        \CONFIG_reg[7][3] ), .B(CoreAPB3_0_APBmslave2_PWDATA[7]), .C(
        \edge_pos[7] ), .Y(N_83_i_0));
    CFG3 #( .INIT(8'hB8) )  
        \xhdl1.GEN_BITS[6].APB_32.INTR_reg_87_0_0_m2_0[6]  (.A(
        \edge_neg[6] ), .B(\CONFIG_reg[6][5] ), .C(\edge_pos[6] ), .Y(
        N_5938));
    CFG4 #( .INIT(16'hA9FF) )  
        \xhdl1.GEN_BITS[30].APB_32.INTR_reg_399_0_o2_0_0[30]  (.A(
        \CONFIG_reg[30][7] ), .B(\CONFIG_reg[30][6] ), .C(
        \CONFIG_reg[30][5] ), .D(\CONFIG_reg[30][3] ), .Y(
        \INTR_reg_399_0_o2_0[30] ));
    CFG2 #( .INIT(4'h2) )  edge_pos_2_sqmuxa_3_i_a2 (.A(\gpin2[5] ), 
        .B(gpin3_5), .Y(N_406));
    CFG2 #( .INIT(4'h6) )  
        \xhdl1.GEN_BITS[6].APB_32.edge_both_93_iv_i_0_i_x2[6]  (.A(
        \gpin2[6] ), .B(gpin3_6), .Y(N_252_i));
    CFG2 #( .INIT(4'hB) )  edge_both_2_sqmuxa_28_i (.A(edge_N_5_mux), 
        .B(\CONFIG_reg[27][3] ), .Y(N_161));
    CFG4 #( .INIT(16'h0F35) )  
        \xhdl1.GEN_BITS[2].REG_GEN.CONFIG_reg[2]_RNIM8I61[7]  (.A(
        \CONFIG_reg[2][7] ), .B(\CONFIG_reg[18][7] ), .C(
        CoreAPB3_0_APBmslave2_PADDR[6]), .D(
        CoreAPB3_0_APBmslave2_PADDR[5]), .Y(\CONFIG_reg_o_2_10_1_1[7] )
        );
    SLE \xhdl1.GEN_BITS[18].REG_GEN.CONFIG_reg[18][2]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[2]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[18]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[18][2] ));
    SLE \xhdl1.GEN_BITS[3].REG_GEN.CONFIG_reg[3][4]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[4]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[3]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[3][4] ));
    SLE \xhdl1.GEN_BITS[9].REG_GEN.CONFIG_reg[9][6]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[6]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[9]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[9][6] ));
    CFG2 #( .INIT(4'h2) )  edge_pos_2_sqmuxa_18_i_a2 (.A(\gpin2[3] ), 
        .B(gpin3_3), .Y(N_687));
    CFG2 #( .INIT(4'h8) )  
        \xhdl1.GEN_BITS[8].REG_GEN.CONFIG_reg[8]2_0_a4_0_a2  (.A(N_678)
        , .B(N_610), .Y(\CONFIG_reg[8]2 ));
    CFG4 #( .INIT(16'hAA08) )  
        \xhdl1.GEN_BITS[1].APB_32.edge_neg_23_iv_i_0[1]  (.A(
        \CONFIG_reg[1][3] ), .B(\edge_neg[1] ), .C(
        CoreAPB3_0_APBmslave2_PWDATA[1]), .D(N_399), .Y(N_121));
    CFG4 #( .INIT(16'hA9FF) )  
        \xhdl1.GEN_BITS[27].APB_32.INTR_reg_360_0_o2_0_0[27]  (.A(
        \CONFIG_reg[27][7] ), .B(\CONFIG_reg[27][6] ), .C(
        \CONFIG_reg[27][5] ), .D(\CONFIG_reg[27][3] ), .Y(
        \INTR_reg_360_0_o2_0[27] ));
    SLE \xhdl1.GEN_BITS[5].REG_GEN.CONFIG_reg[5][1]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[1]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[5]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[5]_1 ));
    CFG3 #( .INIT(8'hFB) )  edge_both_2_sqmuxa_i_0 (.A(edge_N_5_mux), 
        .B(\CONFIG_reg[2][3] ), .C(N_144_i), .Y(N_86));
    SLE \xhdl1.GEN_BITS[8].REG_GEN.CONFIG_reg[8][6]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[6]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[8]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[8][6] ));
    CFG4 #( .INIT(16'h8000) )  
        \xhdl1.GEN_BITS[27].REG_GEN.CONFIG_reg[27]2_0_a4_0_a2  (.A(
        CoreAPB3_0_APBmslave2_PADDR[3]), .B(
        CoreAPB3_0_APBmslave2_PADDR[2]), .C(N_598), .D(N_610), .Y(
        \CONFIG_reg[27]2 ));
    SLE \xhdl1.GEN_BITS[24].REG_GEN.CONFIG_reg[24][2]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[2]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[24]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[24][2] ));
    SLE \xhdl1.GEN_BITS[23].REG_GEN.CONFIG_reg[23][0]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[0]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[23]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[23][0] ));
    CFG3 #( .INIT(8'hFB) )  edge_neg_2_sqmuxa_11_i_0 (.A(edge_N_5_mux), 
        .B(\CONFIG_reg[1][3] ), .C(N_399), .Y(N_54));
    SLE \xhdl1.GEN_BITS[2].APB_32.edge_pos[2]  (.D(N_105), .CLK(
        FCCC_0_GL1), .EN(N_64), .ALn(MSS_RESET_N_F2M_c), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\edge_pos[2] ));
    CFG3 #( .INIT(8'h20) )  
        \xhdl1.GEN_BITS[24].APB_32.edge_both_RNO[24]  (.A(
        \CONFIG_reg[24][3] ), .B(CoreAPB3_0_APBmslave2_PWDATA[24]), .C(
        \edge_pos[24] ), .Y(N_100_i_0));
    SLE \xhdl1.GEN_BITS[1].APB_32.edge_both[1]  (.D(N_95), .CLK(
        FCCC_0_GL1), .EN(N_82), .ALn(MSS_RESET_N_F2M_c), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\edge_both[1] ));
    SLE \xhdl1.GEN_BITS[4].REG_GEN.CONFIG_reg[4][1]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[1]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[4]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[4][1] ));
    CFG4 #( .INIT(16'hAC0F) )  
        \xhdl1.GEN_BITS[26].REG_GEN.CONFIG_reg[26]_RNI0IFS1[0]  (.A(
        \CONFIG_reg[10][0] ), .B(\CONFIG_reg[26][0] ), .C(
        \CONFIG_reg_o_2_10_1_1[0] ), .D(CoreAPB3_0_APBmslave2_PADDR[5])
        , .Y(N_4731));
    SLE \xhdl1.GEN_BITS[17].REG_GEN.CONFIG_reg[17][3]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[3]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[17]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[17][3] ));
    SLE \xhdl1.GEN_BITS[30].APB_32.edge_both[30]  (.D(
        \edge_neg_429[30] ), .CLK(FCCC_0_GL1), .EN(
        edge_neg_2_sqmuxa_6_i_1), .ALn(MSS_RESET_N_F2M_c), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\edge_pos[30] ));
    SLE \xhdl1.GEN_BITS[3].APB_32.INTR_reg[3]  (.D(\INTR_reg_48[3] ), 
        .CLK(FCCC_0_GL1), .EN(VCC_net_1), .ALn(MSS_RESET_N_F2M_c), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\INTR_reg[3] ));
    CFG4 #( .INIT(16'h2000) )  GPOUT_reg_0_sqmuxa_0_a4_0_a2 (.A(
        CoreAPB3_0_APBmslave5_PSELx), .B(N_245), .C(wen_0), .D(N_610), 
        .Y(GPOUT_reg_0_sqmuxa));
    CFG3 #( .INIT(8'h20) )  
        \xhdl1.GEN_BITS[20].APB_32.edge_both_RNO[20]  (.A(
        \CONFIG_reg[20][3] ), .B(CoreAPB3_0_APBmslave2_PWDATA[20]), .C(
        \edge_neg[20] ), .Y(\edge_neg_289[20] ));
    CFG2 #( .INIT(4'h6) )  edge_both_2_sqmuxa_14_i_x2 (.A(\gpin2[1] ), 
        .B(gpin3_1), .Y(N_142_i));
    CFG4 #( .INIT(16'h0F35) )  
        \xhdl1.GEN_BITS[21].REG_GEN.CONFIG_reg[21]_RNIE8H61[6]  (.A(
        \CONFIG_reg[5][6] ), .B(\CONFIG_reg[21][6] ), .C(
        CoreAPB3_0_APBmslave2_PADDR[6]), .D(
        CoreAPB3_0_APBmslave2_PADDR[5]), .Y(\CONFIG_reg_o_2_21_1_1[6] )
        );
    SLE \xhdl1.GEN_BITS[6].REG_GEN.CONFIG_reg[6][4]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[4]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[6]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[6][4] ));
    SLE \xhdl1.GEN_BITS[3].REG_GEN.CONFIG_reg[3][6]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[6]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[3]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[3][6] ));
    CFG4 #( .INIT(16'hAC0F) )  
        \xhdl1.GEN_BITS[11].REG_GEN.CONFIG_reg[11]_RNIOTD72[4]  (.A(
        \CONFIG_reg[11][4] ), .B(\CONFIG_reg[27][4] ), .C(
        \CONFIG_reg_o_2_25_1_1[4] ), .D(CoreAPB3_0_APBmslave2_PADDR[5])
        , .Y(N_4855));
    SLE \xhdl1.GEN_BITS[4].gpin2[4]  (.D(\gpin1[4] ), .CLK(FCCC_0_GL1), 
        .EN(VCC_net_1), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(\gpin2[4] ));
    SLE \xhdl1.GEN_BITS[11].REG_GEN.CONFIG_reg[11][0]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[0]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[11]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[11][0] ));
    CFG4 #( .INIT(16'h0A33) )  
        \xhdl1.GEN_BITS[22].APB_32.INTR_reg_295_0[22]  (.A(INTR_reg_22)
        , .B(\INTR_reg_295_0_o2_1[22] ), .C(
        CoreAPB3_0_APBmslave2_PWDATA[22]), .D(edge_N_5_mux), .Y(
        \INTR_reg_295[22] ));
    CFG4 #( .INIT(16'hF2F3) )  
        \xhdl1.GEN_BITS[26].APB_32.INTR_reg_347_0_o2_1_0[26]  (.A(
        \CONFIG_reg[26][6] ), .B(\edge_pos[26] ), .C(
        \INTR_reg_347_0_o2_0[26] ), .D(\CONFIG_reg[26][5] ), .Y(
        \INTR_reg_347_0_o2_1[26] ));
    CFG4 #( .INIT(16'h0F35) )  
        \xhdl1.GEN_BITS[22].REG_GEN.CONFIG_reg[22]_RNIG3391[5]  (.A(
        \CONFIG_reg[6][5] ), .B(\CONFIG_reg[22][5] ), .C(
        CoreAPB3_0_APBmslave2_PADDR[6]), .D(
        CoreAPB3_0_APBmslave2_PADDR[5]), .Y(\CONFIG_reg_o_2_13_1_1[5] )
        );
    CFG4 #( .INIT(16'hAC0F) )  
        \xhdl1.GEN_BITS[24].REG_GEN.CONFIG_reg[24]_RNII4R22[4]  (.A(
        \CONFIG_reg[8][4] ), .B(\CONFIG_reg[24][4] ), .C(
        \CONFIG_reg_o_2_3_1[4] ), .D(CoreAPB3_0_APBmslave2_PADDR[5]), 
        .Y(N_4679));
    SLE \xhdl1.GEN_BITS[23].REG_GEN.CONFIG_reg[23][3]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[3]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[23]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[23][3] ));
    SLE \xhdl1.GEN_BITS[7].REG_GEN.CONFIG_reg[7][1]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[1]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[7]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[7][1] ));
    SLE \xhdl1.GEN_BITS[24].REG_GEN.CONFIG_reg[24][7]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[7]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[24]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[24][7] ));
    SLE \xhdl1.GEN_BITS[6].gpin1[6]  (.D(GPIO_IN_c[6]), .CLK(
        FCCC_0_GL1), .EN(VCC_net_1), .ALn(MSS_RESET_N_F2M_c), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\gpin1[6] ));
    SLE \xhdl1.GEN_BITS[24].REG_GEN.CONFIG_reg[24][5]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[5]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[24]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[24][5] ));
    CFG4 #( .INIT(16'hAA08) )  
        \xhdl1.GEN_BITS[5].APB_32.edge_pos_79_iv_i_0[5]  (.A(
        \CONFIG_reg[5][3] ), .B(\edge_pos[5] ), .C(
        CoreAPB3_0_APBmslave2_PWDATA[5]), .D(N_406), .Y(N_101));
    SLE \xhdl1.GEN_BITS[16].REG_GEN.CONFIG_reg[16][2]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[2]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[16]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[16][2] ));
    SLE \xhdl1.GEN_BITS[21].APB_32.INTR_reg[21]  (.D(
        \INTR_reg_282[21] ), .CLK(FCCC_0_GL1), .EN(VCC_net_1), .ALn(
        MSS_RESET_N_F2M_c), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(INTR_reg_21));
    SLE \xhdl1.GEN_BITS[27].REG_GEN.CONFIG_reg[27][3]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[3]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[27]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[27][3] ));
    CFG2 #( .INIT(4'hB) )  edge_both_2_sqmuxa_8_i (.A(edge_N_5_mux), 
        .B(\CONFIG_reg[20][3] ), .Y(N_196));
    SLE \xhdl1.GEN_BITS[27].REG_GEN.CONFIG_reg[27][5]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[5]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[27]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[27][5] ));
    CFG4 #( .INIT(16'hF2F3) )  
        \xhdl1.GEN_BITS[17].APB_32.INTR_reg_230_0_o2_1_0[17]  (.A(
        \CONFIG_reg[17][6] ), .B(\edge_neg[17] ), .C(
        \INTR_reg_230_0_o2_0[17] ), .D(\CONFIG_reg[17][5] ), .Y(
        \INTR_reg_230_0_o2_1[17] ));
    CFG4 #( .INIT(16'h0F35) )  
        \xhdl1.GEN_BITS[17].REG_GEN.CONFIG_reg[17]_RNI4TVJ1[0]  (.A(
        \CONFIG_reg[1][0] ), .B(\CONFIG_reg[17][0] ), .C(
        CoreAPB3_0_APBmslave2_PADDR[6]), .D(
        CoreAPB3_0_APBmslave2_PADDR[5]), .Y(\CONFIG_reg_o_2_18_1[0] ));
    SLE \xhdl1.GEN_BITS[13].REG_GEN.CONFIG_reg[13][0]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[0]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[13]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[13][0] ));
    CFG4 #( .INIT(16'hAC0F) )  
        \xhdl1.GEN_BITS[11].REG_GEN.CONFIG_reg[11]_RNI4AE72[7]  (.A(
        \CONFIG_reg[11][7] ), .B(\CONFIG_reg[27][7] ), .C(
        \CONFIG_reg_o_2_25_1_1[7] ), .D(CoreAPB3_0_APBmslave2_PADDR[5])
        , .Y(N_4858));
    CFG4 #( .INIT(16'h0A33) )  
        \xhdl1.GEN_BITS[30].APB_32.INTR_reg_399_0[30]  (.A(INTR_reg_30)
        , .B(\INTR_reg_399_0_o2_1[30] ), .C(
        CoreAPB3_0_APBmslave2_PWDATA[30]), .D(edge_N_5_mux), .Y(
        \INTR_reg_399[30] ));
    SLE \xhdl1.GEN_BITS[9].REG_GEN.CONFIG_reg[9][0]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[0]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[9]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[9][0] ));
    SLE \xhdl1.GEN_BITS[26].APB_32.edge_both[26]  (.D(N_106_i_0), .CLK(
        FCCC_0_GL1), .EN(N_159), .ALn(MSS_RESET_N_F2M_c), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\edge_pos[26] ));
    CFG2 #( .INIT(4'h8) )  
        \xhdl1.GEN_BITS[0].REG_GEN.CONFIG_reg[0]2_0_a4_0_a2  (.A(N_678)
        , .B(N_606), .Y(\CONFIG_reg[0]2 ));
    CFG2 #( .INIT(4'h2) )  edge_pos_2_sqmuxa_5_i_a2 (.A(\gpin2[1] ), 
        .B(gpin3_1), .Y(N_400));
    SLE \xhdl1.GEN_BITS[6].REG_GEN.CONFIG_reg[6][6]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[6]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[6]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[6][6] ));
    SLE \xhdl1.GEN_BITS[26].REG_GEN.CONFIG_reg[26][7]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[7]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[26]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[26][7] ));
    CFG4 #( .INIT(16'hAC0F) )  
        \xhdl1.GEN_BITS[14].REG_GEN.CONFIG_reg[14]_RNIG8Q82[5]  (.A(
        \CONFIG_reg[14][5] ), .B(\CONFIG_reg[30][5] ), .C(
        \CONFIG_reg_o_2_13_1_1[5] ), .D(CoreAPB3_0_APBmslave2_PADDR[5])
        , .Y(N_4760));
    CFG4 #( .INIT(16'hF2F3) )  
        \xhdl1.GEN_BITS[9].APB_32.INTR_reg_126_0_o2_1_0[9]  (.A(
        \CONFIG_reg[9][6] ), .B(\edge_neg[9] ), .C(
        \INTR_reg_126_0_o2_0[9] ), .D(\CONFIG_reg[9][5] ), .Y(
        \INTR_reg_126_0_o2_1[9] ));
    SLE \xhdl1.GEN_BITS[8].REG_GEN.CONFIG_reg[8][0]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[0]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[8]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[8][0] ));
    CFG4 #( .INIT(16'h0800) )  
        \xhdl1.GEN_BITS[4].REG_GEN.CONFIG_reg[4]2_0_a4_0_a2_0_RNIBB9M2  
        (.A(N_603), .B(r_m1_e_1_0), .C(N_245), .D(
        CoreAPB3_0_APBmslave5_PSELx), .Y(
        \CONFIG_reg[4]2_0_a4_0_a2_0_RNIBB9M2 ));
    SLE \xhdl1.GEN_BITS[1].gpin2[1]  (.D(\gpin1[1] ), .CLK(FCCC_0_GL1), 
        .EN(VCC_net_1), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(\gpin2[1] ));
    SLE \xhdl1.GEN_BITS[11].REG_GEN.CONFIG_reg[11][7]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[7]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[11]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[11][7] ));
    SLE \xhdl1.GEN_BITS[15].REG_GEN.CONFIG_reg[15][3]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[3]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[15]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[15][3] ));
    SLE \xhdl1.GEN_BITS[3].gpin2[3]  (.D(\gpin1[3] ), .CLK(FCCC_0_GL1), 
        .EN(VCC_net_1), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(\gpin2[3] ));
    CFG4 #( .INIT(16'hAC0F) )  
        \xhdl1.GEN_BITS[15].REG_GEN.CONFIG_reg[15]_RNIS7O32[6]  (.A(
        \CONFIG_reg[15][6] ), .B(\CONFIG_reg[31][6] ), .C(
        \CONFIG_reg_o_2_28_1_1[6] ), .D(CoreAPB3_0_APBmslave2_PADDR[5])
        , .Y(N_4881));
    SLE \xhdl1.GEN_BITS[31].REG_GEN.CONFIG_reg[31][6]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[6]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[31]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[31][6] ));
    SLE \xhdl1.GEN_BITS[25].REG_GEN.CONFIG_reg[25][0]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[0]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[25]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[25][0] ));
    SLE \xhdl1.GEN_BITS[21].REG_GEN.CONFIG_reg[21][1]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[1]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[21]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[21][1] ));
    CFG4 #( .INIT(16'h0F35) )  
        \xhdl1.GEN_BITS[22].REG_GEN.CONFIG_reg[22]_RNI8R291[1]  (.A(
        \CONFIG_reg[6]_1 ), .B(\CONFIG_reg[22][1] ), .C(
        CoreAPB3_0_APBmslave2_PADDR[6]), .D(
        CoreAPB3_0_APBmslave2_PADDR[5]), .Y(\CONFIG_reg_o_2_13_1_1[1] )
        );
    SLE \xhdl1.GEN_BITS[28].APB_32.edge_both[28]  (.D(N_87_i_0), .CLK(
        FCCC_0_GL1), .EN(N_163), .ALn(MSS_RESET_N_F2M_c), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\edge_pos[28] ));
    SLE \xhdl1.GEN_BITS[23].APB_32.GPOUT_reg[23]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[23]), .CLK(FCCC_0_GL1), .EN(
        GPOUT_reg_0_sqmuxa), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        GPOUT_reg_23));
    SLE \xhdl1.GEN_BITS[0].gpin1[0]  (.D(GPIO_IN_c[0]), .CLK(
        FCCC_0_GL1), .EN(VCC_net_1), .ALn(MSS_RESET_N_F2M_c), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\gpin1[0] ));
    CFG4 #( .INIT(16'hAC0F) )  
        \xhdl1.GEN_BITS[11].REG_GEN.CONFIG_reg[11]_RNIGLD72[2]  (.A(
        \CONFIG_reg[11][2] ), .B(\CONFIG_reg[27][2] ), .C(
        \CONFIG_reg_o_2_25_1_1[2] ), .D(CoreAPB3_0_APBmslave2_PADDR[5])
        , .Y(N_4853));
    CFG3 #( .INIT(8'h20) )  
        \xhdl1.GEN_BITS[19].APB_32.edge_both_RNO[19]  (.A(
        \CONFIG_reg[19][3] ), .B(CoreAPB3_0_APBmslave2_PWDATA[19]), .C(
        \edge_neg[19] ), .Y(\edge_neg_275[19] ));
    CFG4 #( .INIT(16'hAC0F) )  
        \xhdl1.GEN_BITS[28].REG_GEN.CONFIG_reg[28]_RNI2NKA2[1]  (.A(
        \CONFIG_reg[12][1] ), .B(\CONFIG_reg[28][1] ), .C(
        \CONFIG_reg_o_2_6_1_1[1] ), .D(CoreAPB3_0_APBmslave2_PADDR[5]), 
        .Y(N_4700));
    CFG4 #( .INIT(16'hAC0F) )  
        \xhdl1.GEN_BITS[11].REG_GEN.CONFIG_reg[11]_RNICHD72[1]  (.A(
        \CONFIG_reg[11][1] ), .B(\CONFIG_reg[27][1] ), .C(
        \CONFIG_reg_o_2_25_1_1[1] ), .D(CoreAPB3_0_APBmslave2_PADDR[5])
        , .Y(N_4852));
    SLE \xhdl1.GEN_BITS[3].REG_GEN.CONFIG_reg[3][0]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[0]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[3]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[3][0] ));
    CFG2 #( .INIT(4'hB) )  edge_both_2_sqmuxa_18_i (.A(edge_N_5_mux), 
        .B(\CONFIG_reg[10][3] ), .Y(N_184));
    SLE \xhdl1.GEN_BITS[5].gpin3[5]  (.D(\gpin2[5] ), .CLK(FCCC_0_GL1), 
        .EN(VCC_net_1), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(gpin3_5));
    SLE \xhdl1.GEN_BITS[18].APB_32.edge_both[18]  (.D(
        \edge_neg_261[18] ), .CLK(FCCC_0_GL1), .EN(N_192), .ALn(
        MSS_RESET_N_F2M_c), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\edge_neg[18] ));
    CFG4 #( .INIT(16'h0F35) )  
        \xhdl1.GEN_BITS[21].REG_GEN.CONFIG_reg[21]_RNI82H61[3]  (.A(
        \CONFIG_reg[5][3] ), .B(\CONFIG_reg[21][3] ), .C(
        CoreAPB3_0_APBmslave2_PADDR[6]), .D(
        CoreAPB3_0_APBmslave2_PADDR[5]), .Y(\CONFIG_reg_o_2_21_1[3] ));
    CFG4 #( .INIT(16'hF2F3) )  
        \xhdl1.GEN_BITS[8].APB_32.INTR_reg_113_0_o2_1_0[8]  (.A(
        \CONFIG_reg[8][6] ), .B(\edge_pos[8] ), .C(
        \INTR_reg_113_0_o2_0[8] ), .D(\CONFIG_reg[8][5] ), .Y(
        \INTR_reg_113_0_o2_1[8] ));
    SLE \xhdl1.GEN_BITS[0].APB_32.GPOUT_reg[0]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[0]), .CLK(FCCC_0_GL1), .EN(
        GPOUT_reg_0_sqmuxa), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        GPOUT_reg_0));
    CFG2 #( .INIT(4'hB) )  edge_both_2_sqmuxa_29_i (.A(edge_N_5_mux), 
        .B(\CONFIG_reg[26][3] ), .Y(N_159));
    SLE \xhdl1.GEN_BITS[31].REG_GEN.CONFIG_reg[31][7]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[7]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[31]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[31][7] ));
    SLE \xhdl1.GEN_BITS[19].REG_GEN.CONFIG_reg[19][6]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[6]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[19]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[19][6] ));
    CFG4 #( .INIT(16'h0F35) )  
        \xhdl1.GEN_BITS[4].REG_GEN.CONFIG_reg[4]_RNIABV31[6]  (.A(
        \CONFIG_reg[4][6] ), .B(\CONFIG_reg[20][6] ), .C(
        CoreAPB3_0_APBmslave2_PADDR[6]), .D(
        CoreAPB3_0_APBmslave2_PADDR[5]), .Y(\CONFIG_reg_o_2_6_1_1[6] ));
    CFG4 #( .INIT(16'hC5CA) )  
        \xhdl1.GEN_BITS[1].APB_32.INTR_reg_22_0_m2[1]  (.A(gpin3_1), 
        .B(N_174), .C(\CONFIG_reg[1][6] ), .D(\CONFIG_reg[1][5] ), .Y(
        N_177));
    CFG4 #( .INIT(16'hF2F3) )  
        \xhdl1.GEN_BITS[14].APB_32.INTR_reg_191_0_o2_1_0[14]  (.A(
        \CONFIG_reg[14][6] ), .B(\edge_neg[14] ), .C(
        \INTR_reg_191_0_o2_0[14] ), .D(\CONFIG_reg[14][5] ), .Y(
        \INTR_reg_191_0_o2_1[14] ));
    CFG3 #( .INIT(8'h20) )  
        \xhdl1.GEN_BITS[22].APB_32.edge_both_RNO[22]  (.A(
        \CONFIG_reg[22][3] ), .B(CoreAPB3_0_APBmslave2_PWDATA[22]), .C(
        \edge_neg[22] ), .Y(\edge_neg_317[22] ));
    CFG2 #( .INIT(4'h2) )  
        \xhdl1.GEN_BITS[0].APB_32.GPOUT_reg9_0_a2_2_a2_0  (.A(
        CoreAPB3_0_APBmslave2_PADDR[5]), .B(
        CoreAPB3_0_APBmslave2_PADDR[4]), .Y(N_610));
    SLE \xhdl1.GEN_BITS[12].REG_GEN.CONFIG_reg[12][5]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[5]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[12]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[12][5] ));
    SLE \xhdl1.GEN_BITS[19].APB_32.GPOUT_reg[19]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[19]), .CLK(FCCC_0_GL1), .EN(
        GPOUT_reg_0_sqmuxa), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        GPOUT_reg_19));
    SLE \xhdl1.GEN_BITS[18].REG_GEN.CONFIG_reg[18][4]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[4]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[18]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[18][4] ));
    CFG3 #( .INIT(8'h20) )  
        \xhdl1.GEN_BITS[11].APB_32.edge_both_RNO[11]  (.A(
        \CONFIG_reg[11][3] ), .B(CoreAPB3_0_APBmslave2_PWDATA[11]), .C(
        \edge_neg[11] ), .Y(\edge_neg_163[11] ));
    SLE \xhdl1.GEN_BITS[6].APB_32.INTR_reg[6]  (.D(\INTR_reg_87[6] ), 
        .CLK(FCCC_0_GL1), .EN(VCC_net_1), .ALn(MSS_RESET_N_F2M_c), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(INTR_reg_6));
    SLE \xhdl1.GEN_BITS[0].REG_GEN.CONFIG_reg[0][5]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[5]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[0]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[0][5] ));
    SLE \xhdl1.GEN_BITS[3].APB_32.edge_pos[3]  (.D(N_73), .CLK(
        FCCC_0_GL1), .EN(N_79), .ALn(MSS_RESET_N_F2M_c), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\edge_pos[3] ));
    SLE \xhdl1.GEN_BITS[9].APB_32.edge_both[9]  (.D(\edge_neg_135[9] ), 
        .CLK(FCCC_0_GL1), .EN(N_182), .ALn(MSS_RESET_N_F2M_c), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\edge_neg[9] ));
    SLE \xhdl1.GEN_BITS[6].REG_GEN.CONFIG_reg[6][0]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[0]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[6]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[6][0] ));
    CFG4 #( .INIT(16'hA9FF) )  
        \xhdl1.GEN_BITS[22].APB_32.INTR_reg_295_0_o2_0_0[22]  (.A(
        \CONFIG_reg[22][7] ), .B(\CONFIG_reg[22][6] ), .C(
        \CONFIG_reg[22][5] ), .D(\CONFIG_reg[22][3] ), .Y(
        \INTR_reg_295_0_o2_0[22] ));
    CFG2 #( .INIT(4'h6) )  
        \xhdl1.GEN_BITS[3].APB_32.edge_both_51_iv_0_x2[3]  (.A(
        \gpin2[3] ), .B(gpin3_3), .Y(N_253_i));
    SLE \xhdl1.GEN_BITS[15].REG_GEN.CONFIG_reg[15][6]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[6]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[15]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[15][6] ));
    SLE \xhdl1.GEN_BITS[5].REG_GEN.CONFIG_reg[5][2]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[2]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[5]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[5][2] ));
    SLE \xhdl1.GEN_BITS[27].APB_32.INTR_reg[27]  (.D(
        \INTR_reg_360[27] ), .CLK(FCCC_0_GL1), .EN(VCC_net_1), .ALn(
        MSS_RESET_N_F2M_c), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(INTR_reg_27));
    CFG4 #( .INIT(16'hAC0F) )  
        \xhdl1.GEN_BITS[24].REG_GEN.CONFIG_reg[24]_RNIE0R22[3]  (.A(
        \CONFIG_reg[8][3] ), .B(\CONFIG_reg[24][3] ), .C(
        \CONFIG_reg_o_2_3_1[3] ), .D(CoreAPB3_0_APBmslave2_PADDR[5]), 
        .Y(N_4678));
    CFG4 #( .INIT(16'hAC0F) )  
        \xhdl1.GEN_BITS[26].REG_GEN.CONFIG_reg[26]_RNIOAGS1[6]  (.A(
        \CONFIG_reg[10][6] ), .B(\CONFIG_reg[26][6] ), .C(
        \CONFIG_reg_o_2_10_1_1[6] ), .D(CoreAPB3_0_APBmslave2_PADDR[5])
        , .Y(N_4737));
    CFG3 #( .INIT(8'h20) )  
        \xhdl1.GEN_BITS[13].APB_32.edge_both_RNO[13]  (.A(
        \CONFIG_reg[13][3] ), .B(CoreAPB3_0_APBmslave2_PWDATA[13]), .C(
        \edge_neg[13] ), .Y(\edge_neg_191[13] ));
    CFG3 #( .INIT(8'hFB) )  edge_neg_2_sqmuxa_i_0_0 (.A(edge_N_5_mux), 
        .B(\CONFIG_reg[6][3] ), .C(N_688), .Y(N_62));
    CFG3 #( .INIT(8'h04) )  
        \xhdl1.GEN_BITS[6].APB_32.INTR_reg_87_0_0_0_tz_1[6]  (.A(
        \CONFIG_reg[6][5] ), .B(\edge_both[6] ), .C(\CONFIG_reg[6][6] )
        , .Y(\INTR_reg_87_0_0_0_tz_1[6] ));
    SLE \xhdl1.GEN_BITS[19].APB_32.edge_both[19]  (.D(
        \edge_neg_275[19] ), .CLK(FCCC_0_GL1), .EN(N_194), .ALn(
        MSS_RESET_N_F2M_c), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\edge_neg[19] ));
    CFG4 #( .INIT(16'hF2F3) )  
        \xhdl1.GEN_BITS[15].APB_32.INTR_reg_204_0_o2_1_0[15]  (.A(
        \CONFIG_reg[15][6] ), .B(\edge_neg[15] ), .C(
        \INTR_reg_204_0_o2_0[15] ), .D(\CONFIG_reg[15][5] ), .Y(
        \INTR_reg_204_0_o2_1[15] ));
    CFG4 #( .INIT(16'h0F35) )  
        \xhdl1.GEN_BITS[16].REG_GEN.CONFIG_reg[16]_RNIAAE11[5]  (.A(
        \CONFIG_reg[0][5] ), .B(\CONFIG_reg[16][5] ), .C(
        CoreAPB3_0_APBmslave2_PADDR[6]), .D(
        CoreAPB3_0_APBmslave2_PADDR[5]), .Y(\CONFIG_reg_o_2_3_1_1[5] ));
    SLE \xhdl1.GEN_BITS[4].REG_GEN.CONFIG_reg[4][2]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[2]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[4]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[4][2] ));
    CFG2 #( .INIT(4'hB) )  edge_both_2_sqmuxa_24_i (.A(edge_N_5_mux), 
        .B(\CONFIG_reg[31][3] ), .Y(edge_pos_2_sqmuxa_19_i_1));
    CFG4 #( .INIT(16'h0A33) )  
        \xhdl1.GEN_BITS[15].APB_32.INTR_reg_204_0[15]  (.A(INTR_reg_15)
        , .B(\INTR_reg_204_0_o2_1[15] ), .C(
        CoreAPB3_0_APBmslave2_PWDATA[15]), .D(edge_N_5_mux), .Y(
        \INTR_reg_204[15] ));
    SLE \xhdl1.GEN_BITS[28].REG_GEN.CONFIG_reg[28][6]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[6]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[28]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[28][6] ));
    SLE \xhdl1.GEN_BITS[11].REG_GEN.CONFIG_reg[11][4]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[4]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[11]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[11][4] ));
    SLE \xhdl1.GEN_BITS[28].REG_GEN.CONFIG_reg[28][3]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[3]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[28]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[28][3] ));
    SLE \xhdl1.GEN_BITS[23].REG_GEN.CONFIG_reg[23][5]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[5]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[23]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[23][5] ));
    SLE \xhdl1.GEN_BITS[4].gpin1[4]  (.D(GPIO_IN_c[4]), .CLK(
        FCCC_0_GL1), .EN(VCC_net_1), .ALn(MSS_RESET_N_F2M_c), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\gpin1[4] ));
    CFG4 #( .INIT(16'hAA08) )  
        \xhdl1.GEN_BITS[5].APB_32.edge_neg_79_iv_i_0[5]  (.A(
        \CONFIG_reg[5][3] ), .B(\edge_neg[5] ), .C(
        CoreAPB3_0_APBmslave2_PWDATA[5]), .D(N_405), .Y(N_115));
    CFG4 #( .INIT(16'h0F35) )  
        \xhdl1.GEN_BITS[22].REG_GEN.CONFIG_reg[22]_RNICV291[3]  (.A(
        \CONFIG_reg[6][3] ), .B(\CONFIG_reg[22][3] ), .C(
        CoreAPB3_0_APBmslave2_PADDR[6]), .D(
        CoreAPB3_0_APBmslave2_PADDR[5]), .Y(\CONFIG_reg_o_2_13_1_1[3] )
        );
    SLE \xhdl1.GEN_BITS[9].REG_GEN.CONFIG_reg[9][1]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[1]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[9]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[9][1] ));
    CFG4 #( .INIT(16'hAC0F) )  
        \xhdl1.GEN_BITS[29].REG_GEN.CONFIG_reg[29]_RNI6EI52[0]  (.A(
        \CONFIG_reg[13][0] ), .B(\CONFIG_reg[29][0] ), .C(
        \CONFIG_reg_o_2_21_1[0] ), .D(CoreAPB3_0_APBmslave2_PADDR[5]), 
        .Y(N_4819));
    SLE \xhdl1.GEN_BITS[18].REG_GEN.CONFIG_reg[18][1]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[1]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[18]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[18][1] ));
    SLE \xhdl1.GEN_BITS[10].APB_32.INTR_reg[10]  (.D(
        \INTR_reg_139[10] ), .CLK(FCCC_0_GL1), .EN(VCC_net_1), .ALn(
        MSS_RESET_N_F2M_c), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(INTR_reg_10));
    SLE \xhdl1.GEN_BITS[12].REG_GEN.CONFIG_reg[12][3]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[3]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[12]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[12][3] ));
    SLE \xhdl1.GEN_BITS[18].REG_GEN.CONFIG_reg[18][5]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[5]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[18]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[18][5] ));
    SLE \xhdl1.GEN_BITS[4].APB_32.edge_neg[4]  (.D(N_117), .CLK(
        FCCC_0_GL1), .EN(N_58), .ALn(MSS_RESET_N_F2M_c), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\edge_neg[4] ));
    SLE \xhdl1.GEN_BITS[20].APB_32.edge_both[20]  (.D(
        \edge_neg_289[20] ), .CLK(FCCC_0_GL1), .EN(N_196), .ALn(
        MSS_RESET_N_F2M_c), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\edge_neg[20] ));
    SLE \xhdl1.GEN_BITS[17].APB_32.GPOUT_reg[17]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[17]), .CLK(FCCC_0_GL1), .EN(
        GPOUT_reg_0_sqmuxa), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        GPOUT_reg_17));
    SLE \xhdl1.GEN_BITS[8].REG_GEN.CONFIG_reg[8][1]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[1]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[8]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[8][1] ));
    SLE \xhdl1.GEN_BITS[7].REG_GEN.CONFIG_reg[7][2]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[2]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[7]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[7][2] ));
    CFG3 #( .INIT(8'h20) )  
        \xhdl1.GEN_BITS[27].APB_32.edge_both_RNO[27]  (.A(
        \CONFIG_reg[27][3] ), .B(CoreAPB3_0_APBmslave2_PWDATA[27]), .C(
        \edge_neg[27] ), .Y(N_5912_i_0));
    CFG4 #( .INIT(16'hAC0F) )  
        \xhdl1.GEN_BITS[29].REG_GEN.CONFIG_reg[29]_RNIQ2J52[5]  (.A(
        \CONFIG_reg[13][5] ), .B(\CONFIG_reg[29][5] ), .C(
        \CONFIG_reg_o_2_21_1_1[5] ), .D(CoreAPB3_0_APBmslave2_PADDR[5])
        , .Y(N_4824));
    CFG4 #( .INIT(16'h0F35) )  
        \xhdl1.GEN_BITS[21].REG_GEN.CONFIG_reg[21]_RNI60H61[2]  (.A(
        \CONFIG_reg[5][2] ), .B(\CONFIG_reg[21][2] ), .C(
        CoreAPB3_0_APBmslave2_PADDR[6]), .D(
        CoreAPB3_0_APBmslave2_PADDR[5]), .Y(\CONFIG_reg_o_2_21_1_1[2] )
        );
    SLE \xhdl1.GEN_BITS[21].REG_GEN.CONFIG_reg[21][5]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[5]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[21]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[21][5] ));
    CFG4 #( .INIT(16'h0F35) )  
        \xhdl1.GEN_BITS[18].REG_GEN.CONFIG_reg[18]_RNIASH61[1]  (.A(
        \CONFIG_reg[2]_1 ), .B(\CONFIG_reg[18][1] ), .C(
        CoreAPB3_0_APBmslave2_PADDR[6]), .D(
        CoreAPB3_0_APBmslave2_PADDR[5]), .Y(\CONFIG_reg_o_2_10_1_1[1] )
        );
    CFG4 #( .INIT(16'h1000) )  
        \xhdl1.GEN_BITS[16].REG_GEN.CONFIG_reg[16]2_0_a4_0_a2  (.A(
        CoreAPB3_0_APBmslave2_PADDR[3]), .B(
        CoreAPB3_0_APBmslave2_PADDR[2]), .C(N_598), .D(N_606), .Y(
        \CONFIG_reg[16]2 ));
    SLE \xhdl1.GEN_BITS[14].REG_GEN.CONFIG_reg[14][2]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[2]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[14]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[14][2] ));
    SLE \xhdl1.GEN_BITS[24].APB_32.INTR_reg[24]  (.D(
        \INTR_reg_321[24] ), .CLK(FCCC_0_GL1), .EN(VCC_net_1), .ALn(
        MSS_RESET_N_F2M_c), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(INTR_reg_24));
    CFG4 #( .INIT(16'hAC0F) )  
        \xhdl1.GEN_BITS[28].REG_GEN.CONFIG_reg[28]_RNIE3LA2[4]  (.A(
        \CONFIG_reg[12][4] ), .B(\CONFIG_reg[28][4] ), .C(
        \CONFIG_reg_o_2_6_1[4] ), .D(CoreAPB3_0_APBmslave2_PADDR[5]), 
        .Y(N_4703));
    CFG4 #( .INIT(16'h0A33) )  
        \xhdl1.GEN_BITS[25].APB_32.INTR_reg_334_0[25]  (.A(INTR_reg_25)
        , .B(\INTR_reg_334_0_o2_1[25] ), .C(
        CoreAPB3_0_APBmslave2_PWDATA[25]), .D(edge_N_5_mux), .Y(
        \INTR_reg_334[25] ));
    CFG2 #( .INIT(4'hB) )  edge_both_2_sqmuxa_26_i (.A(edge_N_5_mux), 
        .B(\CONFIG_reg[23][3] ), .Y(edge_pos_2_sqmuxa_26_i_1));
    SLE \xhdl1.GEN_BITS[0].APB_32.edge_both[0]  (.D(N_97), .CLK(
        FCCC_0_GL1), .EN(N_80), .ALn(MSS_RESET_N_F2M_c), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\edge_both[0] ));
    SLE \xhdl1.GEN_BITS[14].APB_32.edge_both[14]  (.D(
        \edge_neg_205[14] ), .CLK(FCCC_0_GL1), .EN(
        edge_pos_2_sqmuxa_8_i_1), .ALn(MSS_RESET_N_F2M_c), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\edge_neg[14] ));
    SLE \xhdl1.GEN_BITS[8].APB_32.INTR_reg[8]  (.D(\INTR_reg_113[8] ), 
        .CLK(FCCC_0_GL1), .EN(VCC_net_1), .ALn(MSS_RESET_N_F2M_c), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(INTR_reg_8));
    SLE \xhdl1.GEN_BITS[22].REG_GEN.CONFIG_reg[22][0]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[0]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[22]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[22][0] ));
    SLE \xhdl1.GEN_BITS[3].REG_GEN.CONFIG_reg[3][1]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[1]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[3]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[3]_1 ));
    CFG4 #( .INIT(16'h0F35) )  
        \xhdl1.GEN_BITS[7].REG_GEN.CONFIG_reg[7]_RNIAMKB1[0]  (.A(
        \CONFIG_reg[7][0] ), .B(\CONFIG_reg[23][0] ), .C(
        CoreAPB3_0_APBmslave2_PADDR[6]), .D(
        CoreAPB3_0_APBmslave2_PADDR[5]), .Y(\CONFIG_reg_o_2_28_1_1[0] )
        );
    SLE \xhdl1.GEN_BITS[13].APB_32.edge_both[13]  (.D(
        \edge_neg_191[13] ), .CLK(FCCC_0_GL1), .EN(
        edge_pos_2_sqmuxa_9_i_1), .ALn(MSS_RESET_N_F2M_c), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\edge_neg[13] ));
    CFG2 #( .INIT(4'hB) )  edge_both_2_sqmuxa_19_i (.A(edge_N_5_mux), 
        .B(\CONFIG_reg[9][3] ), .Y(N_182));
    SLE \xhdl1.GEN_BITS[11].REG_GEN.CONFIG_reg[11][2]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[2]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[11]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[11][2] ));
    CFG4 #( .INIT(16'hAA08) )  
        \xhdl1.GEN_BITS[0].APB_32.edge_neg_9_iv_i_0[0]  (.A(
        \CONFIG_reg[0][3] ), .B(\edge_neg[0] ), .C(
        CoreAPB3_0_APBmslave2_PWDATA[0]), .D(N_401), .Y(N_123));
    SLE \xhdl1.GEN_BITS[17].REG_GEN.CONFIG_reg[17][7]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[7]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[17]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[17][7] ));
    SLE \xhdl1.GEN_BITS[5].APB_32.edge_pos[5]  (.D(N_101), .CLK(
        FCCC_0_GL1), .EN(N_70), .ALn(MSS_RESET_N_F2M_c), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\edge_pos[5] ));
    SLE \xhdl1.GEN_BITS[29].REG_GEN.CONFIG_reg[29][4]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[4]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[29]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[29][4] ));
    CFG4 #( .INIT(16'hF2F3) )  
        \xhdl1.GEN_BITS[21].APB_32.INTR_reg_282_0_o2_1_0[21]  (.A(
        \CONFIG_reg[21][6] ), .B(\edge_neg[21] ), .C(
        \INTR_reg_282_0_o2_0[21] ), .D(\CONFIG_reg[21][5] ), .Y(
        \INTR_reg_282_0_o2_1[21] ));
    SLE \xhdl1.GEN_BITS[15].REG_GEN.CONFIG_reg[15][1]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[1]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[15]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[15][1] ));
    CFG4 #( .INIT(16'hAC0F) )  
        \xhdl1.GEN_BITS[28].REG_GEN.CONFIG_reg[28]_RNIMBLA2[6]  (.A(
        \CONFIG_reg[12][6] ), .B(\CONFIG_reg[28][6] ), .C(
        \CONFIG_reg_o_2_6_1_1[6] ), .D(CoreAPB3_0_APBmslave2_PADDR[5]), 
        .Y(N_4705));
    CFG4 #( .INIT(16'h4000) )  
        \xhdl1.GEN_BITS[25].REG_GEN.CONFIG_reg[25]2_0_a4_0_a2  (.A(
        CoreAPB3_0_APBmslave2_PADDR[3]), .B(
        CoreAPB3_0_APBmslave2_PADDR[2]), .C(N_598), .D(N_610), .Y(
        \CONFIG_reg[25]2 ));
    CFG3 #( .INIT(8'h20) )  
        \xhdl1.GEN_BITS[26].APB_32.edge_both_RNO[26]  (.A(
        \CONFIG_reg[26][3] ), .B(CoreAPB3_0_APBmslave2_PWDATA[26]), .C(
        \edge_pos[26] ), .Y(N_106_i_0));
    CFG4 #( .INIT(16'h8000) )  
        \xhdl1.GEN_BITS[31].REG_GEN.CONFIG_reg[31]2_0_a4_0_a2  (.A(
        CoreAPB3_0_APBmslave2_PADDR[3]), .B(
        CoreAPB3_0_APBmslave2_PADDR[2]), .C(N_598), .D(N_605), .Y(
        \CONFIG_reg[31]2 ));
    SLE \xhdl1.GEN_BITS[31].REG_GEN.CONFIG_reg[31][0]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[0]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[31]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[31][0] ));
    SLE \xhdl1.GEN_BITS[5].gpin1[5]  (.D(GPIO_IN_c[5]), .CLK(
        FCCC_0_GL1), .EN(VCC_net_1), .ALn(MSS_RESET_N_F2M_c), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\gpin1[5] ));
    SLE \xhdl1.GEN_BITS[11].REG_GEN.CONFIG_reg[11][5]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[5]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[11]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[11][5] ));
    SLE \xhdl1.GEN_BITS[6].REG_GEN.CONFIG_reg[6][1]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[1]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[6]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[6]_1 ));
    SLE \xhdl1.GEN_BITS[2].APB_32.INTR_reg[2]  (.D(\INTR_reg_35[2] ), 
        .CLK(FCCC_0_GL1), .EN(VCC_net_1), .ALn(MSS_RESET_N_F2M_c), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(INTR_reg_2));
    CFG4 #( .INIT(16'h0F35) )  
        \xhdl1.GEN_BITS[17].REG_GEN.CONFIG_reg[17]_RNI810K1[2]  (.A(
        \CONFIG_reg[1][2] ), .B(\CONFIG_reg[17][2] ), .C(
        CoreAPB3_0_APBmslave2_PADDR[6]), .D(
        CoreAPB3_0_APBmslave2_PADDR[5]), .Y(\CONFIG_reg_o_2_18_1_1[2] )
        );
    CFG3 #( .INIT(8'h20) )  
        \xhdl1.GEN_BITS[18].APB_32.edge_both_RNO[18]  (.A(
        \CONFIG_reg[18][3] ), .B(CoreAPB3_0_APBmslave2_PWDATA[18]), .C(
        \edge_neg[18] ), .Y(\edge_neg_261[18] ));
    CFG3 #( .INIT(8'h20) )  
        \xhdl1.GEN_BITS[29].APB_32.edge_both_RNO[29]  (.A(
        \CONFIG_reg[29][3] ), .B(CoreAPB3_0_APBmslave2_PWDATA[29]), .C(
        \edge_pos[29] ), .Y(\edge_neg_415[29] ));
    CFG4 #( .INIT(16'h0ACC) )  
        \xhdl1.GEN_BITS[1].APB_32.INTR_reg_22_0_0[1]  (.A(INTR_reg_1), 
        .B(\INTR_reg_22_0_0_0_tz[1] ), .C(
        CoreAPB3_0_APBmslave2_PWDATA[1]), .D(edge_N_5_mux), .Y(
        \INTR_reg_22[1] ));
    CFG4 #( .INIT(16'h0A33) )  
        \xhdl1.GEN_BITS[11].APB_32.INTR_reg_152_0[11]  (.A(INTR_reg_11)
        , .B(\INTR_reg_152_0_o2_1[11] ), .C(
        CoreAPB3_0_APBmslave2_PWDATA[11]), .D(edge_N_5_mux), .Y(
        \INTR_reg_152[11] ));
    SLE \xhdl1.GEN_BITS[28].APB_32.INTR_reg[28]  (.D(
        \INTR_reg_373[28] ), .CLK(FCCC_0_GL1), .EN(VCC_net_1), .ALn(
        MSS_RESET_N_F2M_c), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(INTR_reg_28));
    CFG4 #( .INIT(16'hAC0F) )  
        \xhdl1.GEN_BITS[14].REG_GEN.CONFIG_reg[14]_RNIOGQ82[7]  (.A(
        \CONFIG_reg[14][7] ), .B(\CONFIG_reg[30][7] ), .C(
        \CONFIG_reg_o_2_13_1_1[7] ), .D(CoreAPB3_0_APBmslave2_PADDR[5])
        , .Y(N_4762));
    CFG4 #( .INIT(16'h0200) )  
        \xhdl1.GEN_BITS[0].APB_32.un5_PRDATA_o_0_a2_0_o2_s_RNIBS2P2  (
        .A(CoreAPB3_0_APBmslave5_PSELx), .B(N_245), .C(
        un5_PRDATA_o_0_a2_0_o2_out), .D(wen_0), .Y(edge_N_5_mux));
    CFG4 #( .INIT(16'hA9FF) )  
        \xhdl1.GEN_BITS[25].APB_32.INTR_reg_334_0_o2_0_0[25]  (.A(
        \CONFIG_reg[25][7] ), .B(\CONFIG_reg[25][6] ), .C(
        \CONFIG_reg[25][5] ), .D(\CONFIG_reg[25][3] ), .Y(
        \INTR_reg_334_0_o2_0[25] ));
    CFG4 #( .INIT(16'h0F35) )  
        \xhdl1.GEN_BITS[16].REG_GEN.CONFIG_reg[16]_RNI22E11[1]  (.A(
        \CONFIG_reg[0]_1 ), .B(\CONFIG_reg[16][1] ), .C(
        CoreAPB3_0_APBmslave2_PADDR[6]), .D(
        CoreAPB3_0_APBmslave2_PADDR[5]), .Y(\CONFIG_reg_o_2_3_1_1[1] ));
    SLE \xhdl1.GEN_BITS[17].APB_32.edge_both[17]  (.D(
        \edge_neg_247[17] ), .CLK(FCCC_0_GL1), .EN(
        edge_pos_2_sqmuxa_30_i_1), .ALn(MSS_RESET_N_F2M_c), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\edge_neg[17] ));
    CFG3 #( .INIT(8'h04) )  
        \xhdl1.GEN_BITS[2].APB_32.INTR_reg_35_0_0_0_tz_1[2]  (.A(
        \CONFIG_reg[2][5] ), .B(\edge_both[2] ), .C(\CONFIG_reg[2][6] )
        , .Y(\INTR_reg_35_0_0_0_tz_1[2] ));
    SLE \xhdl1.GEN_BITS[5].gpin2[5]  (.D(\gpin1[5] ), .CLK(FCCC_0_GL1), 
        .EN(VCC_net_1), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(\gpin2[5] ));
    SLE \xhdl1.GEN_BITS[26].REG_GEN.CONFIG_reg[26][3]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[3]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[26]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[26][3] ));
    CFG2 #( .INIT(4'h2) )  edge_pos_2_sqmuxa_6_i_a2 (.A(\gpin2[2] ), 
        .B(gpin3_2), .Y(N_396));
    SLE \xhdl1.GEN_BITS[12].APB_32.edge_both[12]  (.D(
        \edge_neg_177[12] ), .CLK(FCCC_0_GL1), .EN(N_188), .ALn(
        MSS_RESET_N_F2M_c), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\edge_neg[12] ));
    SLE \xhdl1.GEN_BITS[27].REG_GEN.CONFIG_reg[27][1]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[1]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[27]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[27][1] ));
    CFG4 #( .INIT(16'h0ACC) )  
        \xhdl1.GEN_BITS[0].APB_32.INTR_reg_9_0_0[0]  (.A(INTR_reg_0), 
        .B(\INTR_reg_9_0_0_0_tz[0] ), .C(
        CoreAPB3_0_APBmslave2_PWDATA[0]), .D(edge_N_5_mux), .Y(
        \INTR_reg_9[0] ));
    CFG4 #( .INIT(16'hAC0F) )  
        \xhdl1.GEN_BITS[28].REG_GEN.CONFIG_reg[28]_RNII7LA2[5]  (.A(
        \CONFIG_reg[12][5] ), .B(\CONFIG_reg[28][5] ), .C(
        \CONFIG_reg_o_2_6_1_1[5] ), .D(CoreAPB3_0_APBmslave2_PADDR[5]), 
        .Y(N_4704));
    SLE \xhdl1.GEN_BITS[20].REG_GEN.CONFIG_reg[20][2]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[2]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[20]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[20][2] ));
    CFG3 #( .INIT(8'h04) )  
        \xhdl1.GEN_BITS[5].APB_32.INTR_reg_74_0_0_0_tz_1[5]  (.A(
        \CONFIG_reg[5][5] ), .B(\edge_both[5] ), .C(\CONFIG_reg[5][6] )
        , .Y(\INTR_reg_74_0_0_0_tz_1[5] ));
    SLE \xhdl1.GEN_BITS[29].REG_GEN.CONFIG_reg[29][1]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[1]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[29]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[29][1] ));
    CFG2 #( .INIT(4'h4) )  edge_neg_2_sqmuxa_7_i_a2 (.A(\gpin2[5] ), 
        .B(gpin3_5), .Y(N_405));
    CFG4 #( .INIT(16'h0F35) )  
        \xhdl1.GEN_BITS[2].REG_GEN.CONFIG_reg[2]_RNIG2I61[4]  (.A(
        \CONFIG_reg[2][4] ), .B(\CONFIG_reg[18][4] ), .C(
        CoreAPB3_0_APBmslave2_PADDR[6]), .D(
        CoreAPB3_0_APBmslave2_PADDR[5]), .Y(\CONFIG_reg_o_2_10_1_1[4] )
        );
    CFG4 #( .INIT(16'h0F35) )  
        \xhdl1.GEN_BITS[22].REG_GEN.CONFIG_reg[22]_RNI6P291[0]  (.A(
        \CONFIG_reg[6][0] ), .B(\CONFIG_reg[22][0] ), .C(
        CoreAPB3_0_APBmslave2_PADDR[6]), .D(
        CoreAPB3_0_APBmslave2_PADDR[5]), .Y(\CONFIG_reg_o_2_13_1_1[0] )
        );
    SLE \xhdl1.GEN_BITS[4].APB_32.edge_pos[4]  (.D(N_103), .CLK(
        FCCC_0_GL1), .EN(N_68), .ALn(MSS_RESET_N_F2M_c), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\edge_pos[4] ));
    CFG4 #( .INIT(16'h0F35) )  
        \xhdl1.GEN_BITS[17].REG_GEN.CONFIG_reg[17]_RNIA30K1[3]  (.A(
        \CONFIG_reg[1][3] ), .B(\CONFIG_reg[17][3] ), .C(
        CoreAPB3_0_APBmslave2_PADDR[6]), .D(
        CoreAPB3_0_APBmslave2_PADDR[5]), .Y(\CONFIG_reg_o_2_18_1[3] ));
    CFG3 #( .INIT(8'h20) )  
        \xhdl1.GEN_BITS[31].APB_32.edge_both_RNO[31]  (.A(
        \CONFIG_reg[31][3] ), .B(CoreAPB3_0_APBmslave2_PWDATA[31]), .C(
        \edge_pos[31] ), .Y(\edge_neg_443[31] ));
    CFG4 #( .INIT(16'hAC0F) )  
        \xhdl1.GEN_BITS[26].REG_GEN.CONFIG_reg[26]_RNI4MFS1[1]  (.A(
        \CONFIG_reg[10][1] ), .B(\CONFIG_reg[26][1] ), .C(
        \CONFIG_reg_o_2_10_1_1[1] ), .D(CoreAPB3_0_APBmslave2_PADDR[5])
        , .Y(N_4732));
    SLE \xhdl1.GEN_BITS[8].APB_32.edge_both[8]  (.D(\edge_neg_121[8] ), 
        .CLK(FCCC_0_GL1), .EN(edge_neg_2_sqmuxa_4_i_1), .ALn(
        MSS_RESET_N_F2M_c), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\edge_pos[8] ));
    CFG4 #( .INIT(16'hAC0F) )  
        \xhdl1.GEN_BITS[28].REG_GEN.CONFIG_reg[28]_RNIAVKA2[3]  (.A(
        \CONFIG_reg[12][3] ), .B(\CONFIG_reg[28][3] ), .C(
        \CONFIG_reg_o_2_6_1[3] ), .D(CoreAPB3_0_APBmslave2_PADDR[5]), 
        .Y(N_4702));
    SLE \xhdl1.GEN_BITS[0].REG_GEN.CONFIG_reg[0][3]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[3]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[0]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[0][3] ));
    SLE \xhdl1.GEN_BITS[23].REG_GEN.CONFIG_reg[23][1]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[1]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[23]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[23][1] ));
    SLE \xhdl1.GEN_BITS[13].REG_GEN.CONFIG_reg[13][3]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[3]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[13]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[13][3] ));
    CFG3 #( .INIT(8'hFB) )  edge_pos_2_sqmuxa_i_0 (.A(edge_N_5_mux), 
        .B(\CONFIG_reg[0][3] ), .C(N_402), .Y(N_74));
    CFG3 #( .INIT(8'hFB) )  edge_both_2_sqmuxa_11_i_0 (.A(edge_N_5_mux)
        , .B(\CONFIG_reg[4][3] ), .C(N_143_i), .Y(N_84));
    CFG3 #( .INIT(8'h20) )  
        \xhdl1.GEN_BITS[21].APB_32.edge_both_RNO[21]  (.A(
        \CONFIG_reg[21][3] ), .B(CoreAPB3_0_APBmslave2_PWDATA[21]), .C(
        \edge_neg[21] ), .Y(\edge_neg_303[21] ));
    CFG4 #( .INIT(16'h0F35) )  
        \xhdl1.GEN_BITS[20].REG_GEN.CONFIG_reg[20]_RNI45V31[3]  (.A(
        \CONFIG_reg[4][3] ), .B(\CONFIG_reg[20][3] ), .C(
        CoreAPB3_0_APBmslave2_PADDR[6]), .D(
        CoreAPB3_0_APBmslave2_PADDR[5]), .Y(\CONFIG_reg_o_2_6_1[3] ));
    SLE \xhdl1.GEN_BITS[18].REG_GEN.CONFIG_reg[18][7]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[7]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[18]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[18][7] ));
    CFG4 #( .INIT(16'h0F35) )  
        \xhdl1.GEN_BITS[17].REG_GEN.CONFIG_reg[17]_RNIG90K1[6]  (.A(
        \CONFIG_reg[1][6] ), .B(\CONFIG_reg[17][6] ), .C(
        CoreAPB3_0_APBmslave2_PADDR[6]), .D(
        CoreAPB3_0_APBmslave2_PADDR[5]), .Y(\CONFIG_reg_o_2_18_1_1[6] )
        );
    SLE \xhdl1.GEN_BITS[0].REG_GEN.CONFIG_reg[0][7]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[7]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[0]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[0][7] ));
    SLE \xhdl1.GEN_BITS[24].REG_GEN.CONFIG_reg[24][1]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[1]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[24]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[24][1] ));
    SLE \xhdl1.GEN_BITS[10].REG_GEN.CONFIG_reg[10][1]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[1]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[10]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[10][1] ));
    SLE \xhdl1.GEN_BITS[2].REG_GEN.CONFIG_reg[2][4]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[4]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[2]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[2][4] ));
    SLE \xhdl1.GEN_BITS[26].REG_GEN.CONFIG_reg[26][0]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[0]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[26]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[26][0] ));
    SLE \xhdl1.GEN_BITS[21].REG_GEN.CONFIG_reg[21][0]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[0]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[21]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[21][0] ));
    CFG4 #( .INIT(16'hA9FF) )  
        \xhdl1.GEN_BITS[20].APB_32.INTR_reg_269_0_o2_0_0[20]  (.A(
        \CONFIG_reg[20][7] ), .B(\CONFIG_reg[20][6] ), .C(
        \CONFIG_reg[20][5] ), .D(\CONFIG_reg[20][3] ), .Y(
        \INTR_reg_269_0_o2_0[20] ));
    CFG4 #( .INIT(16'h0F35) )  
        \xhdl1.GEN_BITS[19].REG_GEN.CONFIG_reg[19]_RNIM1491[5]  (.A(
        \CONFIG_reg[3][5] ), .B(\CONFIG_reg[19][5] ), .C(
        CoreAPB3_0_APBmslave2_PADDR[6]), .D(
        CoreAPB3_0_APBmslave2_PADDR[5]), .Y(\CONFIG_reg_o_2_25_1_1[5] )
        );
    CFG3 #( .INIT(8'hFB) )  edge_both_2_sqmuxa_12_i_0 (.A(edge_N_5_mux)
        , .B(\CONFIG_reg[3][3] ), .C(N_253_i), .Y(
        edge_both_2_sqmuxa_12_i_1));
    SLE \xhdl1.GEN_BITS[25].REG_GEN.CONFIG_reg[25][2]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[2]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[25]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[25][2] ));
    SLE \xhdl1.GEN_BITS[6].gpin3[6]  (.D(\gpin2[6] ), .CLK(FCCC_0_GL1), 
        .EN(VCC_net_1), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(gpin3_6));
    CFG4 #( .INIT(16'h0F35) )  
        \xhdl1.GEN_BITS[4].REG_GEN.CONFIG_reg[4]_RNI23V31[2]  (.A(
        \CONFIG_reg[4][2] ), .B(\CONFIG_reg[20][2] ), .C(
        CoreAPB3_0_APBmslave2_PADDR[6]), .D(
        CoreAPB3_0_APBmslave2_PADDR[5]), .Y(\CONFIG_reg_o_2_6_1_1[2] ));
    CFG4 #( .INIT(16'hAC0F) )  
        \xhdl1.GEN_BITS[29].REG_GEN.CONFIG_reg[29]_RNIU6J52[6]  (.A(
        \CONFIG_reg[13][6] ), .B(\CONFIG_reg[29][6] ), .C(
        \CONFIG_reg_o_2_21_1_1[6] ), .D(CoreAPB3_0_APBmslave2_PADDR[5])
        , .Y(N_4825));
    CFG4 #( .INIT(16'hC480) )  
        \xhdl1.GEN_BITS[1].APB_32.INTR_reg_22_0_0_0_tz[1]  (.A(
        \CONFIG_reg[1][7] ), .B(\CONFIG_reg[1][3] ), .C(
        \INTR_reg_22_0_0_0_tz_1[1] ), .D(N_177), .Y(
        \INTR_reg_22_0_0_0_tz[1] ));
    SLE \xhdl1.GEN_BITS[14].REG_GEN.CONFIG_reg[14][0]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[0]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[14]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[14][0] ));
    SLE \xhdl1.GEN_BITS[26].REG_GEN.CONFIG_reg[26][2]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[2]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[26]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[26][2] ));
    CFG2 #( .INIT(4'hB) )  edge_both_2_sqmuxa_16_i (.A(edge_N_5_mux), 
        .B(\CONFIG_reg[12][3] ), .Y(N_188));
    CFG4 #( .INIT(16'hA9FF) )  
        \xhdl1.GEN_BITS[31].APB_32.INTR_reg_412_0_o2_0_0[31]  (.A(
        \CONFIG_reg[31][7] ), .B(\CONFIG_reg[31][6] ), .C(
        \CONFIG_reg[31][5] ), .D(\CONFIG_reg[31][3] ), .Y(
        \INTR_reg_412_0_o2_0[31] ));
    SLE \xhdl1.GEN_BITS[23].REG_GEN.CONFIG_reg[23][6]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[6]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[23]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[23][6] ));
    CFG2 #( .INIT(4'h8) )  
        \xhdl1.GEN_BITS[3].REG_GPOUT.un34_GPIO_OUT_i  (.A(
        \GPOUT_reg[3] ), .B(\CONFIG_reg[3][0] ), .Y(GPIO_OUT_net_2[3]));
    CFG4 #( .INIT(16'hAC0F) )  
        \xhdl1.GEN_BITS[11].REG_GEN.CONFIG_reg[11]_RNIS1E72[5]  (.A(
        \CONFIG_reg[11][5] ), .B(\CONFIG_reg[27][5] ), .C(
        \CONFIG_reg_o_2_25_1_1[5] ), .D(CoreAPB3_0_APBmslave2_PADDR[5])
        , .Y(N_4856));
    CFG4 #( .INIT(16'hAC0F) )  
        \xhdl1.GEN_BITS[26].REG_GEN.CONFIG_reg[26]_RNI8QFS1[2]  (.A(
        \CONFIG_reg[10][2] ), .B(\CONFIG_reg[26][2] ), .C(
        \CONFIG_reg_o_2_10_1_1[2] ), .D(CoreAPB3_0_APBmslave2_PADDR[5])
        , .Y(N_4733));
    SLE \xhdl1.GEN_BITS[9].REG_GEN.CONFIG_reg[9][2]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[2]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[9]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[9][2] ));
    CFG4 #( .INIT(16'h0A33) )  
        \xhdl1.GEN_BITS[31].APB_32.INTR_reg_412_0[31]  (.A(INTR_reg_31)
        , .B(\INTR_reg_412_0_o2_1[31] ), .C(
        CoreAPB3_0_APBmslave2_PWDATA[31]), .D(edge_N_5_mux), .Y(
        \INTR_reg_412[31] ));
    SLE \xhdl1.GEN_BITS[5].REG_GEN.CONFIG_reg[5][5]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[5]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[5]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[5][5] ));
    CFG4 #( .INIT(16'hAC0F) )  
        \xhdl1.GEN_BITS[14].REG_GEN.CONFIG_reg[14]_RNIKCQ82[6]  (.A(
        \CONFIG_reg[14][6] ), .B(\CONFIG_reg[30][6] ), .C(
        \CONFIG_reg_o_2_13_1_1[6] ), .D(CoreAPB3_0_APBmslave2_PADDR[5])
        , .Y(N_4761));
    SLE \xhdl1.GEN_BITS[10].REG_GEN.CONFIG_reg[10][3]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[3]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[10]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[10][3] ));
    CFG3 #( .INIT(8'h04) )  
        \xhdl1.GEN_BITS[0].APB_32.INTR_reg_9_0_0_0_tz_1[0]  (.A(
        \CONFIG_reg[0][5] ), .B(\edge_both[0] ), .C(\CONFIG_reg[0][6] )
        , .Y(\INTR_reg_9_0_0_0_tz_1[0] ));
    SLE \xhdl1.GEN_BITS[23].APB_32.INTR_reg[23]  (.D(
        \INTR_reg_308[23] ), .CLK(FCCC_0_GL1), .EN(VCC_net_1), .ALn(
        MSS_RESET_N_F2M_c), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(INTR_reg_23));
    SLE \xhdl1.GEN_BITS[8].REG_GEN.CONFIG_reg[8][2]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[2]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[8]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[8][2] ));
    SLE \xhdl1.GEN_BITS[17].REG_GEN.CONFIG_reg[17][4]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[4]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[17]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[17][4] ));
    SLE \xhdl1.GEN_BITS[2].APB_32.edge_both[2]  (.D(N_93), .CLK(
        FCCC_0_GL1), .EN(N_86), .ALn(MSS_RESET_N_F2M_c), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\edge_both[2] ));
    SLE \xhdl1.GEN_BITS[1].gpin3[1]  (.D(\gpin2[1] ), .CLK(FCCC_0_GL1), 
        .EN(VCC_net_1), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(gpin3_1));
    CFG4 #( .INIT(16'h0ACC) )  
        \xhdl1.GEN_BITS[4].APB_32.INTR_reg_61_0_0[4]  (.A(INTR_reg_4), 
        .B(\INTR_reg_61_0_0_0_tz[4] ), .C(
        CoreAPB3_0_APBmslave2_PWDATA[4]), .D(edge_N_5_mux), .Y(
        \INTR_reg_61[4] ));
    SLE \xhdl1.GEN_BITS[20].REG_GEN.CONFIG_reg[20][0]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[0]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[20]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[20][0] ));
    SLE \xhdl1.GEN_BITS[23].REG_GEN.CONFIG_reg[23][2]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[2]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[23]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[23][2] ));
    SLE \xhdl1.GEN_BITS[4].REG_GEN.CONFIG_reg[4][5]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[5]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[4]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[4][5] ));
    SLE \xhdl1.GEN_BITS[2].REG_GEN.CONFIG_reg[2][6]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[6]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[2]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[2][6] ));
    CFG4 #( .INIT(16'hAA08) )  
        \xhdl1.GEN_BITS[4].APB_32.edge_pos_65_iv_i_0[4]  (.A(
        \CONFIG_reg[4][3] ), .B(\edge_pos[4] ), .C(
        CoreAPB3_0_APBmslave2_PWDATA[4]), .D(N_398), .Y(N_103));
    SLE \xhdl1.GEN_BITS[16].REG_GEN.CONFIG_reg[16][7]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[7]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[16]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[16][7] ));
    SLE \xhdl1.GEN_BITS[29].REG_GEN.CONFIG_reg[29][0]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[0]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[29]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[29][0] ));
    CFG4 #( .INIT(16'h4000) )  
        \xhdl1.GEN_BITS[9].REG_GEN.CONFIG_reg[9]2_0_a4_0_a2  (.A(
        CoreAPB3_0_APBmslave2_PADDR[3]), .B(
        CoreAPB3_0_APBmslave2_PADDR[2]), .C(N_604), .D(N_610), .Y(
        \CONFIG_reg[9]2 ));
    SLE \xhdl1.GEN_BITS[2].gpin3[2]  (.D(\gpin2[2] ), .CLK(FCCC_0_GL1), 
        .EN(VCC_net_1), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(gpin3_2));
    CFG3 #( .INIT(8'h20) )  
        \xhdl1.GEN_BITS[15].APB_32.edge_pos_RNO[15]  (.A(
        \CONFIG_reg[15][3] ), .B(CoreAPB3_0_APBmslave2_PWDATA[15]), .C(
        \edge_neg[15] ), .Y(\edge_pos_219[15] ));
    CFG4 #( .INIT(16'hAA08) )  
        \xhdl1.GEN_BITS[6].APB_32.edge_both_RNO[6]  (.A(
        \CONFIG_reg[6][3] ), .B(\edge_both[6] ), .C(
        CoreAPB3_0_APBmslave2_PWDATA[6]), .D(N_252_i), .Y(N_22_i_0));
    SLE \xhdl1.GEN_BITS[1].REG_GEN.CONFIG_reg[1][4]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[4]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[1]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[1][4] ));
    SLE \xhdl1.GEN_BITS[30].REG_GEN.CONFIG_reg[30][7]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[7]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[30]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[30][7] ));
    CFG4 #( .INIT(16'hAC0F) )  
        \xhdl1.GEN_BITS[15].REG_GEN.CONFIG_reg[15]_RNICNN32[2]  (.A(
        \CONFIG_reg[15][2] ), .B(\CONFIG_reg[31][2] ), .C(
        \CONFIG_reg_o_2_28_1_1[2] ), .D(CoreAPB3_0_APBmslave2_PADDR[5])
        , .Y(N_4877));
    CFG4 #( .INIT(16'hAC0F) )  
        \xhdl1.GEN_BITS[9].REG_GEN.CONFIG_reg[9]_RNIIMU72[2]  (.A(
        \CONFIG_reg[9][2] ), .B(\CONFIG_reg[25][2] ), .C(
        \CONFIG_reg_o_2_18_1_1[2] ), .D(CoreAPB3_0_APBmslave2_PADDR[5])
        , .Y(N_4797));
    CFG4 #( .INIT(16'h0A33) )  
        \xhdl1.GEN_BITS[23].APB_32.INTR_reg_308_0[23]  (.A(INTR_reg_23)
        , .B(\INTR_reg_308_0_o2_1[23] ), .C(
        CoreAPB3_0_APBmslave2_PWDATA[23]), .D(edge_N_5_mux), .Y(
        \INTR_reg_308[23] ));
    CFG4 #( .INIT(16'hAC0F) )  
        \xhdl1.GEN_BITS[9].REG_GEN.CONFIG_reg[9]_RNIQUU72[4]  (.A(
        \CONFIG_reg[9][4] ), .B(\CONFIG_reg[25][4] ), .C(
        \CONFIG_reg_o_2_18_1[4] ), .D(CoreAPB3_0_APBmslave2_PADDR[5]), 
        .Y(N_4799));
    SLE \xhdl1.GEN_BITS[19].REG_GEN.CONFIG_reg[19][1]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[1]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[19]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[19][1] ));
    SLE \xhdl1.GEN_BITS[3].REG_GEN.CONFIG_reg[3][2]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[2]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[3]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[3][2] ));
    CFG4 #( .INIT(16'h0F35) )  
        \xhdl1.GEN_BITS[2].REG_GEN.CONFIG_reg[2]_RNIK6I61[6]  (.A(
        \CONFIG_reg[2][6] ), .B(\CONFIG_reg[18][6] ), .C(
        CoreAPB3_0_APBmslave2_PADDR[6]), .D(
        CoreAPB3_0_APBmslave2_PADDR[5]), .Y(\CONFIG_reg_o_2_10_1_1[6] )
        );
    SLE \xhdl1.GEN_BITS[12].REG_GEN.CONFIG_reg[12][0]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[0]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[12]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[12][0] ));
    SLE \xhdl1.GEN_BITS[7].REG_GEN.CONFIG_reg[7][5]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[5]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[7]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[7][5] ));
    CFG4 #( .INIT(16'hAA08) )  
        \xhdl1.GEN_BITS[2].APB_32.edge_pos_37_iv_i_0[2]  (.A(
        \CONFIG_reg[2][3] ), .B(\edge_pos[2] ), .C(
        CoreAPB3_0_APBmslave2_PWDATA[2]), .D(N_396), .Y(N_105));
    CFG4 #( .INIT(16'h0A33) )  
        \xhdl1.GEN_BITS[26].APB_32.INTR_reg_347_0[26]  (.A(INTR_reg_26)
        , .B(\INTR_reg_347_0_o2_1[26] ), .C(
        CoreAPB3_0_APBmslave2_PWDATA[26]), .D(edge_N_5_mux), .Y(
        \INTR_reg_347[26] ));
    CFG4 #( .INIT(16'h4000) )  
        \xhdl1.GEN_BITS[6].REG_GEN.CONFIG_reg[6]2_0_a4_0_a2  (.A(
        CoreAPB3_0_APBmslave2_PADDR[2]), .B(
        CoreAPB3_0_APBmslave2_PADDR[3]), .C(N_603), .D(N_604), .Y(
        \CONFIG_reg[6]2 ));
    SLE \xhdl1.GEN_BITS[24].APB_32.edge_both[24]  (.D(N_100_i_0), .CLK(
        FCCC_0_GL1), .EN(N_155), .ALn(MSS_RESET_N_F2M_c), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\edge_pos[24] ));
    CFG3 #( .INIT(8'hFE) )  
        \xhdl1.GEN_BITS[0].REG_GEN.CONFIG_reg[0]2_0_a4_0_o2  (.A(
        CoreAPB3_0_APBmslave2_PADDR[2]), .B(
        CoreAPB3_0_APBmslave2_PADDR[3]), .C(
        CoreAPB3_0_APBmslave2_PADDR[6]), .Y(N_243));
    CFG4 #( .INIT(16'h4000) )  
        \xhdl1.GEN_BITS[21].REG_GEN.CONFIG_reg[21]2_0_a4_0_a2  (.A(
        CoreAPB3_0_APBmslave2_PADDR[3]), .B(
        CoreAPB3_0_APBmslave2_PADDR[2]), .C(N_598), .D(N_603), .Y(
        \CONFIG_reg[21]2 ));
    CFG4 #( .INIT(16'hAC0F) )  
        \xhdl1.GEN_BITS[29].REG_GEN.CONFIG_reg[29]_RNIMUI52[4]  (.A(
        \CONFIG_reg[13][4] ), .B(\CONFIG_reg[29][4] ), .C(
        \CONFIG_reg_o_2_21_1[4] ), .D(CoreAPB3_0_APBmslave2_PADDR[5]), 
        .Y(N_4823));
    SLE \xhdl1.GEN_BITS[11].REG_GEN.CONFIG_reg[11][3]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[3]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[11]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[11][3] ));
    SLE \xhdl1.GEN_BITS[3].APB_32.GPOUT_reg[3]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[3]), .CLK(FCCC_0_GL1), .EN(
        GPOUT_reg_0_sqmuxa), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \GPOUT_reg[3] ));
    SLE \xhdl1.GEN_BITS[30].REG_GEN.CONFIG_reg[30][6]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[6]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[30]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[30][6] ));
    CFG3 #( .INIT(8'hFB) )  edge_pos_2_sqmuxa_18_i_0 (.A(edge_N_5_mux), 
        .B(\CONFIG_reg[3][3] ), .C(N_687), .Y(N_79));
    CFG4 #( .INIT(16'h0A33) )  
        \xhdl1.GEN_BITS[19].APB_32.INTR_reg_256_0[19]  (.A(INTR_reg_19)
        , .B(\INTR_reg_256_0_o2_1[19] ), .C(
        CoreAPB3_0_APBmslave2_PWDATA[19]), .D(edge_N_5_mux), .Y(
        \INTR_reg_256[19] ));
    SLE \xhdl1.GEN_BITS[5].APB_32.edge_both[5]  (.D(N_89), .CLK(
        FCCC_0_GL1), .EN(N_76), .ALn(MSS_RESET_N_F2M_c), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\edge_both[5] ));
    SLE \xhdl1.GEN_BITS[19].APB_32.INTR_reg[19]  (.D(
        \INTR_reg_256[19] ), .CLK(FCCC_0_GL1), .EN(VCC_net_1), .ALn(
        MSS_RESET_N_F2M_c), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(INTR_reg_19));
    SLE \xhdl1.GEN_BITS[1].REG_GEN.CONFIG_reg[1][6]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[6]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[1]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[1][6] ));
    CFG3 #( .INIT(8'hFB) )  edge_neg_2_sqmuxa_7_i_0 (.A(edge_N_5_mux), 
        .B(\CONFIG_reg[5][3] ), .C(N_405), .Y(N_60));
    SLE \xhdl1.GEN_BITS[15].APB_32.INTR_reg[15]  (.D(
        \INTR_reg_204[15] ), .CLK(FCCC_0_GL1), .EN(VCC_net_1), .ALn(
        MSS_RESET_N_F2M_c), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(INTR_reg_15));
    SLE \xhdl1.GEN_BITS[16].APB_32.INTR_reg[16]  (.D(
        \INTR_reg_217[16] ), .CLK(FCCC_0_GL1), .EN(VCC_net_1), .ALn(
        MSS_RESET_N_F2M_c), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(INTR_reg_16));
    SLE \xhdl1.GEN_BITS[6].REG_GEN.CONFIG_reg[6][2]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[2]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[6]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[6][2] ));
    SLE \xhdl1.GEN_BITS[19].REG_GEN.CONFIG_reg[19][3]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[3]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[19]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[19][3] ));
    CFG2 #( .INIT(4'h8) )  
        \xhdl1.GEN_BITS[14].REG_GEN.CONFIG_reg[14]2_0_a4_0_a2_0  (.A(
        CoreAPB3_0_APBmslave2_PADDR[5]), .B(
        CoreAPB3_0_APBmslave2_PADDR[4]), .Y(N_605));
    CFG4 #( .INIT(16'h0F35) )  
        \xhdl1.GEN_BITS[7].REG_GEN.CONFIG_reg[7]_RNIK0LB1[5]  (.A(
        \CONFIG_reg[7][5] ), .B(\CONFIG_reg[23][5] ), .C(
        CoreAPB3_0_APBmslave2_PADDR[6]), .D(
        CoreAPB3_0_APBmslave2_PADDR[5]), .Y(\CONFIG_reg_o_2_28_1_1[5] )
        );
    SLE \xhdl1.GEN_BITS[21].REG_GEN.CONFIG_reg[21][6]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[6]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[21]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[21][6] ));
    SLE \xhdl1.GEN_BITS[14].REG_GEN.CONFIG_reg[14][5]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[5]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[14]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[14][5] ));
    CFG2 #( .INIT(4'h4) )  edge_neg_2_sqmuxa_11_i_a2 (.A(\gpin2[1] ), 
        .B(gpin3_1), .Y(N_399));
    CFG3 #( .INIT(8'hFB) )  edge_pos_2_sqmuxa_6_i_0 (.A(edge_N_5_mux), 
        .B(\CONFIG_reg[2][3] ), .C(N_396), .Y(N_64));
    CFG4 #( .INIT(16'hAA08) )  
        \xhdl1.GEN_BITS[4].APB_32.edge_neg_65_iv_i_0[4]  (.A(
        \CONFIG_reg[4][3] ), .B(\edge_neg[4] ), .C(
        CoreAPB3_0_APBmslave2_PWDATA[4]), .D(N_397), .Y(N_117));
    CFG2 #( .INIT(4'hB) )  edge_both_2_sqmuxa_3_i (.A(edge_N_5_mux), 
        .B(\CONFIG_reg[16][3] ), .Y(edge_pos_2_sqmuxa_29_i_1));
    CFG4 #( .INIT(16'hAA08) )  
        \xhdl1.GEN_BITS[2].APB_32.edge_neg_37_iv_i_0[2]  (.A(
        \CONFIG_reg[2][3] ), .B(\edge_neg[2] ), .C(
        CoreAPB3_0_APBmslave2_PWDATA[2]), .D(N_395), .Y(N_119));
    CFG3 #( .INIT(8'h20) )  
        \xhdl1.GEN_BITS[16].APB_32.edge_both_RNO[16]  (.A(
        \CONFIG_reg[16][3] ), .B(CoreAPB3_0_APBmslave2_PWDATA[16]), .C(
        \edge_neg[16] ), .Y(\edge_neg_233[16] ));
    SLE \xhdl1.GEN_BITS[2].REG_GEN.CONFIG_reg[2][0]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[0]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[2]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[2][0] ));
    SLE \xhdl1.GEN_BITS[21].REG_GEN.CONFIG_reg[21][4]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[4]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[21]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[21][4] ));
    CFG4 #( .INIT(16'hF2F3) )  
        \xhdl1.GEN_BITS[12].APB_32.INTR_reg_165_0_o2_1_0[12]  (.A(
        \CONFIG_reg[12][6] ), .B(\edge_neg[12] ), .C(
        \INTR_reg_165_0_o2_0[12] ), .D(\CONFIG_reg[12][5] ), .Y(
        \INTR_reg_165_0_o2_1[12] ));
    SLE \xhdl1.GEN_BITS[30].REG_GEN.CONFIG_reg[30][4]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[4]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[30]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[30][4] ));
    SLE \xhdl1.GEN_BITS[28].REG_GEN.CONFIG_reg[28][0]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[0]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[28]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[28][0] ));
    CFG4 #( .INIT(16'h0F35) )  
        \xhdl1.GEN_BITS[16].REG_GEN.CONFIG_reg[16]_RNICCE11[6]  (.A(
        \CONFIG_reg[0][6] ), .B(\CONFIG_reg[16][6] ), .C(
        CoreAPB3_0_APBmslave2_PADDR[6]), .D(
        CoreAPB3_0_APBmslave2_PADDR[5]), .Y(\CONFIG_reg_o_2_3_1_1[6] ));
    SLE \xhdl1.GEN_BITS[22].APB_32.INTR_reg[22]  (.D(
        \INTR_reg_295[22] ), .CLK(FCCC_0_GL1), .EN(VCC_net_1), .ALn(
        MSS_RESET_N_F2M_c), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(INTR_reg_22));
    CFG2 #( .INIT(4'h4) )  edge_neg_2_sqmuxa_9_i_a2 (.A(\gpin2[3] ), 
        .B(gpin3_3), .Y(N_686));
    SLE \xhdl1.GEN_BITS[1].APB_32.INTR_reg[1]  (.D(\INTR_reg_22[1] ), 
        .CLK(FCCC_0_GL1), .EN(VCC_net_1), .ALn(MSS_RESET_N_F2M_c), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(INTR_reg_1));
    CFG4 #( .INIT(16'hAC0F) )  
        \xhdl1.GEN_BITS[26].REG_GEN.CONFIG_reg[26]_RNISEGS1[7]  (.A(
        \CONFIG_reg[10][7] ), .B(\CONFIG_reg[26][7] ), .C(
        \CONFIG_reg_o_2_10_1_1[7] ), .D(CoreAPB3_0_APBmslave2_PADDR[5])
        , .Y(N_4738));
    SLE \xhdl1.GEN_BITS[14].APB_32.GPOUT_reg[14]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[14]), .CLK(FCCC_0_GL1), .EN(
        GPOUT_reg_0_sqmuxa), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        GPOUT_reg_14));
    CFG4 #( .INIT(16'h0F35) )  
        \xhdl1.GEN_BITS[19].REG_GEN.CONFIG_reg[19]_RNIO3491[6]  (.A(
        \CONFIG_reg[3][6] ), .B(\CONFIG_reg[19][6] ), .C(
        CoreAPB3_0_APBmslave2_PADDR[6]), .D(
        CoreAPB3_0_APBmslave2_PADDR[5]), .Y(\CONFIG_reg_o_2_25_1_1[6] )
        );
    CFG4 #( .INIT(16'hAC0F) )  
        \xhdl1.GEN_BITS[15].REG_GEN.CONFIG_reg[15]_RNIO3O32[5]  (.A(
        \CONFIG_reg[15][5] ), .B(\CONFIG_reg[31][5] ), .C(
        \CONFIG_reg_o_2_28_1_1[5] ), .D(CoreAPB3_0_APBmslave2_PADDR[5])
        , .Y(N_4880));
    SLE \xhdl1.GEN_BITS[24].REG_GEN.CONFIG_reg[24][6]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[6]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[24]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[24][6] ));
    SLE \xhdl1.GEN_BITS[16].REG_GEN.CONFIG_reg[16][0]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[0]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[16]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[16][0] ));
    CFG4 #( .INIT(16'hF2F3) )  
        \xhdl1.GEN_BITS[22].APB_32.INTR_reg_295_0_o2_1_0[22]  (.A(
        \CONFIG_reg[22][6] ), .B(\edge_neg[22] ), .C(
        \INTR_reg_295_0_o2_0[22] ), .D(\CONFIG_reg[22][5] ), .Y(
        \INTR_reg_295_0_o2_1[22] ));
    CFG4 #( .INIT(16'h0F35) )  
        \xhdl1.GEN_BITS[22].REG_GEN.CONFIG_reg[22]_RNIK7391[7]  (.A(
        \CONFIG_reg[6][7] ), .B(\CONFIG_reg[22][7] ), .C(
        CoreAPB3_0_APBmslave2_PADDR[6]), .D(
        CoreAPB3_0_APBmslave2_PADDR[5]), .Y(\CONFIG_reg_o_2_13_1_1[7] )
        );
    CFG4 #( .INIT(16'hAA08) )  
        \xhdl1.GEN_BITS[3].APB_32.edge_both_51_iv_i[3]  (.A(
        \CONFIG_reg[3][3] ), .B(\edge_both[3] ), .C(
        CoreAPB3_0_APBmslave2_PWDATA[3]), .D(N_253_i), .Y(
        \edge_both_51_iv_i_0[3] ));
    SLE \xhdl1.GEN_BITS[9].APB_32.GPOUT_reg[9]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[9]), .CLK(FCCC_0_GL1), .EN(
        GPOUT_reg_0_sqmuxa), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        GPOUT_reg_9));
    CFG4 #( .INIT(16'hAA08) )  
        \xhdl1.GEN_BITS[4].APB_32.edge_both_65_iv_i_0[4]  (.A(
        \CONFIG_reg[4][3] ), .B(\edge_both[4] ), .C(
        CoreAPB3_0_APBmslave2_PWDATA[4]), .D(N_143_i), .Y(N_91));
    CFG4 #( .INIT(16'h0F35) )  
        \xhdl1.GEN_BITS[16].REG_GEN.CONFIG_reg[16]_RNI66E11[3]  (.A(
        \CONFIG_reg[0][3] ), .B(\CONFIG_reg[16][3] ), .C(
        CoreAPB3_0_APBmslave2_PADDR[6]), .D(
        CoreAPB3_0_APBmslave2_PADDR[5]), .Y(\CONFIG_reg_o_2_3_1[3] ));
    SLE \xhdl1.GEN_BITS[15].APB_32.GPOUT_reg[15]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[15]), .CLK(FCCC_0_GL1), .EN(
        GPOUT_reg_0_sqmuxa), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        GPOUT_reg_15));
    CFG4 #( .INIT(16'h0F35) )  
        \xhdl1.GEN_BITS[7].REG_GEN.CONFIG_reg[7]_RNIO4LB1[7]  (.A(
        \CONFIG_reg[7][7] ), .B(\CONFIG_reg[23][7] ), .C(
        CoreAPB3_0_APBmslave2_PADDR[6]), .D(
        CoreAPB3_0_APBmslave2_PADDR[5]), .Y(\CONFIG_reg_o_2_28_1_1[7] )
        );
    CFG4 #( .INIT(16'hAC0F) )  
        \xhdl1.GEN_BITS[9].REG_GEN.CONFIG_reg[9]_RNIU2V72[5]  (.A(
        \CONFIG_reg[9][5] ), .B(\CONFIG_reg[25][5] ), .C(
        \CONFIG_reg_o_2_18_1_1[5] ), .D(CoreAPB3_0_APBmslave2_PADDR[5])
        , .Y(N_4800));
    SLE \xhdl1.GEN_BITS[24].REG_GEN.CONFIG_reg[24][0]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[0]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[24]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[24][0] ));
    SLE \xhdl1.GEN_BITS[17].REG_GEN.CONFIG_reg[17][6]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[6]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[17]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[17][6] ));
    CFG3 #( .INIT(8'h04) )  
        \xhdl1.GEN_BITS[1].APB_32.INTR_reg_22_0_0_0_tz_1[1]  (.A(
        \CONFIG_reg[1][5] ), .B(\edge_both[1] ), .C(\CONFIG_reg[1][6] )
        , .Y(\INTR_reg_22_0_0_0_tz_1[1] ));
    CFG3 #( .INIT(8'hFB) )  edge_pos_2_sqmuxa_2_i_0_0 (.A(edge_N_5_mux)
        , .B(\CONFIG_reg[6][3] ), .C(N_689), .Y(N_72));
    CFG4 #( .INIT(16'hC480) )  
        \xhdl1.GEN_BITS[4].APB_32.INTR_reg_61_0_0_0_tz[4]  (.A(
        \CONFIG_reg[4][7] ), .B(\CONFIG_reg[4][3] ), .C(
        \INTR_reg_61_0_0_0_tz_1[4] ), .D(N_179), .Y(
        \INTR_reg_61_0_0_0_tz[4] ));
    SLE \xhdl1.GEN_BITS[19].REG_GEN.CONFIG_reg[19][4]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[4]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[19]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[19][4] ));
    CFG2 #( .INIT(4'h8) )  
        \xhdl1.GEN_BITS[6].REG_GPOUT.un64_GPIO_OUT_i  (.A(GPOUT_reg_6), 
        .B(\CONFIG_reg[6][0] ), .Y(GPIO_OUT_net_2[6]));
    SLE \xhdl1.GEN_BITS[9].APB_32.INTR_reg[9]  (.D(\INTR_reg_126[9] ), 
        .CLK(FCCC_0_GL1), .EN(VCC_net_1), .ALn(MSS_RESET_N_F2M_c), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(INTR_reg_9));
    CFG4 #( .INIT(16'hAC0F) )  
        \xhdl1.GEN_BITS[29].REG_GEN.CONFIG_reg[29]_RNI2BJ52[7]  (.A(
        \CONFIG_reg[13][7] ), .B(\CONFIG_reg[29][7] ), .C(
        \CONFIG_reg_o_2_21_1_1[7] ), .D(CoreAPB3_0_APBmslave2_PADDR[5])
        , .Y(N_4826));
    CFG4 #( .INIT(16'h0A33) )  
        \xhdl1.GEN_BITS[27].APB_32.INTR_reg_360_0[27]  (.A(INTR_reg_27)
        , .B(\INTR_reg_360_0_o2_1[27] ), .C(
        CoreAPB3_0_APBmslave2_PWDATA[27]), .D(edge_N_5_mux), .Y(
        \INTR_reg_360[27] ));
    SLE \xhdl1.GEN_BITS[1].REG_GEN.CONFIG_reg[1][0]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[0]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[1]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[1][0] ));
    CFG2 #( .INIT(4'h4) )  edge_neg_2_sqmuxa_25_i_a2 (.A(\gpin2[0] ), 
        .B(gpin3_0), .Y(N_401));
    CFG4 #( .INIT(16'hC5CA) )  
        \xhdl1.GEN_BITS[2].APB_32.INTR_reg_35_0_m2[2]  (.A(gpin3_2), 
        .B(N_173), .C(\CONFIG_reg[2][6] ), .D(\CONFIG_reg[2][5] ), .Y(
        N_178));
    CFG4 #( .INIT(16'hAC0F) )  
        \xhdl1.GEN_BITS[11].REG_GEN.CONFIG_reg[11]_RNI06E72[6]  (.A(
        \CONFIG_reg[11][6] ), .B(\CONFIG_reg[27][6] ), .C(
        \CONFIG_reg_o_2_25_1_1[6] ), .D(CoreAPB3_0_APBmslave2_PADDR[5])
        , .Y(N_4857));
    SLE \xhdl1.GEN_BITS[20].APB_32.GPOUT_reg[20]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[20]), .CLK(FCCC_0_GL1), .EN(
        GPOUT_reg_0_sqmuxa), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        GPOUT_reg_20));
    SLE \xhdl1.GEN_BITS[29].APB_32.GPOUT_reg[29]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[29]), .CLK(FCCC_0_GL1), .EN(
        GPOUT_reg_0_sqmuxa), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        GPOUT_reg_29));
    CFG4 #( .INIT(16'h0F35) )  
        \xhdl1.GEN_BITS[7].REG_GEN.CONFIG_reg[7]_RNIM2LB1[6]  (.A(
        \CONFIG_reg[7][6] ), .B(\CONFIG_reg[23][6] ), .C(
        CoreAPB3_0_APBmslave2_PADDR[6]), .D(
        CoreAPB3_0_APBmslave2_PADDR[5]), .Y(\CONFIG_reg_o_2_28_1_1[6] )
        );
    CFG2 #( .INIT(4'h8) )  
        \xhdl1.GEN_BITS[4].REG_GPOUT.un44_GPIO_OUT_i  (.A(GPOUT_reg_4), 
        .B(\CONFIG_reg[4][0] ), .Y(GPIO_OUT_net_2[4]));
    CFG4 #( .INIT(16'hAA08) )  
        \xhdl1.GEN_BITS[5].APB_32.edge_both_79_iv_i_0[5]  (.A(
        \CONFIG_reg[5][3] ), .B(\edge_both[5] ), .C(
        CoreAPB3_0_APBmslave2_PWDATA[5]), .D(N_139_i), .Y(N_89));
    CFG4 #( .INIT(16'hAC0F) )  
        \xhdl1.GEN_BITS[24].REG_GEN.CONFIG_reg[24]_RNI6OQ22[1]  (.A(
        \CONFIG_reg[8][1] ), .B(\CONFIG_reg[24][1] ), .C(
        \CONFIG_reg_o_2_3_1_1[1] ), .D(CoreAPB3_0_APBmslave2_PADDR[5]), 
        .Y(N_4676));
    SLE \xhdl1.GEN_BITS[24].REG_GEN.CONFIG_reg[24][3]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[3]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[24]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[24][3] ));
    CFG4 #( .INIT(16'hAC0F) )  
        \xhdl1.GEN_BITS[11].REG_GEN.CONFIG_reg[11]_RNI8DD72[0]  (.A(
        \CONFIG_reg[11][0] ), .B(\CONFIG_reg[27][0] ), .C(
        \CONFIG_reg_o_2_25_1_1[0] ), .D(CoreAPB3_0_APBmslave2_PADDR[5])
        , .Y(N_4851));
    SLE \xhdl1.GEN_BITS[10].APB_32.GPOUT_reg[10]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[10]), .CLK(FCCC_0_GL1), .EN(
        GPOUT_reg_0_sqmuxa), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        GPOUT_reg_10));
    SLE \xhdl1.GEN_BITS[16].REG_GEN.CONFIG_reg[16][1]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[1]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[16]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[16][1] ));
    SLE \xhdl1.GEN_BITS[14].REG_GEN.CONFIG_reg[14][4]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[4]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[14]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[14][4] ));
    SLE \xhdl1.GEN_BITS[7].APB_32.GPOUT_reg[7]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[7]), .CLK(FCCC_0_GL1), .EN(
        GPOUT_reg_0_sqmuxa), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \GPOUT_reg[7] ));
    SLE \xhdl1.GEN_BITS[18].REG_GEN.CONFIG_reg[18][0]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[0]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[18]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[18][0] ));
    CFG4 #( .INIT(16'h0F35) )  
        \xhdl1.GEN_BITS[7].REG_GEN.CONFIG_reg[7]_RNICOKB1[1]  (.A(
        \CONFIG_reg[7][1] ), .B(\CONFIG_reg[23][1] ), .C(
        CoreAPB3_0_APBmslave2_PADDR[6]), .D(
        CoreAPB3_0_APBmslave2_PADDR[5]), .Y(\CONFIG_reg_o_2_28_1_1[1] )
        );
    CFG4 #( .INIT(16'hAC0F) )  
        \xhdl1.GEN_BITS[9].REG_GEN.CONFIG_reg[9]_RNIEIU72[1]  (.A(
        \CONFIG_reg[9][1] ), .B(\CONFIG_reg[25][1] ), .C(
        \CONFIG_reg_o_2_18_1_1[1] ), .D(CoreAPB3_0_APBmslave2_PADDR[5])
        , .Y(N_4796));
    SLE \xhdl1.GEN_BITS[5].REG_GEN.CONFIG_reg[5][3]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[3]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[5]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[5][3] ));
    CFG4 #( .INIT(16'hAC0F) )  
        \xhdl1.GEN_BITS[28].REG_GEN.CONFIG_reg[28]_RNIQFLA2[7]  (.A(
        \CONFIG_reg[12][7] ), .B(\CONFIG_reg[28][7] ), .C(
        \CONFIG_reg_o_2_6_1_1[7] ), .D(CoreAPB3_0_APBmslave2_PADDR[5]), 
        .Y(N_4706));
    CFG4 #( .INIT(16'h8000) )  
        \xhdl1.GEN_BITS[19].REG_GEN.CONFIG_reg[19]2_0_a4_0_a2  (.A(
        CoreAPB3_0_APBmslave2_PADDR[3]), .B(
        CoreAPB3_0_APBmslave2_PADDR[2]), .C(N_598), .D(N_606), .Y(
        \CONFIG_reg[19]2 ));
    CFG4 #( .INIT(16'h0F35) )  
        \xhdl1.GEN_BITS[2].REG_GEN.CONFIG_reg[2]_RNICUH61[2]  (.A(
        \CONFIG_reg[2][2] ), .B(\CONFIG_reg[18][2] ), .C(
        CoreAPB3_0_APBmslave2_PADDR[6]), .D(
        CoreAPB3_0_APBmslave2_PADDR[5]), .Y(\CONFIG_reg_o_2_10_1_1[2] )
        );
    CFG4 #( .INIT(16'hAC0F) )  
        \xhdl1.GEN_BITS[26].REG_GEN.CONFIG_reg[26]_RNICUFS1[3]  (.A(
        \CONFIG_reg[10][3] ), .B(\CONFIG_reg[26][3] ), .C(
        \CONFIG_reg_o_2_10_1_1[3] ), .D(CoreAPB3_0_APBmslave2_PADDR[5])
        , .Y(N_4734));
    SLE \xhdl1.GEN_BITS[5].REG_GEN.CONFIG_reg[5][7]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[7]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[5]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[5][7] ));
    CFG2 #( .INIT(4'hB) )  edge_both_2_sqmuxa_30_i (.A(edge_N_5_mux), 
        .B(\CONFIG_reg[25][3] ), .Y(N_157));
    SLE \xhdl1.GEN_BITS[3].gpin3[3]  (.D(\gpin2[3] ), .CLK(FCCC_0_GL1), 
        .EN(VCC_net_1), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(gpin3_3));
    CFG4 #( .INIT(16'h0A33) )  
        \xhdl1.GEN_BITS[18].APB_32.INTR_reg_243_0[18]  (.A(INTR_reg_18)
        , .B(\INTR_reg_243_0_o2_1[18] ), .C(
        CoreAPB3_0_APBmslave2_PWDATA[18]), .D(edge_N_5_mux), .Y(
        \INTR_reg_243[18] ));
    CFG4 #( .INIT(16'h2000) )  
        \xhdl1.GEN_BITS[10].REG_GEN.CONFIG_reg[10]2_0_a4_0_a2  (.A(
        CoreAPB3_0_APBmslave2_PADDR[3]), .B(
        CoreAPB3_0_APBmslave2_PADDR[2]), .C(N_604), .D(N_610), .Y(
        \CONFIG_reg[10]2 ));
    CFG2 #( .INIT(4'hB) )  edge_both_2_sqmuxa_4_i (.A(edge_N_5_mux), 
        .B(\CONFIG_reg[15][3] ), .Y(edge_pos_2_sqmuxa_7_i_1));
    SLE \xhdl1.GEN_BITS[4].REG_GEN.CONFIG_reg[4][3]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[3]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[4]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[4][3] ));
    SLE \xhdl1.GEN_BITS[9].REG_GEN.CONFIG_reg[9][5]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[5]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[9]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[9][5] ));
    SLE \xhdl1.GEN_BITS[29].REG_GEN.CONFIG_reg[29][5]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[5]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[29]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[29][5] ));
    CFG4 #( .INIT(16'hF2F3) )  
        \xhdl1.GEN_BITS[27].APB_32.INTR_reg_360_0_o2_1_0[27]  (.A(
        \CONFIG_reg[27][6] ), .B(\edge_neg[27] ), .C(
        \INTR_reg_360_0_o2_0[27] ), .D(\CONFIG_reg[27][5] ), .Y(
        \INTR_reg_360_0_o2_1[27] ));
    SLE \xhdl1.GEN_BITS[26].REG_GEN.CONFIG_reg[26][1]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[1]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[26]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[26][1] ));
    SLE \xhdl1.GEN_BITS[22].APB_32.GPOUT_reg[22]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[22]), .CLK(FCCC_0_GL1), .EN(
        GPOUT_reg_0_sqmuxa), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        GPOUT_reg_22));
    CFG2 #( .INIT(4'hB) )  edge_both_2_sqmuxa_20_i (.A(edge_N_5_mux), 
        .B(\CONFIG_reg[8][3] ), .Y(edge_neg_2_sqmuxa_4_i_1));
    SLE \xhdl1.GEN_BITS[27].APB_32.GPOUT_reg[27]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[27]), .CLK(FCCC_0_GL1), .EN(
        GPOUT_reg_0_sqmuxa), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        GPOUT_reg_27));
    SLE \xhdl1.GEN_BITS[31].APB_32.edge_both[31]  (.D(
        \edge_neg_443[31] ), .CLK(FCCC_0_GL1), .EN(
        edge_pos_2_sqmuxa_19_i_1), .ALn(MSS_RESET_N_F2M_c), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\edge_pos[31] ));
    CFG3 #( .INIT(8'h20) )  
        \xhdl1.GEN_BITS[14].APB_32.edge_both_RNO[14]  (.A(
        \CONFIG_reg[14][3] ), .B(CoreAPB3_0_APBmslave2_PWDATA[14]), .C(
        \edge_neg[14] ), .Y(\edge_neg_205[14] ));
    SLE \xhdl1.GEN_BITS[8].REG_GEN.CONFIG_reg[8][5]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[5]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[8]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[8][5] ));
    CFG4 #( .INIT(16'h2000) )  
        \xhdl1.GEN_BITS[26].REG_GEN.CONFIG_reg[26]2_0_a4_0_a2  (.A(
        CoreAPB3_0_APBmslave2_PADDR[3]), .B(
        CoreAPB3_0_APBmslave2_PADDR[2]), .C(N_598), .D(N_610), .Y(
        \CONFIG_reg[26]2 ));
    SLE \xhdl1.GEN_BITS[13].REG_GEN.CONFIG_reg[13][5]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[5]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[13]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[13][5] ));
    CFG4 #( .INIT(16'hAA08) )  
        \xhdl1.GEN_BITS[6].APB_32.edge_neg_93_iv_i_0_0[6]  (.A(
        \CONFIG_reg[6][3] ), .B(\edge_neg[6] ), .C(
        CoreAPB3_0_APBmslave2_PWDATA[6]), .D(N_688), .Y(N_113));
    CFG4 #( .INIT(16'hA9FF) )  
        \xhdl1.GEN_BITS[11].APB_32.INTR_reg_152_0_o2_0_0[11]  (.A(
        \CONFIG_reg[11][7] ), .B(\CONFIG_reg[11][6] ), .C(
        \CONFIG_reg[11][5] ), .D(\CONFIG_reg[11][3] ), .Y(
        \INTR_reg_152_0_o2_0[11] ));
    SLE \xhdl1.GEN_BITS[4].REG_GEN.CONFIG_reg[4][7]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[7]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[4]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[4][7] ));
    CFG4 #( .INIT(16'h0F35) )  
        \xhdl1.GEN_BITS[22].REG_GEN.CONFIG_reg[22]_RNII5391[6]  (.A(
        \CONFIG_reg[6][6] ), .B(\CONFIG_reg[22][6] ), .C(
        CoreAPB3_0_APBmslave2_PADDR[6]), .D(
        CoreAPB3_0_APBmslave2_PADDR[5]), .Y(\CONFIG_reg_o_2_13_1_1[6] )
        );
    CFG4 #( .INIT(16'hC5CA) )  
        \xhdl1.GEN_BITS[0].APB_32.INTR_reg_9_0_0_m2[0]  (.A(gpin3_0), 
        .B(N_175), .C(\CONFIG_reg[0][6] ), .D(\CONFIG_reg[0][5] ), .Y(
        N_5941));
    CFG2 #( .INIT(4'h8) )  
        \xhdl1.GEN_BITS[4].REG_GEN.CONFIG_reg[4]_RNICC9B[1]  (.A(
        \gpin3[4] ), .B(\CONFIG_reg[4][1] ), .Y(r_m1_e_1_0));
    CFG2 #( .INIT(4'h8) )  
        \xhdl1.GEN_BITS[5].REG_GPOUT.un54_GPIO_OUT_i  (.A(GPOUT_reg_5), 
        .B(\CONFIG_reg[5][0] ), .Y(GPIO_OUT_net_2[5]));
    CFG4 #( .INIT(16'h2000) )  
        \xhdl1.GEN_BITS[5].REG_GEN.CONFIG_reg[5]2_0_a4_0_a2  (.A(
        CoreAPB3_0_APBmslave2_PADDR[2]), .B(
        CoreAPB3_0_APBmslave2_PADDR[3]), .C(N_603), .D(N_604), .Y(
        \CONFIG_reg[5]2 ));
    CFG4 #( .INIT(16'hAC0F) )  
        \xhdl1.GEN_BITS[29].REG_GEN.CONFIG_reg[29]_RNIEMI52[2]  (.A(
        \CONFIG_reg[13][2] ), .B(\CONFIG_reg[29][2] ), .C(
        \CONFIG_reg_o_2_21_1_1[2] ), .D(CoreAPB3_0_APBmslave2_PADDR[5])
        , .Y(N_4821));
    CFG4 #( .INIT(16'h0A33) )  
        \xhdl1.GEN_BITS[24].APB_32.INTR_reg_321_0[24]  (.A(INTR_reg_24)
        , .B(\INTR_reg_321_0_o2_1[24] ), .C(
        CoreAPB3_0_APBmslave2_PWDATA[24]), .D(edge_N_5_mux), .Y(
        \INTR_reg_321[24] ));
    CFG2 #( .INIT(4'hB) )  edge_both_2_sqmuxa_27_i (.A(edge_N_5_mux), 
        .B(\CONFIG_reg[28][3] ), .Y(N_163));
    SLE \xhdl1.GEN_BITS[7].REG_GEN.CONFIG_reg[7][3]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[3]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[7]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[7][3] ));
    SLE \xhdl1.GEN_BITS[2].REG_GEN.CONFIG_reg[2][1]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[1]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[2]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[2]_1 ));
    CFG4 #( .INIT(16'h0F35) )  
        \xhdl1.GEN_BITS[18].REG_GEN.CONFIG_reg[18]_RNIE0I61[3]  (.A(
        \CONFIG_reg[2][3] ), .B(\CONFIG_reg[18][3] ), .C(
        CoreAPB3_0_APBmslave2_PADDR[6]), .D(
        CoreAPB3_0_APBmslave2_PADDR[5]), .Y(\CONFIG_reg_o_2_10_1_1[3] )
        );
    SLE \xhdl1.GEN_BITS[6].APB_32.GPOUT_reg[6]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[6]), .CLK(FCCC_0_GL1), .EN(
        GPOUT_reg_0_sqmuxa), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        GPOUT_reg_6));
    VCC VCC (.Y(VCC_net_1));
    SLE \xhdl1.GEN_BITS[21].REG_GEN.CONFIG_reg[21][3]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[3]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[21]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[21][3] ));
    CFG4 #( .INIT(16'hF2F3) )  
        \xhdl1.GEN_BITS[31].APB_32.INTR_reg_412_0_o2_1_0[31]  (.A(
        \CONFIG_reg[31][6] ), .B(\edge_pos[31] ), .C(
        \INTR_reg_412_0_o2_0[31] ), .D(\CONFIG_reg[31][5] ), .Y(
        \INTR_reg_412_0_o2_1[31] ));
    SLE \xhdl1.GEN_BITS[20].REG_GEN.CONFIG_reg[20][1]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[1]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[20]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[20][1] ));
    SLE \xhdl1.GEN_BITS[29].REG_GEN.CONFIG_reg[29][3]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[3]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[29]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[29][3] ));
    SLE \xhdl1.GEN_BITS[7].REG_GEN.CONFIG_reg[7][7]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[7]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[7]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[7][7] ));
    CFG4 #( .INIT(16'hF2F3) )  
        \xhdl1.GEN_BITS[18].APB_32.INTR_reg_243_0_o2_1_0[18]  (.A(
        \CONFIG_reg[18][6] ), .B(\edge_neg[18] ), .C(
        \INTR_reg_243_0_o2_0[18] ), .D(\CONFIG_reg[18][5] ), .Y(
        \INTR_reg_243_0_o2_1[18] ));
    SLE \xhdl1.GEN_BITS[3].REG_GEN.CONFIG_reg[3][5]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[5]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[3]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[3][5] ));
    CFG2 #( .INIT(4'hB) )  edge_both_2_sqmuxa_31_i (.A(edge_N_5_mux), 
        .B(\CONFIG_reg[24][3] ), .Y(N_155));
    CFG2 #( .INIT(4'hB) )  edge_both_2_sqmuxa_25_i (.A(edge_N_5_mux), 
        .B(\CONFIG_reg[30][3] ), .Y(edge_neg_2_sqmuxa_6_i_1));
    CFG4 #( .INIT(16'h0F35) )  
        \xhdl1.GEN_BITS[4].REG_GEN.CONFIG_reg[4]_RNI67V31[4]  (.A(
        \CONFIG_reg[4][4] ), .B(\CONFIG_reg[20][4] ), .C(
        CoreAPB3_0_APBmslave2_PADDR[6]), .D(
        CoreAPB3_0_APBmslave2_PADDR[5]), .Y(\CONFIG_reg_o_2_6_1[4] ));
    CFG2 #( .INIT(4'hB) )  edge_both_2_sqmuxa_21_i (.A(edge_N_5_mux), 
        .B(\CONFIG_reg[7][3] ), .Y(edge_pos_2_sqmuxa_1_i_1));
    CFG4 #( .INIT(16'hF2F3) )  
        \xhdl1.GEN_BITS[20].APB_32.INTR_reg_269_0_o2_1_0[20]  (.A(
        \CONFIG_reg[20][6] ), .B(\edge_neg[20] ), .C(
        \INTR_reg_269_0_o2_0[20] ), .D(\CONFIG_reg[20][5] ), .Y(
        \INTR_reg_269_0_o2_1[20] ));
    CFG4 #( .INIT(16'h0F35) )  
        \xhdl1.GEN_BITS[16].REG_GEN.CONFIG_reg[16]_RNI00E11[0]  (.A(
        \CONFIG_reg[0][0] ), .B(\CONFIG_reg[16][0] ), .C(
        CoreAPB3_0_APBmslave2_PADDR[6]), .D(
        CoreAPB3_0_APBmslave2_PADDR[5]), .Y(\CONFIG_reg_o_2_3_1[0] ));
    CFG4 #( .INIT(16'h4000) )  
        \xhdl1.GEN_BITS[0].REG_GEN.CONFIG_reg[0]2_0_a4_0_a2_1  (.A(
        N_243), .B(wen_0), .C(GEN_m3_e_1), .D(iPSELS_2[5]), .Y(N_678));
    SLE \xhdl1.GEN_BITS[30].REG_GEN.CONFIG_reg[30][5]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[5]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[30]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[30][5] ));
    CFG4 #( .INIT(16'h0A33) )  
        \xhdl1.GEN_BITS[13].APB_32.INTR_reg_178_0[13]  (.A(INTR_reg_13)
        , .B(\INTR_reg_178_0_o2_1[13] ), .C(
        CoreAPB3_0_APBmslave2_PWDATA[13]), .D(edge_N_5_mux), .Y(
        \INTR_reg_178[13] ));
    CFG4 #( .INIT(16'hA9FF) )  
        \xhdl1.GEN_BITS[23].APB_32.INTR_reg_308_0_o2_0_0[23]  (.A(
        \CONFIG_reg[23][7] ), .B(\CONFIG_reg[23][6] ), .C(
        \CONFIG_reg[23][5] ), .D(\CONFIG_reg[23][3] ), .Y(
        \INTR_reg_308_0_o2_0[23] ));
    CFG4 #( .INIT(16'h0A33) )  
        \xhdl1.GEN_BITS[8].APB_32.INTR_reg_113_0[8]  (.A(INTR_reg_8), 
        .B(\INTR_reg_113_0_o2_1[8] ), .C(
        CoreAPB3_0_APBmslave2_PWDATA[8]), .D(edge_N_5_mux), .Y(
        \INTR_reg_113[8] ));
    SLE \xhdl1.GEN_BITS[10].APB_32.edge_both[10]  (.D(
        \edge_neg_149[10] ), .CLK(FCCC_0_GL1), .EN(N_184), .ALn(
        MSS_RESET_N_F2M_c), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\edge_pos[10] ));
    CFG4 #( .INIT(16'hA9FF) )  
        \xhdl1.GEN_BITS[29].APB_32.INTR_reg_386_0_o2_0_0[29]  (.A(
        \CONFIG_reg[29][7] ), .B(\CONFIG_reg[29][6] ), .C(
        \CONFIG_reg[29][5] ), .D(\CONFIG_reg[29][3] ), .Y(
        \INTR_reg_386_0_o2_0[29] ));
    CFG4 #( .INIT(16'h0F35) )  
        \xhdl1.GEN_BITS[22].REG_GEN.CONFIG_reg[22]_RNIAT291[2]  (.A(
        \CONFIG_reg[6][2] ), .B(\CONFIG_reg[22][2] ), .C(
        CoreAPB3_0_APBmslave2_PADDR[6]), .D(
        CoreAPB3_0_APBmslave2_PADDR[5]), .Y(\CONFIG_reg_o_2_13_1_1[2] )
        );
    SLE \xhdl1.GEN_BITS[20].REG_GEN.CONFIG_reg[20][5]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[5]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[20]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[20][5] ));
    SLE \xhdl1.GEN_BITS[15].REG_GEN.CONFIG_reg[15][7]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[7]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[15]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[15][7] ));
    SLE \xhdl1.GEN_BITS[3].APB_32.edge_both[3]  (.D(
        \edge_both_51_iv_i_0[3] ), .CLK(FCCC_0_GL1), .EN(
        edge_both_2_sqmuxa_12_i_1), .ALn(MSS_RESET_N_F2M_c), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\edge_both[3] ));
    CFG4 #( .INIT(16'hAA08) )  
        \xhdl1.GEN_BITS[6].APB_32.edge_pos_93_iv_i_0_0[6]  (.A(
        \CONFIG_reg[6][3] ), .B(\edge_pos[6] ), .C(
        CoreAPB3_0_APBmslave2_PWDATA[6]), .D(N_689), .Y(N_99));
    SLE \xhdl1.GEN_BITS[30].APB_32.INTR_reg[30]  (.D(
        \INTR_reg_399[30] ), .CLK(FCCC_0_GL1), .EN(VCC_net_1), .ALn(
        MSS_RESET_N_F2M_c), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(INTR_reg_30));
    CFG2 #( .INIT(4'hB) )  edge_both_2_sqmuxa_5_i (.A(edge_N_5_mux), 
        .B(\CONFIG_reg[14][3] ), .Y(edge_pos_2_sqmuxa_8_i_1));
    SLE \xhdl1.GEN_BITS[7].APB_32.INTR_reg[7]  (.D(\INTR_reg_100[7] ), 
        .CLK(FCCC_0_GL1), .EN(VCC_net_1), .ALn(MSS_RESET_N_F2M_c), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(INTR_reg_7));
    CFG4 #( .INIT(16'h2000) )  
        \xhdl1.GEN_BITS[2].REG_GEN.CONFIG_reg[2]2_0_a4_0_a2  (.A(
        CoreAPB3_0_APBmslave2_PADDR[3]), .B(
        CoreAPB3_0_APBmslave2_PADDR[2]), .C(N_604), .D(N_606), .Y(
        \CONFIG_reg[2]2 ));
    CFG4 #( .INIT(16'hAA08) )  
        \xhdl1.GEN_BITS[1].APB_32.edge_both_23_iv_i_0[1]  (.A(
        \CONFIG_reg[1][3] ), .B(\edge_both[1] ), .C(
        CoreAPB3_0_APBmslave2_PWDATA[1]), .D(N_142_i), .Y(N_95));
    CFG2 #( .INIT(4'h8) )  
        \xhdl1.GEN_BITS[12].REG_GEN.CONFIG_reg[12]2_0_a4_0_a2  (.A(
        N_678), .B(N_605), .Y(\CONFIG_reg[12]2 ));
    SLE \xhdl1.GEN_BITS[1].REG_GEN.CONFIG_reg[1][1]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[1]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[1]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[1]_1 ));
    SLE \xhdl1.GEN_BITS[6].REG_GEN.CONFIG_reg[6][5]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[5]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[6]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[6][5] ));
    SLE \xhdl1.GEN_BITS[16].APB_32.GPOUT_reg[16]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[16]), .CLK(FCCC_0_GL1), .EN(
        GPOUT_reg_0_sqmuxa), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        GPOUT_reg_16));
    CFG4 #( .INIT(16'h0ACC) )  
        \xhdl1.GEN_BITS[6].APB_32.INTR_reg_87_0_0[6]  (.A(INTR_reg_6), 
        .B(\INTR_reg_87_0_0_0_tz[6] ), .C(
        CoreAPB3_0_APBmslave2_PWDATA[6]), .D(edge_N_5_mux), .Y(
        \INTR_reg_87[6] ));
    SLE \xhdl1.GEN_BITS[4].gpin3[4]  (.D(\gpin2[4] ), .CLK(FCCC_0_GL1), 
        .EN(VCC_net_1), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(\gpin3[4] ));
    CFG4 #( .INIT(16'hC5CA) )  
        \xhdl1.GEN_BITS[6].APB_32.INTR_reg_87_0_0_m2[6]  (.A(gpin3_6), 
        .B(N_5938), .C(\CONFIG_reg[6][6] ), .D(\CONFIG_reg[6][5] ), .Y(
        N_5939));
    CFG4 #( .INIT(16'hF2F3) )  
        \xhdl1.GEN_BITS[7].APB_32.INTR_reg_100_0_o2_1_0[7]  (.A(
        \CONFIG_reg[7][6] ), .B(\edge_pos[7] ), .C(
        \INTR_reg_100_0_o2_0[7] ), .D(\CONFIG_reg[7][5] ), .Y(
        \INTR_reg_100_0_o2_1[7] ));
    CFG3 #( .INIT(8'hB8) )  
        \xhdl1.GEN_BITS[2].APB_32.INTR_reg_35_0_m2_0[2]  (.A(
        \edge_neg[2] ), .B(\CONFIG_reg[2][5] ), .C(\edge_pos[2] ), .Y(
        N_173));
    CFG4 #( .INIT(16'hF2F3) )  
        \xhdl1.GEN_BITS[29].APB_32.INTR_reg_386_0_o2_1_0[29]  (.A(
        \CONFIG_reg[29][6] ), .B(\edge_pos[29] ), .C(
        \INTR_reg_386_0_o2_0[29] ), .D(\CONFIG_reg[29][5] ), .Y(
        \INTR_reg_386_0_o2_1[29] ));
    CFG3 #( .INIT(8'h20) )  
        \xhdl1.GEN_BITS[10].APB_32.edge_both_RNO[10]  (.A(
        \CONFIG_reg[10][3] ), .B(CoreAPB3_0_APBmslave2_PWDATA[10]), .C(
        \edge_pos[10] ), .Y(\edge_neg_149[10] ));
    SLE \xhdl1.GEN_BITS[23].APB_32.edge_both[23]  (.D(N_96_i_0), .CLK(
        FCCC_0_GL1), .EN(edge_pos_2_sqmuxa_26_i_1), .ALn(
        MSS_RESET_N_F2M_c), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\edge_neg[23] ));
    CFG4 #( .INIT(16'hF2F3) )  
        \xhdl1.GEN_BITS[19].APB_32.INTR_reg_256_0_o2_1_0[19]  (.A(
        \CONFIG_reg[19][6] ), .B(\edge_neg[19] ), .C(
        \INTR_reg_256_0_o2_0[19] ), .D(\CONFIG_reg[19][5] ), .Y(
        \INTR_reg_256_0_o2_1[19] ));
    SLE \xhdl1.GEN_BITS[25].REG_GEN.CONFIG_reg[25][3]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[3]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[25]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[25][3] ));
    SLE \xhdl1.GEN_BITS[15].REG_GEN.CONFIG_reg[15][4]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[4]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[15]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[15][4] ));
    CFG3 #( .INIT(8'hFB) )  edge_pos_2_sqmuxa_5_i_0 (.A(edge_N_5_mux), 
        .B(\CONFIG_reg[1][3] ), .C(N_400), .Y(N_66));
    CFG4 #( .INIT(16'hA9FF) )  
        \xhdl1.GEN_BITS[9].APB_32.INTR_reg_126_0_o2_0_0[9]  (.A(
        \CONFIG_reg[9][7] ), .B(\CONFIG_reg[9][6] ), .C(
        \CONFIG_reg[9][5] ), .D(\CONFIG_reg[9][3] ), .Y(
        \INTR_reg_126_0_o2_0[9] ));
    SLE \xhdl1.GEN_BITS[3].APB_32.edge_neg[3]  (.D(
        \edge_neg_51_iv_i_1[3] ), .CLK(FCCC_0_GL1), .EN(N_81), .ALn(
        MSS_RESET_N_F2M_c), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\edge_neg[3] ));
    CFG4 #( .INIT(16'h8000) )  
        \xhdl1.GEN_BITS[11].REG_GEN.CONFIG_reg[11]2_0_a4_0_a2  (.A(
        CoreAPB3_0_APBmslave2_PADDR[3]), .B(
        CoreAPB3_0_APBmslave2_PADDR[2]), .C(N_604), .D(N_610), .Y(
        \CONFIG_reg[11]2 ));
    SLE \xhdl1.GEN_BITS[13].REG_GEN.CONFIG_reg[13][6]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[6]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[13]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[13][6] ));
    SLE \xhdl1.GEN_BITS[11].APB_32.INTR_reg[11]  (.D(
        \INTR_reg_152[11] ), .CLK(FCCC_0_GL1), .EN(VCC_net_1), .ALn(
        MSS_RESET_N_F2M_c), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(INTR_reg_11));
    CFG4 #( .INIT(16'h0F35) )  
        \xhdl1.GEN_BITS[21].REG_GEN.CONFIG_reg[21]_RNI4UG61[1]  (.A(
        \CONFIG_reg[5]_1 ), .B(\CONFIG_reg[21][1] ), .C(
        CoreAPB3_0_APBmslave2_PADDR[6]), .D(
        CoreAPB3_0_APBmslave2_PADDR[5]), .Y(\CONFIG_reg_o_2_21_1_1[1] )
        );
    CFG3 #( .INIT(8'hFB) )  edge_pos_2_sqmuxa_3_i_0 (.A(edge_N_5_mux), 
        .B(\CONFIG_reg[5][3] ), .C(N_406), .Y(N_70));
    CFG4 #( .INIT(16'hAC0F) )  
        \xhdl1.GEN_BITS[15].REG_GEN.CONFIG_reg[15]_RNIKVN32[4]  (.A(
        \CONFIG_reg[15][4] ), .B(\CONFIG_reg[31][4] ), .C(
        \CONFIG_reg_o_2_28_1_1[4] ), .D(CoreAPB3_0_APBmslave2_PADDR[5])
        , .Y(N_4879));
    CFG4 #( .INIT(16'h0A33) )  
        \xhdl1.GEN_BITS[29].APB_32.INTR_reg_386_0[29]  (.A(INTR_reg_29)
        , .B(\INTR_reg_386_0_o2_1[29] ), .C(
        CoreAPB3_0_APBmslave2_PWDATA[29]), .D(edge_N_5_mux), .Y(
        \INTR_reg_386[29] ));
    SLE \xhdl1.GEN_BITS[10].REG_GEN.CONFIG_reg[10][7]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[7]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[10]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[10][7] ));
    CFG2 #( .INIT(4'h4) )  PRDATA_m1_e (.A(N_245), .B(PRDATA_m1_e_1), 
        .Y(N_452));
    CFG4 #( .INIT(16'hA9FF) )  
        \xhdl1.GEN_BITS[26].APB_32.INTR_reg_347_0_o2_0_0[26]  (.A(
        \CONFIG_reg[26][7] ), .B(\CONFIG_reg[26][6] ), .C(
        \CONFIG_reg[26][5] ), .D(\CONFIG_reg[26][3] ), .Y(
        \INTR_reg_347_0_o2_0[26] ));
    SLE \xhdl1.GEN_BITS[14].REG_GEN.CONFIG_reg[14][7]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[7]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[14]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[14][7] ));
    SLE \xhdl1.GEN_BITS[27].REG_GEN.CONFIG_reg[27][6]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[6]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[27]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[27][6] ));
    CFG4 #( .INIT(16'hFFEF) )  \RDATA_32.un12_PRDATA_o_0_o2  (.A(
        CoreAPB3_0_APBmslave2_PADDR[0]), .B(N_243), .C(
        CoreAPB3_0_APBmslave2_PADDR[7]), .D(
        CoreAPB3_0_APBmslave2_PADDR[1]), .Y(N_245));
    CFG2 #( .INIT(4'hB) )  edge_both_2_sqmuxa_10_i (.A(edge_N_5_mux), 
        .B(\CONFIG_reg[18][3] ), .Y(N_192));
    CFG4 #( .INIT(16'hA9FF) )  
        \xhdl1.GEN_BITS[18].APB_32.INTR_reg_243_0_o2_0_0[18]  (.A(
        \CONFIG_reg[18][7] ), .B(\CONFIG_reg[18][6] ), .C(
        \CONFIG_reg[18][5] ), .D(\CONFIG_reg[18][3] ), .Y(
        \INTR_reg_243_0_o2_0[18] ));
    CFG3 #( .INIT(8'h35) )  
        \xhdl1.GEN_BITS[3].APB_32.GPOUT_reg_RNI20L91[3]  (.A(
        \INTR_reg[3] ), .B(\GPOUT_reg[3] ), .C(
        CoreAPB3_0_APBmslave2_PADDR[5]), .Y(PRDATA_N_3_0));
    SLE \xhdl1.GEN_BITS[30].REG_GEN.CONFIG_reg[30][3]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[3]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[30]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[30][3] ));
    CFG2 #( .INIT(4'hB) )  edge_both_2_sqmuxa_1_i (.A(edge_N_5_mux), 
        .B(\CONFIG_reg[17][3] ), .Y(edge_pos_2_sqmuxa_30_i_1));
    CFG2 #( .INIT(4'h6) )  edge_both_2_sqmuxa_15_i_x2 (.A(\gpin2[0] ), 
        .B(gpin3_0), .Y(N_141_i));
    CFG4 #( .INIT(16'h0F35) )  
        \xhdl1.GEN_BITS[19].REG_GEN.CONFIG_reg[19]_RNIKV391[4]  (.A(
        \CONFIG_reg[3][4] ), .B(\CONFIG_reg[19][4] ), .C(
        CoreAPB3_0_APBmslave2_PADDR[6]), .D(
        CoreAPB3_0_APBmslave2_PADDR[5]), .Y(\CONFIG_reg_o_2_25_1_1[4] )
        );
    CFG4 #( .INIT(16'hAC0F) )  
        \xhdl1.GEN_BITS[24].REG_GEN.CONFIG_reg[24]_RNIM8R22[5]  (.A(
        \CONFIG_reg[8][5] ), .B(\CONFIG_reg[24][5] ), .C(
        \CONFIG_reg_o_2_3_1_1[5] ), .D(CoreAPB3_0_APBmslave2_PADDR[5]), 
        .Y(N_4680));
    SLE \xhdl1.GEN_BITS[22].APB_32.edge_both[22]  (.D(
        \edge_neg_317[22] ), .CLK(FCCC_0_GL1), .EN(N_200), .ALn(
        MSS_RESET_N_F2M_c), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\edge_neg[22] ));
    CFG4 #( .INIT(16'h0F35) )  
        \xhdl1.GEN_BITS[7].REG_GEN.CONFIG_reg[7]_RNIGSKB1[3]  (.A(
        \CONFIG_reg[7][3] ), .B(\CONFIG_reg[23][3] ), .C(
        CoreAPB3_0_APBmslave2_PADDR[6]), .D(
        CoreAPB3_0_APBmslave2_PADDR[5]), .Y(\CONFIG_reg_o_2_28_1_1[3] )
        );
    CFG4 #( .INIT(16'h0F35) )  
        \xhdl1.GEN_BITS[18].REG_GEN.CONFIG_reg[18]_RNI8QH61[0]  (.A(
        \CONFIG_reg[2][0] ), .B(\CONFIG_reg[18][0] ), .C(
        CoreAPB3_0_APBmslave2_PADDR[6]), .D(
        CoreAPB3_0_APBmslave2_PADDR[5]), .Y(\CONFIG_reg_o_2_10_1_1[0] )
        );
    CFG3 #( .INIT(8'h20) )  
        \xhdl1.GEN_BITS[28].APB_32.edge_both_RNO[28]  (.A(
        \CONFIG_reg[28][3] ), .B(CoreAPB3_0_APBmslave2_PWDATA[28]), .C(
        \edge_pos[28] ), .Y(N_87_i_0));
    CFG4 #( .INIT(16'h0A33) )  
        \xhdl1.GEN_BITS[20].APB_32.INTR_reg_269_0[20]  (.A(INTR_reg_20)
        , .B(\INTR_reg_269_0_o2_1[20] ), .C(
        CoreAPB3_0_APBmslave2_PWDATA[20]), .D(edge_N_5_mux), .Y(
        \INTR_reg_269[20] ));
    CFG3 #( .INIT(8'h20) )  
        \xhdl1.GEN_BITS[12].APB_32.edge_both_RNO[12]  (.A(
        \CONFIG_reg[12][3] ), .B(CoreAPB3_0_APBmslave2_PWDATA[12]), .C(
        \edge_neg[12] ), .Y(\edge_neg_177[12] ));
    CFG2 #( .INIT(4'hB) )  edge_both_2_sqmuxa_17_i (.A(edge_N_5_mux), 
        .B(\CONFIG_reg[11][3] ), .Y(N_186));
    CFG4 #( .INIT(16'hA9FF) )  
        \xhdl1.GEN_BITS[12].APB_32.INTR_reg_165_0_o2_0_0[12]  (.A(
        \CONFIG_reg[12][7] ), .B(\CONFIG_reg[12][6] ), .C(
        \CONFIG_reg[12][5] ), .D(\CONFIG_reg[12][3] ), .Y(
        \INTR_reg_165_0_o2_0[12] ));
    SLE \xhdl1.GEN_BITS[1].APB_32.GPOUT_reg[1]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[1]), .CLK(FCCC_0_GL1), .EN(
        GPOUT_reg_0_sqmuxa), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        GPOUT_reg_1));
    CFG4 #( .INIT(16'hF2F3) )  
        \xhdl1.GEN_BITS[13].APB_32.INTR_reg_178_0_o2_1_0[13]  (.A(
        \CONFIG_reg[13][6] ), .B(\edge_neg[13] ), .C(
        \INTR_reg_178_0_o2_0[13] ), .D(\CONFIG_reg[13][5] ), .Y(
        \INTR_reg_178_0_o2_1[13] ));
    SLE \xhdl1.GEN_BITS[21].REG_GEN.CONFIG_reg[21][7]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[7]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[21]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[21][7] ));
    CFG3 #( .INIT(8'h20) )  
        \xhdl1.GEN_BITS[9].APB_32.edge_both_RNO[9]  (.A(
        \CONFIG_reg[9][3] ), .B(CoreAPB3_0_APBmslave2_PWDATA[9]), .C(
        \edge_neg[9] ), .Y(\edge_neg_135[9] ));
    CFG2 #( .INIT(4'h8) )  
        \xhdl1.GEN_BITS[2].REG_GPOUT.un24_GPIO_OUT_i  (.A(GPOUT_reg_2), 
        .B(\CONFIG_reg[2][0] ), .Y(GPIO_OUT_net_2[2]));
    CFG4 #( .INIT(16'h0ACC) )  
        \xhdl1.GEN_BITS[2].APB_32.INTR_reg_35_0_0[2]  (.A(INTR_reg_2), 
        .B(\INTR_reg_35_0_0_0_tz[2] ), .C(
        CoreAPB3_0_APBmslave2_PWDATA[2]), .D(edge_N_5_mux), .Y(
        \INTR_reg_35[2] ));
    SLE \xhdl1.GEN_BITS[23].REG_GEN.CONFIG_reg[23][7]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[7]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[23]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[23][7] ));
    SLE \xhdl1.GEN_BITS[12].APB_32.GPOUT_reg[12]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[12]), .CLK(FCCC_0_GL1), .EN(
        GPOUT_reg_0_sqmuxa), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        GPOUT_reg_12));
    CFG2 #( .INIT(4'hE) )  
        \xhdl1.GEN_BITS[0].APB_32.un5_PRDATA_o_0_a2_0_o2_s  (.A(
        CoreAPB3_0_APBmslave2_PADDR[5]), .B(
        CoreAPB3_0_APBmslave2_PADDR[4]), .Y(un5_PRDATA_o_0_a2_0_o2_out)
        );
    SLE \xhdl1.GEN_BITS[19].REG_GEN.CONFIG_reg[19][0]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[0]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[19]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[19][0] ));
    SLE \xhdl1.GEN_BITS[20].REG_GEN.CONFIG_reg[20][3]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[3]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[20]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[20][3] ));
    CFG4 #( .INIT(16'h0A33) )  
        \xhdl1.GEN_BITS[7].APB_32.INTR_reg_100_0[7]  (.A(INTR_reg_7), 
        .B(\INTR_reg_100_0_o2_1[7] ), .C(
        CoreAPB3_0_APBmslave2_PWDATA[7]), .D(edge_N_5_mux), .Y(
        \INTR_reg_100[7] ));
    SLE \xhdl1.GEN_BITS[25].REG_GEN.CONFIG_reg[25][4]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[4]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[25]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[25][4] ));
    SLE \xhdl1.GEN_BITS[12].REG_GEN.CONFIG_reg[12][4]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[4]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[12]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[12][4] ));
    CFG3 #( .INIT(8'h04) )  
        \xhdl1.GEN_BITS[4].APB_32.INTR_reg_61_0_0_0_tz_1[4]  (.A(
        \CONFIG_reg[4][5] ), .B(\edge_both[4] ), .C(\CONFIG_reg[4][6] )
        , .Y(\INTR_reg_61_0_0_0_tz_1[4] ));
    SLE \xhdl1.GEN_BITS[4].APB_32.edge_both[4]  (.D(N_91), .CLK(
        FCCC_0_GL1), .EN(N_84), .ALn(MSS_RESET_N_F2M_c), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\edge_both[4] ));
    SLE \xhdl1.GEN_BITS[9].REG_GEN.CONFIG_reg[9][3]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[3]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[9]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[9][3] ));
    SLE \xhdl1.GEN_BITS[29].REG_GEN.CONFIG_reg[29][7]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[7]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[29]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[29][7] ));
    CFG4 #( .INIT(16'hAC0F) )  
        \xhdl1.GEN_BITS[26].REG_GEN.CONFIG_reg[26]_RNIG2GS1[4]  (.A(
        \CONFIG_reg[10][4] ), .B(\CONFIG_reg[26][4] ), .C(
        \CONFIG_reg_o_2_10_1_1[4] ), .D(CoreAPB3_0_APBmslave2_PADDR[5])
        , .Y(N_4735));
    SLE \xhdl1.GEN_BITS[17].REG_GEN.CONFIG_reg[17][1]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[1]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[17]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[17][1] ));
    CFG4 #( .INIT(16'hF2F3) )  
        \xhdl1.GEN_BITS[25].APB_32.INTR_reg_334_0_o2_1_0[25]  (.A(
        \CONFIG_reg[25][6] ), .B(\edge_neg[25] ), .C(
        \INTR_reg_334_0_o2_0[25] ), .D(\CONFIG_reg[25][5] ), .Y(
        \INTR_reg_334_0_o2_1[25] ));
    CFG4 #( .INIT(16'hAA08) )  
        \xhdl1.GEN_BITS[3].APB_32.edge_neg_51_iv_i_0[3]  (.A(
        \CONFIG_reg[3][3] ), .B(\edge_neg[3] ), .C(
        CoreAPB3_0_APBmslave2_PWDATA[3]), .D(N_686), .Y(
        \edge_neg_51_iv_i_1[3] ));
    CFG4 #( .INIT(16'h0F35) )  
        \xhdl1.GEN_BITS[19].REG_GEN.CONFIG_reg[19]_RNIEP391[1]  (.A(
        \CONFIG_reg[3]_1 ), .B(\CONFIG_reg[19][1] ), .C(
        CoreAPB3_0_APBmslave2_PADDR[6]), .D(
        CoreAPB3_0_APBmslave2_PADDR[5]), .Y(\CONFIG_reg_o_2_25_1_1[1] )
        );
    CFG2 #( .INIT(4'hB) )  edge_both_2_sqmuxa_13_i (.A(edge_N_5_mux), 
        .B(\CONFIG_reg[29][3] ), .Y(N_190));
    CFG4 #( .INIT(16'hA9FF) )  
        \xhdl1.GEN_BITS[17].APB_32.INTR_reg_230_0_o2_0_0[17]  (.A(
        \CONFIG_reg[17][7] ), .B(\CONFIG_reg[17][6] ), .C(
        \CONFIG_reg[17][5] ), .D(\CONFIG_reg[17][3] ), .Y(
        \INTR_reg_230_0_o2_0[17] ));
    SLE \xhdl1.GEN_BITS[8].REG_GEN.CONFIG_reg[8][3]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[3]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[8]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[8][3] ));
    CFG2 #( .INIT(4'hB) )  edge_both_2_sqmuxa_2_i (.A(edge_N_5_mux), 
        .B(\CONFIG_reg[13][3] ), .Y(edge_pos_2_sqmuxa_9_i_1));
    SLE \xhdl1.GEN_BITS[7].APB_32.edge_both[7]  (.D(N_83_i_0), .CLK(
        FCCC_0_GL1), .EN(edge_pos_2_sqmuxa_1_i_1), .ALn(
        MSS_RESET_N_F2M_c), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\edge_pos[7] ));
    CFG4 #( .INIT(16'h0ACC) )  
        \xhdl1.GEN_BITS[5].APB_32.INTR_reg_74_0_0[5]  (.A(INTR_reg_5), 
        .B(\INTR_reg_74_0_0_0_tz[5] ), .C(
        CoreAPB3_0_APBmslave2_PWDATA[5]), .D(edge_N_5_mux), .Y(
        \INTR_reg_74[5] ));
    CFG4 #( .INIT(16'hC480) )  
        \xhdl1.GEN_BITS[2].APB_32.INTR_reg_35_0_0_0_tz[2]  (.A(
        \CONFIG_reg[2][7] ), .B(\CONFIG_reg[2][3] ), .C(
        \INTR_reg_35_0_0_0_tz_1[2] ), .D(N_178), .Y(
        \INTR_reg_35_0_0_0_tz[2] ));
    CFG4 #( .INIT(16'hA9FF) )  
        \xhdl1.GEN_BITS[7].APB_32.INTR_reg_100_0_o2_0_0[7]  (.A(
        \CONFIG_reg[7][7] ), .B(\CONFIG_reg[7][6] ), .C(
        \CONFIG_reg[7][5] ), .D(\CONFIG_reg[7][3] ), .Y(
        \INTR_reg_100_0_o2_0[7] ));
    SLE \xhdl1.GEN_BITS[2].REG_GEN.CONFIG_reg[2][2]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[2]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[2]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[2][2] ));
    SLE \xhdl1.GEN_BITS[9].REG_GEN.CONFIG_reg[9][7]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[7]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[9]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[9][7] ));
    SLE \xhdl1.GEN_BITS[0].gpin3[0]  (.D(\gpin2[0] ), .CLK(FCCC_0_GL1), 
        .EN(VCC_net_1), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(gpin3_0));
    CFG4 #( .INIT(16'h0F35) )  
        \xhdl1.GEN_BITS[20].REG_GEN.CONFIG_reg[20]_RNI01V31[1]  (.A(
        \CONFIG_reg[4][1] ), .B(\CONFIG_reg[20][1] ), .C(
        CoreAPB3_0_APBmslave2_PADDR[6]), .D(
        CoreAPB3_0_APBmslave2_PADDR[5]), .Y(\CONFIG_reg_o_2_6_1_1[1] ));
    SLE \xhdl1.GEN_BITS[8].APB_32.GPOUT_reg[8]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[8]), .CLK(FCCC_0_GL1), .EN(
        GPOUT_reg_0_sqmuxa), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        GPOUT_reg_8));
    SLE \xhdl1.GEN_BITS[19].REG_GEN.CONFIG_reg[19][5]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[5]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[19]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[19][5] ));
    CFG4 #( .INIT(16'h8000) )  
        \xhdl1.GEN_BITS[23].REG_GEN.CONFIG_reg[23]2_0_a4_0_a2  (.A(
        CoreAPB3_0_APBmslave2_PADDR[3]), .B(
        CoreAPB3_0_APBmslave2_PADDR[2]), .C(N_598), .D(N_603), .Y(
        \CONFIG_reg[23]2 ));
    CFG4 #( .INIT(16'h0F35) )  
        \xhdl1.GEN_BITS[17].REG_GEN.CONFIG_reg[17]_RNIE70K1[5]  (.A(
        \CONFIG_reg[1][5] ), .B(\CONFIG_reg[17][5] ), .C(
        CoreAPB3_0_APBmslave2_PADDR[6]), .D(
        CoreAPB3_0_APBmslave2_PADDR[5]), .Y(\CONFIG_reg_o_2_18_1_1[5] )
        );
    SLE \xhdl1.GEN_BITS[15].REG_GEN.CONFIG_reg[15][2]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[2]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[15]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[15][2] ));
    CFG4 #( .INIT(16'h2000) )  
        \xhdl1.GEN_BITS[14].REG_GEN.CONFIG_reg[14]2_0_a4_0_a2  (.A(
        CoreAPB3_0_APBmslave2_PADDR[3]), .B(
        CoreAPB3_0_APBmslave2_PADDR[2]), .C(N_604), .D(N_605), .Y(
        \CONFIG_reg[14]2 ));
    SLE \xhdl1.GEN_BITS[30].APB_32.GPOUT_reg[30]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[30]), .CLK(FCCC_0_GL1), .EN(
        GPOUT_reg_0_sqmuxa), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        GPOUT_reg_30));
    SLE \xhdl1.GEN_BITS[0].REG_GEN.CONFIG_reg[0][4]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[4]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[0]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[0][4] ));
    SLE \xhdl1.GEN_BITS[8].REG_GEN.CONFIG_reg[8][7]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[7]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[8]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[8][7] ));
    CFG3 #( .INIT(8'h20) )  
        \xhdl1.GEN_BITS[17].APB_32.edge_both_RNO[17]  (.A(
        \CONFIG_reg[17][3] ), .B(CoreAPB3_0_APBmslave2_PWDATA[17]), .C(
        \edge_neg[17] ), .Y(\edge_neg_247[17] ));
    SLE \xhdl1.GEN_BITS[15].APB_32.edge_pos[15]  (.D(
        \edge_pos_219[15] ), .CLK(FCCC_0_GL1), .EN(
        edge_pos_2_sqmuxa_7_i_1), .ALn(MSS_RESET_N_F2M_c), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\edge_neg[15] ));
    SLE \xhdl1.GEN_BITS[21].APB_32.GPOUT_reg[21]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[21]), .CLK(FCCC_0_GL1), .EN(
        GPOUT_reg_0_sqmuxa), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        GPOUT_reg_21));
    CFG4 #( .INIT(16'h0F35) )  
        \xhdl1.GEN_BITS[19].REG_GEN.CONFIG_reg[19]_RNIQ5491[7]  (.A(
        \CONFIG_reg[3][7] ), .B(\CONFIG_reg[19][7] ), .C(
        CoreAPB3_0_APBmslave2_PADDR[6]), .D(
        CoreAPB3_0_APBmslave2_PADDR[5]), .Y(\CONFIG_reg_o_2_25_1_1[7] )
        );
    CFG4 #( .INIT(16'hAC0F) )  
        \xhdl1.GEN_BITS[14].REG_GEN.CONFIG_reg[14]_RNISJP82[0]  (.A(
        \CONFIG_reg[14][0] ), .B(\CONFIG_reg[30][0] ), .C(
        \CONFIG_reg_o_2_13_1_1[0] ), .D(CoreAPB3_0_APBmslave2_PADDR[5])
        , .Y(N_4755));
    CFG4 #( .INIT(16'h4000) )  
        \xhdl1.GEN_BITS[2].REG_GEN.CONFIG_reg[2]2_0_a4_0_a2_1  (.A(
        CoreAPB3_0_APBmslave2_PADDR[6]), .B(wen_0), .C(GEN_m3_e_1), .D(
        iPSELS_2[5]), .Y(N_604));
    CFG3 #( .INIT(8'hFB) )  edge_neg_2_sqmuxa_8_i_0 (.A(edge_N_5_mux), 
        .B(\CONFIG_reg[4][3] ), .C(N_397), .Y(N_58));
    SLE \xhdl1.GEN_BITS[25].REG_GEN.CONFIG_reg[25][5]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[5]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[25]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[25][5] ));
    CFG4 #( .INIT(16'h2000) )  
        \xhdl1.GEN_BITS[18].REG_GEN.CONFIG_reg[18]2_0_a4_0_a2  (.A(
        CoreAPB3_0_APBmslave2_PADDR[3]), .B(
        CoreAPB3_0_APBmslave2_PADDR[2]), .C(N_598), .D(N_606), .Y(
        \CONFIG_reg[18]2 ));
    SLE \xhdl1.GEN_BITS[16].REG_GEN.CONFIG_reg[16][6]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[6]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[16]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[16][6] ));
    SLE \xhdl1.GEN_BITS[15].REG_GEN.CONFIG_reg[15][5]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[5]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[15]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[15][5] ));
    SLE \xhdl1.GEN_BITS[17].APB_32.INTR_reg[17]  (.D(
        \INTR_reg_230[17] ), .CLK(FCCC_0_GL1), .EN(VCC_net_1), .ALn(
        MSS_RESET_N_F2M_c), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(INTR_reg_17));
    SLE \xhdl1.GEN_BITS[3].REG_GEN.CONFIG_reg[3][3]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[3]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[3]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[3][3] ));
    SLE \xhdl1.GEN_BITS[29].REG_GEN.CONFIG_reg[29][6]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[6]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[29]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[29][6] ));
    SLE \xhdl1.GEN_BITS[16].REG_GEN.CONFIG_reg[16][4]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[4]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[16]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[16][4] ));
    SLE \xhdl1.GEN_BITS[5].APB_32.edge_neg[5]  (.D(N_115), .CLK(
        FCCC_0_GL1), .EN(N_60), .ALn(MSS_RESET_N_F2M_c), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\edge_neg[5] ));
    SLE \xhdl1.GEN_BITS[21].APB_32.edge_both[21]  (.D(
        \edge_neg_303[21] ), .CLK(FCCC_0_GL1), .EN(N_198), .ALn(
        MSS_RESET_N_F2M_c), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\edge_neg[21] ));
    SLE \xhdl1.GEN_BITS[16].REG_GEN.CONFIG_reg[16][3]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[3]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[16]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[16][3] ));
    CFG3 #( .INIT(8'hFB) )  edge_both_2_sqmuxa_22_i_0_0 (.A(
        edge_N_5_mux), .B(\CONFIG_reg[6][3] ), .C(N_252_i), .Y(N_78));
    SLE \xhdl1.GEN_BITS[6].APB_32.edge_pos[6]  (.D(N_99), .CLK(
        FCCC_0_GL1), .EN(N_72), .ALn(MSS_RESET_N_F2M_c), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\edge_pos[6] ));
    SLE \xhdl1.GEN_BITS[3].REG_GEN.CONFIG_reg[3][7]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[7]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[3]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[3][7] ));
    CFG4 #( .INIT(16'hAC0F) )  
        \xhdl1.GEN_BITS[26].REG_GEN.CONFIG_reg[26]_RNIK6GS1[5]  (.A(
        \CONFIG_reg[10][5] ), .B(\CONFIG_reg[26][5] ), .C(
        \CONFIG_reg_o_2_10_1_1[5] ), .D(CoreAPB3_0_APBmslave2_PADDR[5])
        , .Y(N_4736));
    SLE \xhdl1.GEN_BITS[27].REG_GEN.CONFIG_reg[27][4]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[4]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[27]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[27][4] ));
    SLE \xhdl1.GEN_BITS[1].REG_GEN.CONFIG_reg[1][2]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[2]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[1]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[1][2] ));
    CFG4 #( .INIT(16'hAC0F) )  
        \xhdl1.GEN_BITS[9].REG_GEN.CONFIG_reg[9]_RNI6BV72[7]  (.A(
        \CONFIG_reg[9][7] ), .B(\CONFIG_reg[25][7] ), .C(
        \CONFIG_reg_o_2_18_1_1[7] ), .D(CoreAPB3_0_APBmslave2_PADDR[5])
        , .Y(N_4802));
    CFG4 #( .INIT(16'hAC0F) )  
        \xhdl1.GEN_BITS[29].REG_GEN.CONFIG_reg[29]_RNIIQI52[3]  (.A(
        \CONFIG_reg[13][3] ), .B(\CONFIG_reg[29][3] ), .C(
        \CONFIG_reg_o_2_21_1[3] ), .D(CoreAPB3_0_APBmslave2_PADDR[5]), 
        .Y(N_4822));
    SLE \xhdl1.GEN_BITS[0].REG_GEN.CONFIG_reg[0][6]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[6]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[0]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[0][6] ));
    CFG3 #( .INIT(8'h20) )  
        \xhdl1.GEN_BITS[25].APB_32.edge_both_RNO[25]  (.A(
        \CONFIG_reg[25][3] ), .B(CoreAPB3_0_APBmslave2_PWDATA[25]), .C(
        \edge_neg[25] ), .Y(N_5911_i_0));
    SLE \xhdl1.GEN_BITS[11].REG_GEN.CONFIG_reg[11][6]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[6]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[11]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[11][6] ));
    CFG4 #( .INIT(16'h2000) )  
        \xhdl1.GEN_BITS[22].REG_GEN.CONFIG_reg[22]2_0_a4_0_a2  (.A(
        CoreAPB3_0_APBmslave2_PADDR[3]), .B(
        CoreAPB3_0_APBmslave2_PADDR[2]), .C(N_598), .D(N_603), .Y(
        \CONFIG_reg[22]2 ));
    CFG3 #( .INIT(8'h20) )  
        \xhdl1.GEN_BITS[8].APB_32.edge_both_RNO[8]  (.A(
        \CONFIG_reg[8][3] ), .B(CoreAPB3_0_APBmslave2_PWDATA[8]), .C(
        \edge_pos[8] ), .Y(\edge_neg_121[8] ));
    CFG4 #( .INIT(16'hAA08) )  
        \xhdl1.GEN_BITS[0].APB_32.edge_both_9_iv_i_0[0]  (.A(
        \CONFIG_reg[0][3] ), .B(\edge_both[0] ), .C(
        CoreAPB3_0_APBmslave2_PWDATA[0]), .D(N_141_i), .Y(N_97));
    SLE \xhdl1.GEN_BITS[20].APB_32.INTR_reg[20]  (.D(
        \INTR_reg_269[20] ), .CLK(FCCC_0_GL1), .EN(VCC_net_1), .ALn(
        MSS_RESET_N_F2M_c), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(INTR_reg_20));
    SLE \xhdl1.GEN_BITS[14].REG_GEN.CONFIG_reg[14][6]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[6]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[14]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[14][6] ));
    CFG4 #( .INIT(16'h0F35) )  
        \xhdl1.GEN_BITS[19].REG_GEN.CONFIG_reg[19]_RNIIT391[3]  (.A(
        \CONFIG_reg[3][3] ), .B(\CONFIG_reg[19][3] ), .C(
        CoreAPB3_0_APBmslave2_PADDR[6]), .D(
        CoreAPB3_0_APBmslave2_PADDR[5]), .Y(\CONFIG_reg_o_2_25_1_1[3] )
        );
    CFG4 #( .INIT(16'h0F35) )  
        \xhdl1.GEN_BITS[7].REG_GEN.CONFIG_reg[7]_RNIEQKB1[2]  (.A(
        \CONFIG_reg[7][2] ), .B(\CONFIG_reg[23][2] ), .C(
        CoreAPB3_0_APBmslave2_PADDR[6]), .D(
        CoreAPB3_0_APBmslave2_PADDR[5]), .Y(\CONFIG_reg_o_2_28_1_1[2] )
        );
    SLE \xhdl1.GEN_BITS[6].REG_GEN.CONFIG_reg[6][3]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[3]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[6]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[6][3] ));
    CFG3 #( .INIT(8'hB8) )  \xhdl1.GEN_BITS[3].REG_INT.un34_intr_1  (
        .A(\edge_neg[3] ), .B(\CONFIG_reg[3][5] ), .C(\edge_pos[3] ), 
        .Y(N_4549));
    CFG2 #( .INIT(4'h4) )  
        \xhdl1.GEN_BITS[4].REG_GEN.CONFIG_reg[4]2_0_a4_0_a2_0  (.A(
        CoreAPB3_0_APBmslave2_PADDR[5]), .B(
        CoreAPB3_0_APBmslave2_PADDR[4]), .Y(N_603));
    SLE \xhdl1.GEN_BITS[4].APB_32.INTR_reg[4]  (.D(\INTR_reg_61[4] ), 
        .CLK(FCCC_0_GL1), .EN(VCC_net_1), .ALn(MSS_RESET_N_F2M_c), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(INTR_reg_4));
    CFG4 #( .INIT(16'hAA08) )  
        \xhdl1.GEN_BITS[3].APB_32.edge_pos_51_iv_i_0[3]  (.A(
        \CONFIG_reg[3][3] ), .B(\edge_pos[3] ), .C(
        CoreAPB3_0_APBmslave2_PWDATA[3]), .D(N_687), .Y(N_73));
    CFG4 #( .INIT(16'h0F35) )  
        \xhdl1.GEN_BITS[21].REG_GEN.CONFIG_reg[21]_RNI2SG61[0]  (.A(
        \CONFIG_reg[5][0] ), .B(\CONFIG_reg[21][0] ), .C(
        CoreAPB3_0_APBmslave2_PADDR[6]), .D(
        CoreAPB3_0_APBmslave2_PADDR[5]), .Y(\CONFIG_reg_o_2_21_1[0] ));
    SLE \xhdl1.GEN_BITS[21].REG_GEN.CONFIG_reg[21][2]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[2]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[21]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[21][2] ));
    CFG4 #( .INIT(16'hA9FF) )  
        \xhdl1.GEN_BITS[8].APB_32.INTR_reg_113_0_o2_0_0[8]  (.A(
        \CONFIG_reg[8][7] ), .B(\CONFIG_reg[8][6] ), .C(
        \CONFIG_reg[8][5] ), .D(\CONFIG_reg[8][3] ), .Y(
        \INTR_reg_113_0_o2_0[8] ));
    SLE \xhdl1.GEN_BITS[5].APB_32.INTR_reg[5]  (.D(\INTR_reg_74[5] ), 
        .CLK(FCCC_0_GL1), .EN(VCC_net_1), .ALn(MSS_RESET_N_F2M_c), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(INTR_reg_5));
    SLE \xhdl1.GEN_BITS[12].REG_GEN.CONFIG_reg[12][2]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[2]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[12]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[12][2] ));
    SLE \xhdl1.GEN_BITS[29].REG_GEN.CONFIG_reg[29][2]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[2]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[29]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[29][2] ));
    CFG4 #( .INIT(16'hF2F3) )  
        \xhdl1.GEN_BITS[30].APB_32.INTR_reg_399_0_o2_1_0[30]  (.A(
        \CONFIG_reg[30][6] ), .B(\edge_pos[30] ), .C(
        \INTR_reg_399_0_o2_0[30] ), .D(\CONFIG_reg[30][5] ), .Y(
        \INTR_reg_399_0_o2_1[30] ));
    CFG3 #( .INIT(8'h20) )  
        \xhdl1.GEN_BITS[30].APB_32.edge_both_RNO[30]  (.A(
        \CONFIG_reg[30][3] ), .B(CoreAPB3_0_APBmslave2_PWDATA[30]), .C(
        \edge_pos[30] ), .Y(\edge_neg_429[30] ));
    SLE \xhdl1.GEN_BITS[6].REG_GEN.CONFIG_reg[6][7]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[7]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[6]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[6][7] ));
    SLE \xhdl1.GEN_BITS[15].REG_GEN.CONFIG_reg[15][0]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[0]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[15]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[15][0] ));
    CFG4 #( .INIT(16'hC480) )  
        \xhdl1.GEN_BITS[5].APB_32.INTR_reg_74_0_0_0_tz[5]  (.A(
        \CONFIG_reg[5][7] ), .B(\CONFIG_reg[5][3] ), .C(
        \INTR_reg_74_0_0_0_tz_1[5] ), .D(N_5940), .Y(
        \INTR_reg_74_0_0_0_tz[5] ));
    CFG3 #( .INIT(8'hFB) )  edge_both_2_sqmuxa_15_i_0 (.A(edge_N_5_mux)
        , .B(\CONFIG_reg[0][3] ), .C(N_141_i), .Y(N_80));
    SLE \xhdl1.GEN_BITS[10].REG_GEN.CONFIG_reg[10][0]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[0]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[10]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[10][0] ));
    SLE \xhdl1.GEN_BITS[14].APB_32.INTR_reg[14]  (.D(
        \INTR_reg_191[14] ), .CLK(FCCC_0_GL1), .EN(VCC_net_1), .ALn(
        MSS_RESET_N_F2M_c), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(INTR_reg_14));
    SLE \xhdl1.GEN_BITS[24].APB_32.GPOUT_reg[24]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[24]), .CLK(FCCC_0_GL1), .EN(
        GPOUT_reg_0_sqmuxa), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        GPOUT_reg_24));
    SLE \xhdl1.GEN_BITS[17].REG_GEN.CONFIG_reg[17][5]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[5]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[17]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[17][5] ));
    CFG4 #( .INIT(16'hF2F3) )  
        \xhdl1.GEN_BITS[16].APB_32.INTR_reg_217_0_o2_1_0[16]  (.A(
        \CONFIG_reg[16][6] ), .B(\edge_neg[16] ), .C(
        \INTR_reg_217_0_o2_0[16] ), .D(\CONFIG_reg[16][5] ), .Y(
        \INTR_reg_217_0_o2_1[16] ));
    SLE \xhdl1.GEN_BITS[1].APB_32.edge_pos[1]  (.D(N_107), .CLK(
        FCCC_0_GL1), .EN(N_66), .ALn(MSS_RESET_N_F2M_c), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(\edge_pos[1] ));
    CFG4 #( .INIT(16'h0A33) )  
        \xhdl1.GEN_BITS[9].APB_32.INTR_reg_126_0[9]  (.A(INTR_reg_9), 
        .B(\INTR_reg_126_0_o2_1[9] ), .C(
        CoreAPB3_0_APBmslave2_PWDATA[9]), .D(edge_N_5_mux), .Y(
        \INTR_reg_126[9] ));
    CFG4 #( .INIT(16'h0F35) )  
        \xhdl1.GEN_BITS[21].REG_GEN.CONFIG_reg[21]_RNIA4H61[4]  (.A(
        \CONFIG_reg[5][4] ), .B(\CONFIG_reg[21][4] ), .C(
        CoreAPB3_0_APBmslave2_PADDR[6]), .D(
        CoreAPB3_0_APBmslave2_PADDR[5]), .Y(\CONFIG_reg_o_2_21_1[4] ));
    CFG2 #( .INIT(4'h8) )  
        \xhdl1.GEN_BITS[4].REG_GEN.CONFIG_reg[4]2_0_a4_0_a2  (.A(N_678)
        , .B(N_603), .Y(\CONFIG_reg[4]2 ));
    CFG4 #( .INIT(16'h0F35) )  
        \xhdl1.GEN_BITS[19].REG_GEN.CONFIG_reg[19]_RNICN391[0]  (.A(
        \CONFIG_reg[3][0] ), .B(\CONFIG_reg[19][0] ), .C(
        CoreAPB3_0_APBmslave2_PADDR[6]), .D(
        CoreAPB3_0_APBmslave2_PADDR[5]), .Y(\CONFIG_reg_o_2_25_1_1[0] )
        );
    CFG4 #( .INIT(16'h0A33) )  
        \xhdl1.GEN_BITS[12].APB_32.INTR_reg_165_0[12]  (.A(INTR_reg_12)
        , .B(\INTR_reg_165_0_o2_1[12] ), .C(
        CoreAPB3_0_APBmslave2_PWDATA[12]), .D(edge_N_5_mux), .Y(
        \INTR_reg_165[12] ));
    CFG4 #( .INIT(16'h8000) )  
        \xhdl1.GEN_BITS[3].REG_GEN.CONFIG_reg[3]2_0_a4_0_a2  (.A(
        CoreAPB3_0_APBmslave2_PADDR[3]), .B(
        CoreAPB3_0_APBmslave2_PADDR[2]), .C(N_604), .D(N_606), .Y(
        \CONFIG_reg[3]2 ));
    SLE \xhdl1.GEN_BITS[12].REG_GEN.CONFIG_reg[12][7]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[7]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[12]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[12][7] ));
    CFG4 #( .INIT(16'hAC0F) )  
        \xhdl1.GEN_BITS[24].REG_GEN.CONFIG_reg[24]_RNIASQ22[2]  (.A(
        \CONFIG_reg[8][2] ), .B(\CONFIG_reg[24][2] ), .C(
        \CONFIG_reg_o_2_3_1_1[2] ), .D(CoreAPB3_0_APBmslave2_PADDR[5]), 
        .Y(N_4677));
    CFG4 #( .INIT(16'hAC0F) )  
        \xhdl1.GEN_BITS[9].REG_GEN.CONFIG_reg[9]_RNIAEU72[0]  (.A(
        \CONFIG_reg[9][0] ), .B(\CONFIG_reg[25][0] ), .C(
        \CONFIG_reg_o_2_18_1[0] ), .D(CoreAPB3_0_APBmslave2_PADDR[5]), 
        .Y(N_4795));
    SLE \xhdl1.GEN_BITS[31].REG_GEN.CONFIG_reg[31][3]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[3]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[31]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[31][3] ));
    SLE \xhdl1.GEN_BITS[11].APB_32.GPOUT_reg[11]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[11]), .CLK(FCCC_0_GL1), .EN(
        GPOUT_reg_0_sqmuxa), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        GPOUT_reg_11));
    SLE \xhdl1.GEN_BITS[31].REG_GEN.CONFIG_reg[31][2]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[2]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[31]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[31][2] ));
    CFG4 #( .INIT(16'hAC0F) )  
        \xhdl1.GEN_BITS[15].REG_GEN.CONFIG_reg[15]_RNI8JN32[1]  (.A(
        \CONFIG_reg[15][1] ), .B(\CONFIG_reg[31][1] ), .C(
        \CONFIG_reg_o_2_28_1_1[1] ), .D(CoreAPB3_0_APBmslave2_PADDR[5])
        , .Y(N_4876));
    CFG4 #( .INIT(16'hA9FF) )  
        \xhdl1.GEN_BITS[16].APB_32.INTR_reg_217_0_o2_0_0[16]  (.A(
        \CONFIG_reg[16][7] ), .B(\CONFIG_reg[16][6] ), .C(
        \CONFIG_reg[16][5] ), .D(\CONFIG_reg[16][3] ), .Y(
        \INTR_reg_217_0_o2_0[16] ));
    CFG2 #( .INIT(4'h1) )  
        \xhdl1.GEN_BITS[0].REG_GEN.CONFIG_reg[0]2_0_a4_0_a2_0  (.A(
        CoreAPB3_0_APBmslave2_PADDR[5]), .B(
        CoreAPB3_0_APBmslave2_PADDR[4]), .Y(N_606));
    CFG4 #( .INIT(16'h0F35) )  
        \xhdl1.GEN_BITS[18].REG_GEN.CONFIG_reg[18]_RNII4I61[5]  (.A(
        \CONFIG_reg[2][5] ), .B(\CONFIG_reg[18][5] ), .C(
        CoreAPB3_0_APBmslave2_PADDR[6]), .D(
        CoreAPB3_0_APBmslave2_PADDR[5]), .Y(\CONFIG_reg_o_2_10_1_1[5] )
        );
    SLE \xhdl1.GEN_BITS[0].REG_GEN.CONFIG_reg[0][0]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[0]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[0]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[0][0] ));
    CFG4 #( .INIT(16'hAC0F) )  
        \xhdl1.GEN_BITS[15].REG_GEN.CONFIG_reg[15]_RNI0CO32[7]  (.A(
        \CONFIG_reg[15][7] ), .B(\CONFIG_reg[31][7] ), .C(
        \CONFIG_reg_o_2_28_1_1[7] ), .D(CoreAPB3_0_APBmslave2_PADDR[5])
        , .Y(N_4882));
    SLE \xhdl1.GEN_BITS[24].REG_GEN.CONFIG_reg[24][4]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[4]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[24]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[24][4] ));
    CFG2 #( .INIT(4'h4) )  edge_neg_2_sqmuxa_10_i_a2 (.A(\gpin2[2] ), 
        .B(gpin3_2), .Y(N_395));
    SLE \xhdl1.GEN_BITS[29].APB_32.edge_both[29]  (.D(
        \edge_neg_415[29] ), .CLK(FCCC_0_GL1), .EN(N_190), .ALn(
        MSS_RESET_N_F2M_c), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(\edge_pos[29] ));
    CFG4 #( .INIT(16'hAC0F) )  
        \xhdl1.GEN_BITS[15].REG_GEN.CONFIG_reg[15]_RNIGRN32[3]  (.A(
        \CONFIG_reg[15][3] ), .B(\CONFIG_reg[31][3] ), .C(
        \CONFIG_reg_o_2_28_1_1[3] ), .D(CoreAPB3_0_APBmslave2_PADDR[5])
        , .Y(N_4878));
    SLE \xhdl1.GEN_BITS[22].REG_GEN.CONFIG_reg[22][7]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[7]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[22]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[22][7] ));
    CFG4 #( .INIT(16'hAC0F) )  
        \xhdl1.GEN_BITS[14].REG_GEN.CONFIG_reg[14]_RNI0OP82[1]  (.A(
        \CONFIG_reg[14][1] ), .B(\CONFIG_reg[30][1] ), .C(
        \CONFIG_reg_o_2_13_1_1[1] ), .D(CoreAPB3_0_APBmslave2_PADDR[5])
        , .Y(N_4756));
    SLE \xhdl1.GEN_BITS[10].REG_GEN.CONFIG_reg[10][4]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[4]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[10]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[10][4] ));
    CFG4 #( .INIT(16'hAC0F) )  
        \xhdl1.GEN_BITS[9].REG_GEN.CONFIG_reg[9]_RNIMQU72[3]  (.A(
        \CONFIG_reg[9][3] ), .B(\CONFIG_reg[25][3] ), .C(
        \CONFIG_reg_o_2_18_1[3] ), .D(CoreAPB3_0_APBmslave2_PADDR[5]), 
        .Y(N_4798));
    SLE \xhdl1.GEN_BITS[14].REG_GEN.CONFIG_reg[14][1]  (.D(
        CoreAPB3_0_APBmslave2_PWDATA[1]), .CLK(FCCC_0_GL1), .EN(
        \CONFIG_reg[14]2 ), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \CONFIG_reg[14][1] ));
    CFG3 #( .INIT(8'h08) )  PRDATA_m1_e_1_inst_1 (.A(
        CoreAPB3_0_APBmslave2_PADDR[5]), .B(\GPOUT_reg[7] ), .C(
        CoreAPB3_0_APBmslave2_PADDR[4]), .Y(PRDATA_m1_e_1));
    CFG4 #( .INIT(16'hA820) )  
        \xhdl1.GEN_BITS[3].REG_INT.un34_intr_u_ns  (.A(
        \CONFIG_reg[3][3] ), .B(\CONFIG_reg[3][7] ), .C(un34_intr_u_bm)
        , .D(un34_intr_u_ns_1), .Y(un34_intr));
    CFG3 #( .INIT(8'hFB) )  edge_neg_2_sqmuxa_25_i_0 (.A(edge_N_5_mux), 
        .B(\CONFIG_reg[0][3] ), .C(N_401), .Y(N_52));
    SLE \xhdl1.GEN_BITS[0].gpin2[0]  (.D(\gpin1[0] ), .CLK(FCCC_0_GL1), 
        .EN(VCC_net_1), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(\gpin2[0] ));
    
endmodule


module FIC_COREAPBLSRAM_0_lsram_512to35328x32_512s_32s(
       lsram_width32_PRDATA,
       CoreAPB3_0_APBmslave2_PADDR,
       CoreAPB3_0_APBmslave2_PWDATA,
       FCCC_0_GL1,
       MSS_RESET_N_F2M_c,
       wen
    );
output [31:0] lsram_width32_PRDATA;
input  [8:0] CoreAPB3_0_APBmslave2_PADDR;
input  [31:0] CoreAPB3_0_APBmslave2_PWDATA;
input  FCCC_0_GL1;
input  MSS_RESET_N_F2M_c;
input  wen;

    wire VCC_net_1, GND_net_1;
    
    RAM1K18 block0 (.A_DOUT({nc0, lsram_width32_PRDATA[15], 
        lsram_width32_PRDATA[14], lsram_width32_PRDATA[13], 
        lsram_width32_PRDATA[12], lsram_width32_PRDATA[11], 
        lsram_width32_PRDATA[10], lsram_width32_PRDATA[9], 
        lsram_width32_PRDATA[8], nc1, lsram_width32_PRDATA[7], 
        lsram_width32_PRDATA[6], lsram_width32_PRDATA[5], 
        lsram_width32_PRDATA[4], lsram_width32_PRDATA[3], 
        lsram_width32_PRDATA[2], lsram_width32_PRDATA[1], 
        lsram_width32_PRDATA[0]}), .B_DOUT({nc2, 
        lsram_width32_PRDATA[31], lsram_width32_PRDATA[30], 
        lsram_width32_PRDATA[29], lsram_width32_PRDATA[28], 
        lsram_width32_PRDATA[27], lsram_width32_PRDATA[26], 
        lsram_width32_PRDATA[25], lsram_width32_PRDATA[24], nc3, 
        lsram_width32_PRDATA[23], lsram_width32_PRDATA[22], 
        lsram_width32_PRDATA[21], lsram_width32_PRDATA[20], 
        lsram_width32_PRDATA[19], lsram_width32_PRDATA[18], 
        lsram_width32_PRDATA[17], lsram_width32_PRDATA[16]}), .BUSY(), 
        .A_CLK(FCCC_0_GL1), .A_DOUT_CLK(VCC_net_1), .A_ARST_N(
        MSS_RESET_N_F2M_c), .A_DOUT_EN(VCC_net_1), .A_BLK({VCC_net_1, 
        VCC_net_1, VCC_net_1}), .A_DOUT_ARST_N(VCC_net_1), 
        .A_DOUT_SRST_N(VCC_net_1), .A_DIN({GND_net_1, 
        CoreAPB3_0_APBmslave2_PWDATA[15], 
        CoreAPB3_0_APBmslave2_PWDATA[14], 
        CoreAPB3_0_APBmslave2_PWDATA[13], 
        CoreAPB3_0_APBmslave2_PWDATA[12], 
        CoreAPB3_0_APBmslave2_PWDATA[11], 
        CoreAPB3_0_APBmslave2_PWDATA[10], 
        CoreAPB3_0_APBmslave2_PWDATA[9], 
        CoreAPB3_0_APBmslave2_PWDATA[8], GND_net_1, 
        CoreAPB3_0_APBmslave2_PWDATA[7], 
        CoreAPB3_0_APBmslave2_PWDATA[6], 
        CoreAPB3_0_APBmslave2_PWDATA[5], 
        CoreAPB3_0_APBmslave2_PWDATA[4], 
        CoreAPB3_0_APBmslave2_PWDATA[3], 
        CoreAPB3_0_APBmslave2_PWDATA[2], 
        CoreAPB3_0_APBmslave2_PWDATA[1], 
        CoreAPB3_0_APBmslave2_PWDATA[0]}), .A_ADDR({
        CoreAPB3_0_APBmslave2_PADDR[8], CoreAPB3_0_APBmslave2_PADDR[7], 
        CoreAPB3_0_APBmslave2_PADDR[6], CoreAPB3_0_APBmslave2_PADDR[5], 
        CoreAPB3_0_APBmslave2_PADDR[4], CoreAPB3_0_APBmslave2_PADDR[3], 
        CoreAPB3_0_APBmslave2_PADDR[2], CoreAPB3_0_APBmslave2_PADDR[1], 
        CoreAPB3_0_APBmslave2_PADDR[0], GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1}), .A_WEN({wen, wen}), .B_CLK(
        FCCC_0_GL1), .B_DOUT_CLK(VCC_net_1), .B_ARST_N(
        MSS_RESET_N_F2M_c), .B_DOUT_EN(VCC_net_1), .B_BLK({VCC_net_1, 
        VCC_net_1, VCC_net_1}), .B_DOUT_ARST_N(VCC_net_1), 
        .B_DOUT_SRST_N(VCC_net_1), .B_DIN({GND_net_1, 
        CoreAPB3_0_APBmslave2_PWDATA[31], 
        CoreAPB3_0_APBmslave2_PWDATA[30], 
        CoreAPB3_0_APBmslave2_PWDATA[29], 
        CoreAPB3_0_APBmslave2_PWDATA[28], 
        CoreAPB3_0_APBmslave2_PWDATA[27], 
        CoreAPB3_0_APBmslave2_PWDATA[26], 
        CoreAPB3_0_APBmslave2_PWDATA[25], 
        CoreAPB3_0_APBmslave2_PWDATA[24], GND_net_1, 
        CoreAPB3_0_APBmslave2_PWDATA[23], 
        CoreAPB3_0_APBmslave2_PWDATA[22], 
        CoreAPB3_0_APBmslave2_PWDATA[21], 
        CoreAPB3_0_APBmslave2_PWDATA[20], 
        CoreAPB3_0_APBmslave2_PWDATA[19], 
        CoreAPB3_0_APBmslave2_PWDATA[18], 
        CoreAPB3_0_APBmslave2_PWDATA[17], 
        CoreAPB3_0_APBmslave2_PWDATA[16]}), .B_ADDR({
        CoreAPB3_0_APBmslave2_PADDR[8], CoreAPB3_0_APBmslave2_PADDR[7], 
        CoreAPB3_0_APBmslave2_PADDR[6], CoreAPB3_0_APBmslave2_PADDR[5], 
        CoreAPB3_0_APBmslave2_PADDR[4], CoreAPB3_0_APBmslave2_PADDR[3], 
        CoreAPB3_0_APBmslave2_PADDR[2], CoreAPB3_0_APBmslave2_PADDR[1], 
        CoreAPB3_0_APBmslave2_PADDR[0], GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1}), .B_WEN({wen, wen}), .A_EN(
        VCC_net_1), .A_DOUT_LAT(VCC_net_1), .A_WIDTH({VCC_net_1, 
        GND_net_1, VCC_net_1}), .A_WMODE(GND_net_1), .B_EN(VCC_net_1), 
        .B_DOUT_LAT(VCC_net_1), .B_WIDTH({VCC_net_1, GND_net_1, 
        VCC_net_1}), .B_WMODE(GND_net_1), .SII_LOCK(GND_net_1));
    VCC VCC (.Y(VCC_net_1));
    GND GND (.Y(GND_net_1));
    
endmodule


module FIC_COREAPBLSRAM_0_COREAPBLSRAM_Z2(
       PRDATA_reg,
       lsram_width32_PRDATA,
       CoreAPB3_0_APBmslave2_PADDR,
       CoreAPB3_0_APBmslave2_PWDATA,
       MSS_RESET_N_F2M_c,
       FCCC_0_GL1,
       CoreAPB3_0_APBmslave2_PREADY,
       CoreAPB3_0_APBmslave2_PENABLE,
       CoreAPB3_0_APBmslave2_PWRITE,
       wen_0,
       PRDATA4_out,
       iPRDATA29
    );
output [31:0] PRDATA_reg;
output [31:0] lsram_width32_PRDATA;
input  [8:0] CoreAPB3_0_APBmslave2_PADDR;
input  [31:0] CoreAPB3_0_APBmslave2_PWDATA;
input  MSS_RESET_N_F2M_c;
input  FCCC_0_GL1;
output CoreAPB3_0_APBmslave2_PREADY;
input  CoreAPB3_0_APBmslave2_PENABLE;
input  CoreAPB3_0_APBmslave2_PWRITE;
output wen_0;
output PRDATA4_out;
input  iPRDATA29;

    wire VCC_net_1, PRDATA4_net_1, GND_net_1, PREADY_reg6_i_0, 
        wen_net_1;
    
    SLE \PRDATA_reg[13]  (.D(lsram_width32_PRDATA[13]), .CLK(
        FCCC_0_GL1), .EN(PRDATA4_net_1), .ALn(MSS_RESET_N_F2M_c), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(PRDATA_reg[13]));
    FIC_COREAPBLSRAM_0_lsram_512to35328x32_512s_32s 
        \genblk1.genblk1.lsram_512to35328x32_block0  (
        .lsram_width32_PRDATA({lsram_width32_PRDATA[31], 
        lsram_width32_PRDATA[30], lsram_width32_PRDATA[29], 
        lsram_width32_PRDATA[28], lsram_width32_PRDATA[27], 
        lsram_width32_PRDATA[26], lsram_width32_PRDATA[25], 
        lsram_width32_PRDATA[24], lsram_width32_PRDATA[23], 
        lsram_width32_PRDATA[22], lsram_width32_PRDATA[21], 
        lsram_width32_PRDATA[20], lsram_width32_PRDATA[19], 
        lsram_width32_PRDATA[18], lsram_width32_PRDATA[17], 
        lsram_width32_PRDATA[16], lsram_width32_PRDATA[15], 
        lsram_width32_PRDATA[14], lsram_width32_PRDATA[13], 
        lsram_width32_PRDATA[12], lsram_width32_PRDATA[11], 
        lsram_width32_PRDATA[10], lsram_width32_PRDATA[9], 
        lsram_width32_PRDATA[8], lsram_width32_PRDATA[7], 
        lsram_width32_PRDATA[6], lsram_width32_PRDATA[5], 
        lsram_width32_PRDATA[4], lsram_width32_PRDATA[3], 
        lsram_width32_PRDATA[2], lsram_width32_PRDATA[1], 
        lsram_width32_PRDATA[0]}), .CoreAPB3_0_APBmslave2_PADDR({
        CoreAPB3_0_APBmslave2_PADDR[8], CoreAPB3_0_APBmslave2_PADDR[7], 
        CoreAPB3_0_APBmslave2_PADDR[6], CoreAPB3_0_APBmslave2_PADDR[5], 
        CoreAPB3_0_APBmslave2_PADDR[4], CoreAPB3_0_APBmslave2_PADDR[3], 
        CoreAPB3_0_APBmslave2_PADDR[2], CoreAPB3_0_APBmslave2_PADDR[1], 
        CoreAPB3_0_APBmslave2_PADDR[0]}), 
        .CoreAPB3_0_APBmslave2_PWDATA({
        CoreAPB3_0_APBmslave2_PWDATA[31], 
        CoreAPB3_0_APBmslave2_PWDATA[30], 
        CoreAPB3_0_APBmslave2_PWDATA[29], 
        CoreAPB3_0_APBmslave2_PWDATA[28], 
        CoreAPB3_0_APBmslave2_PWDATA[27], 
        CoreAPB3_0_APBmslave2_PWDATA[26], 
        CoreAPB3_0_APBmslave2_PWDATA[25], 
        CoreAPB3_0_APBmslave2_PWDATA[24], 
        CoreAPB3_0_APBmslave2_PWDATA[23], 
        CoreAPB3_0_APBmslave2_PWDATA[22], 
        CoreAPB3_0_APBmslave2_PWDATA[21], 
        CoreAPB3_0_APBmslave2_PWDATA[20], 
        CoreAPB3_0_APBmslave2_PWDATA[19], 
        CoreAPB3_0_APBmslave2_PWDATA[18], 
        CoreAPB3_0_APBmslave2_PWDATA[17], 
        CoreAPB3_0_APBmslave2_PWDATA[16], 
        CoreAPB3_0_APBmslave2_PWDATA[15], 
        CoreAPB3_0_APBmslave2_PWDATA[14], 
        CoreAPB3_0_APBmslave2_PWDATA[13], 
        CoreAPB3_0_APBmslave2_PWDATA[12], 
        CoreAPB3_0_APBmslave2_PWDATA[11], 
        CoreAPB3_0_APBmslave2_PWDATA[10], 
        CoreAPB3_0_APBmslave2_PWDATA[9], 
        CoreAPB3_0_APBmslave2_PWDATA[8], 
        CoreAPB3_0_APBmslave2_PWDATA[7], 
        CoreAPB3_0_APBmslave2_PWDATA[6], 
        CoreAPB3_0_APBmslave2_PWDATA[5], 
        CoreAPB3_0_APBmslave2_PWDATA[4], 
        CoreAPB3_0_APBmslave2_PWDATA[3], 
        CoreAPB3_0_APBmslave2_PWDATA[2], 
        CoreAPB3_0_APBmslave2_PWDATA[1], 
        CoreAPB3_0_APBmslave2_PWDATA[0]}), .FCCC_0_GL1(FCCC_0_GL1), 
        .MSS_RESET_N_F2M_c(MSS_RESET_N_F2M_c), .wen(wen_net_1));
    SLE \PRDATA_reg[26]  (.D(lsram_width32_PRDATA[26]), .CLK(
        FCCC_0_GL1), .EN(PRDATA4_net_1), .ALn(MSS_RESET_N_F2M_c), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(PRDATA_reg[26]));
    CFG2 #( .INIT(4'h8) )  wen_0_inst_1 (.A(
        CoreAPB3_0_APBmslave2_PENABLE), .B(
        CoreAPB3_0_APBmslave2_PWRITE), .Y(wen_0));
    SLE \PRDATA_reg[6]  (.D(lsram_width32_PRDATA[6]), .CLK(FCCC_0_GL1), 
        .EN(PRDATA4_net_1), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        PRDATA_reg[6]));
    SLE \PRDATA_reg[14]  (.D(lsram_width32_PRDATA[14]), .CLK(
        FCCC_0_GL1), .EN(PRDATA4_net_1), .ALn(MSS_RESET_N_F2M_c), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(PRDATA_reg[14]));
    SLE \PRDATA_reg[17]  (.D(lsram_width32_PRDATA[17]), .CLK(
        FCCC_0_GL1), .EN(PRDATA4_net_1), .ALn(MSS_RESET_N_F2M_c), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(PRDATA_reg[17]));
    SLE \PRDATA_reg[15]  (.D(lsram_width32_PRDATA[15]), .CLK(
        FCCC_0_GL1), .EN(PRDATA4_net_1), .ALn(MSS_RESET_N_F2M_c), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(PRDATA_reg[15]));
    VCC VCC (.Y(VCC_net_1));
    SLE \PRDATA_reg[9]  (.D(lsram_width32_PRDATA[9]), .CLK(FCCC_0_GL1), 
        .EN(PRDATA4_net_1), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        PRDATA_reg[9]));
    CFG2 #( .INIT(4'h8) )  PRDATA4 (.A(iPRDATA29), .B(PRDATA4_out), .Y(
        PRDATA4_net_1));
    SLE \PRDATA_reg[10]  (.D(lsram_width32_PRDATA[10]), .CLK(
        FCCC_0_GL1), .EN(PRDATA4_net_1), .ALn(MSS_RESET_N_F2M_c), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(PRDATA_reg[10]));
    SLE \PRDATA_reg[23]  (.D(lsram_width32_PRDATA[23]), .CLK(
        FCCC_0_GL1), .EN(PRDATA4_net_1), .ALn(MSS_RESET_N_F2M_c), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(PRDATA_reg[23]));
    CFG2 #( .INIT(4'h8) )  wen (.A(iPRDATA29), .B(wen_0), .Y(wen_net_1)
        );
    SLE \PRDATA_reg[4]  (.D(lsram_width32_PRDATA[4]), .CLK(FCCC_0_GL1), 
        .EN(PRDATA4_net_1), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        PRDATA_reg[4]));
    GND GND (.Y(GND_net_1));
    SLE \PRDATA_reg[24]  (.D(lsram_width32_PRDATA[24]), .CLK(
        FCCC_0_GL1), .EN(PRDATA4_net_1), .ALn(MSS_RESET_N_F2M_c), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(PRDATA_reg[24]));
    SLE \PRDATA_reg[27]  (.D(lsram_width32_PRDATA[27]), .CLK(
        FCCC_0_GL1), .EN(PRDATA4_net_1), .ALn(MSS_RESET_N_F2M_c), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(PRDATA_reg[27]));
    SLE \PRDATA_reg[19]  (.D(lsram_width32_PRDATA[19]), .CLK(
        FCCC_0_GL1), .EN(PRDATA4_net_1), .ALn(MSS_RESET_N_F2M_c), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(PRDATA_reg[19]));
    SLE \PRDATA_reg[2]  (.D(lsram_width32_PRDATA[2]), .CLK(FCCC_0_GL1), 
        .EN(PRDATA4_net_1), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        PRDATA_reg[2]));
    SLE \PRDATA_reg[25]  (.D(lsram_width32_PRDATA[25]), .CLK(
        FCCC_0_GL1), .EN(PRDATA4_net_1), .ALn(MSS_RESET_N_F2M_c), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(PRDATA_reg[25]));
    SLE \PRDATA_reg[3]  (.D(lsram_width32_PRDATA[3]), .CLK(FCCC_0_GL1), 
        .EN(PRDATA4_net_1), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        PRDATA_reg[3]));
    SLE \PRDATA_reg[11]  (.D(lsram_width32_PRDATA[11]), .CLK(
        FCCC_0_GL1), .EN(PRDATA4_net_1), .ALn(MSS_RESET_N_F2M_c), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(PRDATA_reg[11]));
    SLE \PRDATA_reg[18]  (.D(lsram_width32_PRDATA[18]), .CLK(
        FCCC_0_GL1), .EN(PRDATA4_net_1), .ALn(MSS_RESET_N_F2M_c), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(PRDATA_reg[18]));
    SLE \PRDATA_reg[20]  (.D(lsram_width32_PRDATA[20]), .CLK(
        FCCC_0_GL1), .EN(PRDATA4_net_1), .ALn(MSS_RESET_N_F2M_c), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(PRDATA_reg[20]));
    SLE \PRDATA_reg[30]  (.D(lsram_width32_PRDATA[30]), .CLK(
        FCCC_0_GL1), .EN(PRDATA4_net_1), .ALn(MSS_RESET_N_F2M_c), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(PRDATA_reg[30]));
    SLE \PRDATA_reg[12]  (.D(lsram_width32_PRDATA[12]), .CLK(
        FCCC_0_GL1), .EN(PRDATA4_net_1), .ALn(MSS_RESET_N_F2M_c), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(PRDATA_reg[12]));
    CFG4 #( .INIT(16'hFFBF) )  PREADY_reg6_i (.A(
        CoreAPB3_0_APBmslave2_PWRITE), .B(CoreAPB3_0_APBmslave2_PREADY)
        , .C(iPRDATA29), .D(CoreAPB3_0_APBmslave2_PENABLE), .Y(
        PREADY_reg6_i_0));
    SLE \PRDATA_reg[5]  (.D(lsram_width32_PRDATA[5]), .CLK(FCCC_0_GL1), 
        .EN(PRDATA4_net_1), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        PRDATA_reg[5]));
    SLE \PRDATA_reg[1]  (.D(lsram_width32_PRDATA[1]), .CLK(FCCC_0_GL1), 
        .EN(PRDATA4_net_1), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        PRDATA_reg[1]));
    SLE \PRDATA_reg[16]  (.D(lsram_width32_PRDATA[16]), .CLK(
        FCCC_0_GL1), .EN(PRDATA4_net_1), .ALn(MSS_RESET_N_F2M_c), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(PRDATA_reg[16]));
    SLE \PRDATA_reg[8]  (.D(lsram_width32_PRDATA[8]), .CLK(FCCC_0_GL1), 
        .EN(PRDATA4_net_1), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        PRDATA_reg[8]));
    SLE \PRDATA_reg[29]  (.D(lsram_width32_PRDATA[29]), .CLK(
        FCCC_0_GL1), .EN(PRDATA4_net_1), .ALn(MSS_RESET_N_F2M_c), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(PRDATA_reg[29]));
    SLE \PRDATA_reg[0]  (.D(lsram_width32_PRDATA[0]), .CLK(FCCC_0_GL1), 
        .EN(PRDATA4_net_1), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        PRDATA_reg[0]));
    SLE \PRDATA_reg[21]  (.D(lsram_width32_PRDATA[21]), .CLK(
        FCCC_0_GL1), .EN(PRDATA4_net_1), .ALn(MSS_RESET_N_F2M_c), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(PRDATA_reg[21]));
    SLE \PRDATA_reg[31]  (.D(lsram_width32_PRDATA[31]), .CLK(
        FCCC_0_GL1), .EN(PRDATA4_net_1), .ALn(MSS_RESET_N_F2M_c), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(PRDATA_reg[31]));
    SLE \PRDATA_reg[7]  (.D(lsram_width32_PRDATA[7]), .CLK(FCCC_0_GL1), 
        .EN(PRDATA4_net_1), .ALn(MSS_RESET_N_F2M_c), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        PRDATA_reg[7]));
    CFG2 #( .INIT(4'h2) )  PRDATA4_s (.A(CoreAPB3_0_APBmslave2_PENABLE)
        , .B(CoreAPB3_0_APBmslave2_PWRITE), .Y(PRDATA4_out));
    SLE PREADY_reg (.D(PREADY_reg6_i_0), .CLK(FCCC_0_GL1), .EN(
        VCC_net_1), .ALn(MSS_RESET_N_F2M_c), .ADn(GND_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        CoreAPB3_0_APBmslave2_PREADY));
    SLE \PRDATA_reg[28]  (.D(lsram_width32_PRDATA[28]), .CLK(
        FCCC_0_GL1), .EN(PRDATA4_net_1), .ALn(MSS_RESET_N_F2M_c), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(PRDATA_reg[28]));
    SLE \PRDATA_reg[22]  (.D(lsram_width32_PRDATA[22]), .CLK(
        FCCC_0_GL1), .EN(PRDATA4_net_1), .ALn(MSS_RESET_N_F2M_c), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(PRDATA_reg[22]));
    
endmodule


module FIC(
       GPIO_IN,
       GPIO_OUT,
       MMUART_0_RXD,
       MSS_RESET_N_F2M,
       MMUART_0_TXD
    );
input  [0:6] GPIO_IN;
output [0:6] GPIO_OUT;
input  MMUART_0_RXD;
input  MSS_RESET_N_F2M;
output MMUART_0_TXD;

    wire \GPIO_OUT_net_2[6] , \GPIO_OUT_net_2[5] , \GPIO_OUT_net_2[4] , 
        \GPIO_OUT_net_2[3] , \GPIO_OUT_net_2[2] , \GPIO_OUT_net_2[1] , 
        \GPIO_OUT_net_2[0] , GND_net_1, 
        \CoreAPB3_0_APBmslave2_PADDR[0] , 
        \CoreAPB3_0_APBmslave2_PADDR[1] , 
        \CoreAPB3_0_APBmslave2_PADDR[2] , 
        \CoreAPB3_0_APBmslave2_PADDR[3] , 
        \CoreAPB3_0_APBmslave2_PADDR[4] , 
        \CoreAPB3_0_APBmslave2_PADDR[5] , 
        \CoreAPB3_0_APBmslave2_PADDR[6] , 
        \CoreAPB3_0_APBmslave2_PADDR[7] , 
        \CoreAPB3_0_APBmslave2_PADDR[8] , 
        \FIC_MSS_0_FIC_0_APB_MASTER_PADDR[28] , 
        \FIC_MSS_0_FIC_0_APB_MASTER_PADDR[29] , 
        \FIC_MSS_0_FIC_0_APB_MASTER_PADDR[30] , 
        \FIC_MSS_0_FIC_0_APB_MASTER_PADDR[31] , 
        CoreAPB3_0_APBmslave2_PWRITE, CoreAPB3_0_APBmslave2_PENABLE, 
        FIC_MSS_0_FIC_0_APB_MASTER_PSELx, 
        \CoreAPB3_0_APBmslave2_PWDATA[0] , 
        \CoreAPB3_0_APBmslave2_PWDATA[1] , 
        \CoreAPB3_0_APBmslave2_PWDATA[2] , 
        \CoreAPB3_0_APBmslave2_PWDATA[3] , 
        \CoreAPB3_0_APBmslave2_PWDATA[4] , 
        \CoreAPB3_0_APBmslave2_PWDATA[5] , 
        \CoreAPB3_0_APBmslave2_PWDATA[6] , 
        \CoreAPB3_0_APBmslave2_PWDATA[7] , 
        \CoreAPB3_0_APBmslave2_PWDATA[8] , 
        \CoreAPB3_0_APBmslave2_PWDATA[9] , 
        \CoreAPB3_0_APBmslave2_PWDATA[10] , 
        \CoreAPB3_0_APBmslave2_PWDATA[11] , 
        \CoreAPB3_0_APBmslave2_PWDATA[12] , 
        \CoreAPB3_0_APBmslave2_PWDATA[13] , 
        \CoreAPB3_0_APBmslave2_PWDATA[14] , 
        \CoreAPB3_0_APBmslave2_PWDATA[15] , 
        \CoreAPB3_0_APBmslave2_PWDATA[16] , 
        \CoreAPB3_0_APBmslave2_PWDATA[17] , 
        \CoreAPB3_0_APBmslave2_PWDATA[18] , 
        \CoreAPB3_0_APBmslave2_PWDATA[19] , 
        \CoreAPB3_0_APBmslave2_PWDATA[20] , 
        \CoreAPB3_0_APBmslave2_PWDATA[21] , 
        \CoreAPB3_0_APBmslave2_PWDATA[22] , 
        \CoreAPB3_0_APBmslave2_PWDATA[23] , 
        \CoreAPB3_0_APBmslave2_PWDATA[24] , 
        \CoreAPB3_0_APBmslave2_PWDATA[25] , 
        \CoreAPB3_0_APBmslave2_PWDATA[26] , 
        \CoreAPB3_0_APBmslave2_PWDATA[27] , 
        \CoreAPB3_0_APBmslave2_PWDATA[28] , 
        \CoreAPB3_0_APBmslave2_PWDATA[29] , 
        \CoreAPB3_0_APBmslave2_PWDATA[30] , 
        \CoreAPB3_0_APBmslave2_PWDATA[31] , 
        \FIC_MSS_0_FIC_0_APB_MASTER_PRDATA[3] , 
        \FIC_MSS_0_FIC_0_APB_MASTER_PRDATA[4] , 
        \FIC_MSS_0_FIC_0_APB_MASTER_PRDATA[7] , 
        \FIC_MSS_0_FIC_0_APB_MASTER_PRDATA[8] , 
        \FIC_MSS_0_FIC_0_APB_MASTER_PRDATA[9] , 
        \FIC_MSS_0_FIC_0_APB_MASTER_PRDATA[10] , 
        \FIC_MSS_0_FIC_0_APB_MASTER_PRDATA[11] , 
        \FIC_MSS_0_FIC_0_APB_MASTER_PRDATA[12] , 
        \FIC_MSS_0_FIC_0_APB_MASTER_PRDATA[13] , 
        \FIC_MSS_0_FIC_0_APB_MASTER_PRDATA[14] , 
        \FIC_MSS_0_FIC_0_APB_MASTER_PRDATA[15] , 
        \FIC_MSS_0_FIC_0_APB_MASTER_PRDATA[16] , 
        \FIC_MSS_0_FIC_0_APB_MASTER_PRDATA[17] , 
        \FIC_MSS_0_FIC_0_APB_MASTER_PRDATA[18] , 
        \FIC_MSS_0_FIC_0_APB_MASTER_PRDATA[19] , 
        \FIC_MSS_0_FIC_0_APB_MASTER_PRDATA[20] , 
        \FIC_MSS_0_FIC_0_APB_MASTER_PRDATA[21] , 
        \FIC_MSS_0_FIC_0_APB_MASTER_PRDATA[22] , 
        \FIC_MSS_0_FIC_0_APB_MASTER_PRDATA[23] , 
        \FIC_MSS_0_FIC_0_APB_MASTER_PRDATA[24] , 
        \FIC_MSS_0_FIC_0_APB_MASTER_PRDATA[25] , 
        \FIC_MSS_0_FIC_0_APB_MASTER_PRDATA[26] , 
        \FIC_MSS_0_FIC_0_APB_MASTER_PRDATA[27] , 
        \FIC_MSS_0_FIC_0_APB_MASTER_PRDATA[28] , 
        \FIC_MSS_0_FIC_0_APB_MASTER_PRDATA[29] , 
        \FIC_MSS_0_FIC_0_APB_MASTER_PRDATA[30] , 
        \FIC_MSS_0_FIC_0_APB_MASTER_PRDATA[31] , 
        \CoreAPB3_0_APBmslave3_PRDATA[0] , 
        \CoreAPB3_0_APBmslave3_PRDATA[1] , 
        \CoreAPB3_0_APBmslave3_PRDATA[2] , 
        \CoreAPB3_0_APBmslave3_PRDATA[3] , 
        \CoreAPB3_0_APBmslave3_PRDATA[4] , 
        \CoreAPB3_0_APBmslave3_PRDATA[5] , 
        \CoreAPB3_0_APBmslave3_PRDATA[6] , 
        \CoreAPB3_0_APBmslave3_PRDATA[7] , 
        CoreAPB3_0_APBmslave2_PREADY, CoreAPB3_0_APBmslave3_PREADY, 
        FCCC_0_GL1, OSC_0_RCOSC_25_50MHZ_CCC_OUT_RCOSC_25_50MHZ_CCC, 
        FCCC_0_LOCK, VCC_net_1, 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[0] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[1] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[2] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[3] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[4] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[5] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[6] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[7] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[8] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[9] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[10] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[11] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[12] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[13] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[14] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[15] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[16] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[17] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[18] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[19] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[20] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[21] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[22] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[23] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[24] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[25] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[26] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[27] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[28] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[29] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[30] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[31] , 
        \COREAPBLSRAM_0.PRDATA_reg[0] , \COREAPBLSRAM_0.PRDATA_reg[1] , 
        \COREAPBLSRAM_0.PRDATA_reg[2] , \COREAPBLSRAM_0.PRDATA_reg[3] , 
        \COREAPBLSRAM_0.PRDATA_reg[4] , \COREAPBLSRAM_0.PRDATA_reg[5] , 
        \COREAPBLSRAM_0.PRDATA_reg[6] , \COREAPBLSRAM_0.PRDATA_reg[7] , 
        \COREAPBLSRAM_0.PRDATA_reg[8] , \COREAPBLSRAM_0.PRDATA_reg[9] , 
        \COREAPBLSRAM_0.PRDATA_reg[10] , 
        \COREAPBLSRAM_0.PRDATA_reg[11] , 
        \COREAPBLSRAM_0.PRDATA_reg[12] , 
        \COREAPBLSRAM_0.PRDATA_reg[13] , 
        \COREAPBLSRAM_0.PRDATA_reg[14] , 
        \COREAPBLSRAM_0.PRDATA_reg[15] , 
        \COREAPBLSRAM_0.PRDATA_reg[16] , 
        \COREAPBLSRAM_0.PRDATA_reg[17] , 
        \COREAPBLSRAM_0.PRDATA_reg[18] , 
        \COREAPBLSRAM_0.PRDATA_reg[19] , 
        \COREAPBLSRAM_0.PRDATA_reg[20] , 
        \COREAPBLSRAM_0.PRDATA_reg[21] , 
        \COREAPBLSRAM_0.PRDATA_reg[22] , 
        \COREAPBLSRAM_0.PRDATA_reg[23] , 
        \COREAPBLSRAM_0.PRDATA_reg[24] , 
        \COREAPBLSRAM_0.PRDATA_reg[25] , 
        \COREAPBLSRAM_0.PRDATA_reg[26] , 
        \COREAPBLSRAM_0.PRDATA_reg[27] , 
        \COREAPBLSRAM_0.PRDATA_reg[28] , 
        \COREAPBLSRAM_0.PRDATA_reg[29] , 
        \COREAPBLSRAM_0.PRDATA_reg[30] , 
        \COREAPBLSRAM_0.PRDATA_reg[31] , 
        \CoreGPIO_0.xhdl1.GEN_BITS[0].gpin3[0] , 
        \CoreGPIO_0.xhdl1.GEN_BITS[1].gpin3[1] , 
        \CoreGPIO_0.xhdl1.GEN_BITS[2].gpin3[2] , 
        \CoreGPIO_0.xhdl1.GEN_BITS[3].gpin3[3] , 
        \CoreGPIO_0.xhdl1.GEN_BITS[5].gpin3[5] , 
        \CoreGPIO_0.xhdl1.GEN_BITS[6].gpin3[6] , 
        \CoreGPIO_0.xhdl1.GEN_BITS[0].APB_32.INTR_reg[0] , 
        \CoreGPIO_0.xhdl1.GEN_BITS[1].APB_32.INTR_reg[1] , 
        \CoreGPIO_0.xhdl1.GEN_BITS[2].APB_32.INTR_reg[2] , 
        \CoreGPIO_0.xhdl1.GEN_BITS[4].APB_32.INTR_reg[4] , 
        \CoreGPIO_0.xhdl1.GEN_BITS[5].APB_32.INTR_reg[5] , 
        \CoreGPIO_0.xhdl1.GEN_BITS[6].APB_32.INTR_reg[6] , 
        \CoreGPIO_0.xhdl1.GEN_BITS[7].APB_32.INTR_reg[7] , 
        \CoreGPIO_0.xhdl1.GEN_BITS[8].APB_32.INTR_reg[8] , 
        \CoreGPIO_0.xhdl1.GEN_BITS[9].APB_32.INTR_reg[9] , 
        \CoreGPIO_0.xhdl1.GEN_BITS[10].APB_32.INTR_reg[10] , 
        \CoreGPIO_0.xhdl1.GEN_BITS[11].APB_32.INTR_reg[11] , 
        \CoreGPIO_0.xhdl1.GEN_BITS[12].APB_32.INTR_reg[12] , 
        \CoreGPIO_0.xhdl1.GEN_BITS[13].APB_32.INTR_reg[13] , 
        \CoreGPIO_0.xhdl1.GEN_BITS[14].APB_32.INTR_reg[14] , 
        \CoreGPIO_0.xhdl1.GEN_BITS[15].APB_32.INTR_reg[15] , 
        \CoreGPIO_0.xhdl1.GEN_BITS[16].APB_32.INTR_reg[16] , 
        \CoreGPIO_0.xhdl1.GEN_BITS[17].APB_32.INTR_reg[17] , 
        \CoreGPIO_0.xhdl1.GEN_BITS[18].APB_32.INTR_reg[18] , 
        \CoreGPIO_0.xhdl1.GEN_BITS[19].APB_32.INTR_reg[19] , 
        \CoreGPIO_0.xhdl1.GEN_BITS[20].APB_32.INTR_reg[20] , 
        \CoreGPIO_0.xhdl1.GEN_BITS[21].APB_32.INTR_reg[21] , 
        \CoreGPIO_0.xhdl1.GEN_BITS[22].APB_32.INTR_reg[22] , 
        \CoreGPIO_0.xhdl1.GEN_BITS[23].APB_32.INTR_reg[23] , 
        \CoreGPIO_0.xhdl1.GEN_BITS[24].APB_32.INTR_reg[24] , 
        \CoreGPIO_0.xhdl1.GEN_BITS[25].APB_32.INTR_reg[25] , 
        \CoreGPIO_0.xhdl1.GEN_BITS[26].APB_32.INTR_reg[26] , 
        \CoreGPIO_0.xhdl1.GEN_BITS[27].APB_32.INTR_reg[27] , 
        \CoreGPIO_0.xhdl1.GEN_BITS[28].APB_32.INTR_reg[28] , 
        \CoreGPIO_0.xhdl1.GEN_BITS[29].APB_32.INTR_reg[29] , 
        \CoreGPIO_0.xhdl1.GEN_BITS[30].APB_32.INTR_reg[30] , 
        \CoreGPIO_0.xhdl1.GEN_BITS[31].APB_32.INTR_reg[31] , 
        \CoreGPIO_0.xhdl1.GEN_BITS[0].REG_GEN.CONFIG_reg[0][1] , 
        \CoreGPIO_0.xhdl1.GEN_BITS[1].REG_GEN.CONFIG_reg[1][1] , 
        \CoreGPIO_0.xhdl1.GEN_BITS[2].REG_GEN.CONFIG_reg[2][1] , 
        \CoreGPIO_0.xhdl1.GEN_BITS[3].REG_GEN.CONFIG_reg[3][1] , 
        \CoreGPIO_0.xhdl1.GEN_BITS[5].REG_GEN.CONFIG_reg[5][1] , 
        \CoreGPIO_0.xhdl1.GEN_BITS[6].REG_GEN.CONFIG_reg[6][1] , 
        \CoreGPIO_0.xhdl1.GEN_BITS[0].APB_32.GPOUT_reg[0] , 
        \CoreGPIO_0.xhdl1.GEN_BITS[1].APB_32.GPOUT_reg[1] , 
        \CoreGPIO_0.xhdl1.GEN_BITS[2].APB_32.GPOUT_reg[2] , 
        \CoreGPIO_0.xhdl1.GEN_BITS[4].APB_32.GPOUT_reg[4] , 
        \CoreGPIO_0.xhdl1.GEN_BITS[5].APB_32.GPOUT_reg[5] , 
        \CoreGPIO_0.xhdl1.GEN_BITS[6].APB_32.GPOUT_reg[6] , 
        \CoreGPIO_0.xhdl1.GEN_BITS[8].APB_32.GPOUT_reg[8] , 
        \CoreGPIO_0.xhdl1.GEN_BITS[9].APB_32.GPOUT_reg[9] , 
        \CoreGPIO_0.xhdl1.GEN_BITS[10].APB_32.GPOUT_reg[10] , 
        \CoreGPIO_0.xhdl1.GEN_BITS[11].APB_32.GPOUT_reg[11] , 
        \CoreGPIO_0.xhdl1.GEN_BITS[12].APB_32.GPOUT_reg[12] , 
        \CoreGPIO_0.xhdl1.GEN_BITS[13].APB_32.GPOUT_reg[13] , 
        \CoreGPIO_0.xhdl1.GEN_BITS[14].APB_32.GPOUT_reg[14] , 
        \CoreGPIO_0.xhdl1.GEN_BITS[15].APB_32.GPOUT_reg[15] , 
        \CoreGPIO_0.xhdl1.GEN_BITS[16].APB_32.GPOUT_reg[16] , 
        \CoreGPIO_0.xhdl1.GEN_BITS[17].APB_32.GPOUT_reg[17] , 
        \CoreGPIO_0.xhdl1.GEN_BITS[18].APB_32.GPOUT_reg[18] , 
        \CoreGPIO_0.xhdl1.GEN_BITS[19].APB_32.GPOUT_reg[19] , 
        \CoreGPIO_0.xhdl1.GEN_BITS[20].APB_32.GPOUT_reg[20] , 
        \CoreGPIO_0.xhdl1.GEN_BITS[21].APB_32.GPOUT_reg[21] , 
        \CoreGPIO_0.xhdl1.GEN_BITS[22].APB_32.GPOUT_reg[22] , 
        \CoreGPIO_0.xhdl1.GEN_BITS[23].APB_32.GPOUT_reg[23] , 
        \CoreGPIO_0.xhdl1.GEN_BITS[24].APB_32.GPOUT_reg[24] , 
        \CoreGPIO_0.xhdl1.GEN_BITS[25].APB_32.GPOUT_reg[25] , 
        \CoreGPIO_0.xhdl1.GEN_BITS[26].APB_32.GPOUT_reg[26] , 
        \CoreGPIO_0.xhdl1.GEN_BITS[27].APB_32.GPOUT_reg[27] , 
        \CoreGPIO_0.xhdl1.GEN_BITS[28].APB_32.GPOUT_reg[28] , 
        \CoreGPIO_0.xhdl1.GEN_BITS[29].APB_32.GPOUT_reg[29] , 
        \CoreGPIO_0.xhdl1.GEN_BITS[30].APB_32.GPOUT_reg[30] , 
        \CoreGPIO_0.xhdl1.GEN_BITS[31].APB_32.GPOUT_reg[31] , 
        \GPIO_IN_c[6] , \GPIO_IN_c[5] , \GPIO_IN_c[4] , \GPIO_IN_c[3] , 
        \GPIO_IN_c[2] , \GPIO_IN_c[1] , \GPIO_IN_c[0] , 
        MSS_RESET_N_F2M_c, \CoreGPIO_0.N_4682 , \CoreGPIO_0.N_4706 , 
        \CoreGPIO_0.N_4738 , \CoreGPIO_0.N_4762 , \CoreGPIO_0.N_4802 , 
        \CoreGPIO_0.N_4826 , \CoreGPIO_0.N_4858 , \CoreGPIO_0.N_4882 , 
        CoreAPB3_0_APBmslave3_PSELx, \CoreGPIO_0.N_4681 , 
        \CoreGPIO_0.N_4705 , \CoreGPIO_0.N_4737 , \CoreGPIO_0.N_4761 , 
        \CoreGPIO_0.N_4801 , \CoreGPIO_0.N_4825 , \CoreGPIO_0.N_4857 , 
        \CoreGPIO_0.N_4881 , \CoreGPIO_0.N_247 , 
        \CoreAPB3_0.u_mux_p_to_b3.iPRDATA29 , 
        CoreAPB3_0_APBmslave5_PSELx, \CoreGPIO_0.N_452 , 
        \CoreGPIO_0.N_245 , \CoreGPIO_0.N_603 , \CoreGPIO_0.N_4856 , 
        \CoreGPIO_0.N_4880 , \CoreGPIO_0.N_4855 , \CoreGPIO_0.N_4879 , 
        \CoreGPIO_0.N_4854 , \CoreGPIO_0.N_4878 , \CoreGPIO_0.N_4853 , 
        \CoreGPIO_0.N_4877 , \CoreGPIO_0.N_4852 , \CoreGPIO_0.N_4876 , 
        \CoreGPIO_0.N_4851 , \CoreGPIO_0.N_4875 , \CoreGPIO_0.N_4800 , 
        \CoreGPIO_0.N_4824 , \CoreGPIO_0.N_4799 , \CoreGPIO_0.N_4823 , 
        \CoreGPIO_0.N_4798 , \CoreGPIO_0.N_4822 , \CoreGPIO_0.N_4797 , 
        \CoreGPIO_0.N_4821 , \CoreGPIO_0.N_4796 , \CoreGPIO_0.N_4820 , 
        \CoreGPIO_0.N_4795 , \CoreGPIO_0.N_4819 , \CoreGPIO_0.N_4736 , 
        \CoreGPIO_0.N_4760 , \CoreGPIO_0.N_4735 , \CoreGPIO_0.N_4759 , 
        \CoreGPIO_0.N_4734 , \CoreGPIO_0.N_4758 , \CoreGPIO_0.N_4733 , 
        \CoreGPIO_0.N_4757 , \CoreGPIO_0.N_4732 , \CoreGPIO_0.N_4756 , 
        \CoreGPIO_0.N_4731 , \CoreGPIO_0.N_4755 , \CoreGPIO_0.N_4680 , 
        \CoreGPIO_0.N_4704 , \CoreGPIO_0.N_4679 , \CoreGPIO_0.N_4703 , 
        \CoreGPIO_0.N_4678 , \CoreGPIO_0.N_4702 , \CoreGPIO_0.N_4677 , 
        \CoreGPIO_0.N_4701 , \CoreGPIO_0.N_4676 , \CoreGPIO_0.N_4700 , 
        \CoreGPIO_0.N_4675 , \CoreGPIO_0.N_4699 , 
        \CoreAPB3_0.iPSELS_2[5] , \COREAPBLSRAM_0.PRDATA4_out , 
        \xhdl1.GEN_BITS[4].REG_GEN.CONFIG_reg[4]2_0_a4_0_a2_0_RNIBB9M2 , 
        \CoreGPIO_0.PRDATA_m1_e_1 , \COREAPBLSRAM_0.wen_0 , 
        \CoreGPIO_0.N_610 , \CoreAPB3_0.CoreAPB3_N_8_i_0 , 
        \CoreAPB3_0.CoreAPB3_N_8_2_i_0 , 
        \CoreAPB3_0.CoreAPB3_N_8_3_i_0 , 
        \CoreAPB3_0.CoreAPB3_N_8_1_i_0 , 
        \CoreAPB3_0.CoreAPB3_N_8_0_i_0 , 
        \CoreAPB3_0.u_mux_p_to_b3.PREADY_0_iv_i_0 , 
        \CoreGPIO_0.PRDATA_N_3_0 , MSS_RESET_N_F2M_ibuf_net_1;
    
    INBUF MSS_RESET_N_F2M_ibuf (.PAD(MSS_RESET_N_F2M), .Y(
        MSS_RESET_N_F2M_ibuf_net_1));
    CoreAPB3_Z1 CoreAPB3_0 (.FIC_MSS_0_FIC_0_APB_MASTER_PADDR({
        \FIC_MSS_0_FIC_0_APB_MASTER_PADDR[31] , 
        \FIC_MSS_0_FIC_0_APB_MASTER_PADDR[30] , 
        \FIC_MSS_0_FIC_0_APB_MASTER_PADDR[29] , 
        \FIC_MSS_0_FIC_0_APB_MASTER_PADDR[28] }), .iPSELS_2({
        \CoreAPB3_0.iPSELS_2[5] }), .\CONFIG_reg[3] ({
        \CoreGPIO_0.xhdl1.GEN_BITS[3].REG_GEN.CONFIG_reg[3][1] }), 
        .\CONFIG_reg[5] ({
        \CoreGPIO_0.xhdl1.GEN_BITS[5].REG_GEN.CONFIG_reg[5][1] }), 
        .\CONFIG_reg[6] ({
        \CoreGPIO_0.xhdl1.GEN_BITS[6].REG_GEN.CONFIG_reg[6][1] }), 
        .\CONFIG_reg[2] ({
        \CoreGPIO_0.xhdl1.GEN_BITS[2].REG_GEN.CONFIG_reg[2][1] }), 
        .\CONFIG_reg[1] ({
        \CoreGPIO_0.xhdl1.GEN_BITS[1].REG_GEN.CONFIG_reg[1][1] }), 
        .\CONFIG_reg[0] ({
        \CoreGPIO_0.xhdl1.GEN_BITS[0].REG_GEN.CONFIG_reg[0][1] }), 
        .CoreAPB3_0_APBmslave3_PRDATA({
        \CoreAPB3_0_APBmslave3_PRDATA[7] , 
        \CoreAPB3_0_APBmslave3_PRDATA[6] , 
        \CoreAPB3_0_APBmslave3_PRDATA[5] , 
        \CoreAPB3_0_APBmslave3_PRDATA[4] , 
        \CoreAPB3_0_APBmslave3_PRDATA[3] , 
        \CoreAPB3_0_APBmslave3_PRDATA[2] , 
        \CoreAPB3_0_APBmslave3_PRDATA[1] , 
        \CoreAPB3_0_APBmslave3_PRDATA[0] }), .PRDATA_reg({
        \COREAPBLSRAM_0.PRDATA_reg[31] , 
        \COREAPBLSRAM_0.PRDATA_reg[30] , 
        \COREAPBLSRAM_0.PRDATA_reg[29] , 
        \COREAPBLSRAM_0.PRDATA_reg[28] , 
        \COREAPBLSRAM_0.PRDATA_reg[27] , 
        \COREAPBLSRAM_0.PRDATA_reg[26] , 
        \COREAPBLSRAM_0.PRDATA_reg[25] , 
        \COREAPBLSRAM_0.PRDATA_reg[24] , 
        \COREAPBLSRAM_0.PRDATA_reg[23] , 
        \COREAPBLSRAM_0.PRDATA_reg[22] , 
        \COREAPBLSRAM_0.PRDATA_reg[21] , 
        \COREAPBLSRAM_0.PRDATA_reg[20] , 
        \COREAPBLSRAM_0.PRDATA_reg[19] , 
        \COREAPBLSRAM_0.PRDATA_reg[18] , 
        \COREAPBLSRAM_0.PRDATA_reg[17] , 
        \COREAPBLSRAM_0.PRDATA_reg[16] , 
        \COREAPBLSRAM_0.PRDATA_reg[15] , 
        \COREAPBLSRAM_0.PRDATA_reg[14] , 
        \COREAPBLSRAM_0.PRDATA_reg[13] , 
        \COREAPBLSRAM_0.PRDATA_reg[12] , 
        \COREAPBLSRAM_0.PRDATA_reg[11] , 
        \COREAPBLSRAM_0.PRDATA_reg[10] , 
        \COREAPBLSRAM_0.PRDATA_reg[9] , \COREAPBLSRAM_0.PRDATA_reg[8] , 
        \COREAPBLSRAM_0.PRDATA_reg[7] , \COREAPBLSRAM_0.PRDATA_reg[6] , 
        \COREAPBLSRAM_0.PRDATA_reg[5] , \COREAPBLSRAM_0.PRDATA_reg[4] , 
        \COREAPBLSRAM_0.PRDATA_reg[3] , \COREAPBLSRAM_0.PRDATA_reg[2] , 
        \COREAPBLSRAM_0.PRDATA_reg[1] , \COREAPBLSRAM_0.PRDATA_reg[0] })
        , .lsram_width32_PRDATA({
        \COREAPBLSRAM_0.lsram_width32_PRDATA[31] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[30] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[29] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[28] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[27] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[26] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[25] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[24] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[23] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[22] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[21] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[20] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[19] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[18] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[17] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[16] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[15] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[14] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[13] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[12] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[11] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[10] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[9] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[8] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[7] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[6] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[5] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[4] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[3] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[2] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[1] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[0] }), 
        .CoreAPB3_0_APBmslave2_PADDR_5(
        \CoreAPB3_0_APBmslave2_PADDR[7] ), 
        .CoreAPB3_0_APBmslave2_PADDR_2(
        \CoreAPB3_0_APBmslave2_PADDR[4] ), 
        .CoreAPB3_0_APBmslave2_PADDR_1(
        \CoreAPB3_0_APBmslave2_PADDR[3] ), 
        .CoreAPB3_0_APBmslave2_PADDR_0(
        \CoreAPB3_0_APBmslave2_PADDR[2] ), 
        .CoreAPB3_0_APBmslave2_PADDR_3(
        \CoreAPB3_0_APBmslave2_PADDR[5] ), .gpin3_3(
        \CoreGPIO_0.xhdl1.GEN_BITS[3].gpin3[3] ), .gpin3_5(
        \CoreGPIO_0.xhdl1.GEN_BITS[5].gpin3[5] ), .gpin3_6(
        \CoreGPIO_0.xhdl1.GEN_BITS[6].gpin3[6] ), .gpin3_2(
        \CoreGPIO_0.xhdl1.GEN_BITS[2].gpin3[2] ), .gpin3_1(
        \CoreGPIO_0.xhdl1.GEN_BITS[1].gpin3[1] ), .gpin3_0(
        \CoreGPIO_0.xhdl1.GEN_BITS[0].gpin3[0] ), .GPOUT_reg_4(
        \CoreGPIO_0.xhdl1.GEN_BITS[4].APB_32.GPOUT_reg[4] ), 
        .GPOUT_reg_0(
        \CoreGPIO_0.xhdl1.GEN_BITS[0].APB_32.GPOUT_reg[0] ), 
        .GPOUT_reg_6(
        \CoreGPIO_0.xhdl1.GEN_BITS[6].APB_32.GPOUT_reg[6] ), 
        .GPOUT_reg_5(
        \CoreGPIO_0.xhdl1.GEN_BITS[5].APB_32.GPOUT_reg[5] ), 
        .GPOUT_reg_1(
        \CoreGPIO_0.xhdl1.GEN_BITS[1].APB_32.GPOUT_reg[1] ), 
        .GPOUT_reg_2(
        \CoreGPIO_0.xhdl1.GEN_BITS[2].APB_32.GPOUT_reg[2] ), 
        .GPOUT_reg_8(
        \CoreGPIO_0.xhdl1.GEN_BITS[8].APB_32.GPOUT_reg[8] ), 
        .GPOUT_reg_9(
        \CoreGPIO_0.xhdl1.GEN_BITS[9].APB_32.GPOUT_reg[9] ), 
        .GPOUT_reg_10(
        \CoreGPIO_0.xhdl1.GEN_BITS[10].APB_32.GPOUT_reg[10] ), 
        .GPOUT_reg_11(
        \CoreGPIO_0.xhdl1.GEN_BITS[11].APB_32.GPOUT_reg[11] ), 
        .GPOUT_reg_12(
        \CoreGPIO_0.xhdl1.GEN_BITS[12].APB_32.GPOUT_reg[12] ), 
        .GPOUT_reg_13(
        \CoreGPIO_0.xhdl1.GEN_BITS[13].APB_32.GPOUT_reg[13] ), 
        .GPOUT_reg_14(
        \CoreGPIO_0.xhdl1.GEN_BITS[14].APB_32.GPOUT_reg[14] ), 
        .GPOUT_reg_15(
        \CoreGPIO_0.xhdl1.GEN_BITS[15].APB_32.GPOUT_reg[15] ), 
        .GPOUT_reg_16(
        \CoreGPIO_0.xhdl1.GEN_BITS[16].APB_32.GPOUT_reg[16] ), 
        .GPOUT_reg_17(
        \CoreGPIO_0.xhdl1.GEN_BITS[17].APB_32.GPOUT_reg[17] ), 
        .GPOUT_reg_18(
        \CoreGPIO_0.xhdl1.GEN_BITS[18].APB_32.GPOUT_reg[18] ), 
        .GPOUT_reg_19(
        \CoreGPIO_0.xhdl1.GEN_BITS[19].APB_32.GPOUT_reg[19] ), 
        .GPOUT_reg_20(
        \CoreGPIO_0.xhdl1.GEN_BITS[20].APB_32.GPOUT_reg[20] ), 
        .GPOUT_reg_21(
        \CoreGPIO_0.xhdl1.GEN_BITS[21].APB_32.GPOUT_reg[21] ), 
        .GPOUT_reg_22(
        \CoreGPIO_0.xhdl1.GEN_BITS[22].APB_32.GPOUT_reg[22] ), 
        .GPOUT_reg_23(
        \CoreGPIO_0.xhdl1.GEN_BITS[23].APB_32.GPOUT_reg[23] ), 
        .GPOUT_reg_24(
        \CoreGPIO_0.xhdl1.GEN_BITS[24].APB_32.GPOUT_reg[24] ), 
        .GPOUT_reg_25(
        \CoreGPIO_0.xhdl1.GEN_BITS[25].APB_32.GPOUT_reg[25] ), 
        .GPOUT_reg_26(
        \CoreGPIO_0.xhdl1.GEN_BITS[26].APB_32.GPOUT_reg[26] ), 
        .GPOUT_reg_27(
        \CoreGPIO_0.xhdl1.GEN_BITS[27].APB_32.GPOUT_reg[27] ), 
        .GPOUT_reg_28(
        \CoreGPIO_0.xhdl1.GEN_BITS[28].APB_32.GPOUT_reg[28] ), 
        .GPOUT_reg_29(
        \CoreGPIO_0.xhdl1.GEN_BITS[29].APB_32.GPOUT_reg[29] ), 
        .GPOUT_reg_30(
        \CoreGPIO_0.xhdl1.GEN_BITS[30].APB_32.GPOUT_reg[30] ), 
        .GPOUT_reg_31(
        \CoreGPIO_0.xhdl1.GEN_BITS[31].APB_32.GPOUT_reg[31] ), 
        .INTR_reg_2(\CoreGPIO_0.xhdl1.GEN_BITS[2].APB_32.INTR_reg[2] ), 
        .INTR_reg_1(\CoreGPIO_0.xhdl1.GEN_BITS[1].APB_32.INTR_reg[1] ), 
        .INTR_reg_5(\CoreGPIO_0.xhdl1.GEN_BITS[5].APB_32.INTR_reg[5] ), 
        .INTR_reg_6(\CoreGPIO_0.xhdl1.GEN_BITS[6].APB_32.INTR_reg[6] ), 
        .INTR_reg_0(\CoreGPIO_0.xhdl1.GEN_BITS[0].APB_32.INTR_reg[0] ), 
        .INTR_reg_4(\CoreGPIO_0.xhdl1.GEN_BITS[4].APB_32.INTR_reg[4] ), 
        .INTR_reg_7(\CoreGPIO_0.xhdl1.GEN_BITS[7].APB_32.INTR_reg[7] ), 
        .INTR_reg_8(\CoreGPIO_0.xhdl1.GEN_BITS[8].APB_32.INTR_reg[8] ), 
        .INTR_reg_9(\CoreGPIO_0.xhdl1.GEN_BITS[9].APB_32.INTR_reg[9] ), 
        .INTR_reg_10(
        \CoreGPIO_0.xhdl1.GEN_BITS[10].APB_32.INTR_reg[10] ), 
        .INTR_reg_11(
        \CoreGPIO_0.xhdl1.GEN_BITS[11].APB_32.INTR_reg[11] ), 
        .INTR_reg_12(
        \CoreGPIO_0.xhdl1.GEN_BITS[12].APB_32.INTR_reg[12] ), 
        .INTR_reg_13(
        \CoreGPIO_0.xhdl1.GEN_BITS[13].APB_32.INTR_reg[13] ), 
        .INTR_reg_14(
        \CoreGPIO_0.xhdl1.GEN_BITS[14].APB_32.INTR_reg[14] ), 
        .INTR_reg_15(
        \CoreGPIO_0.xhdl1.GEN_BITS[15].APB_32.INTR_reg[15] ), 
        .INTR_reg_16(
        \CoreGPIO_0.xhdl1.GEN_BITS[16].APB_32.INTR_reg[16] ), 
        .INTR_reg_17(
        \CoreGPIO_0.xhdl1.GEN_BITS[17].APB_32.INTR_reg[17] ), 
        .INTR_reg_18(
        \CoreGPIO_0.xhdl1.GEN_BITS[18].APB_32.INTR_reg[18] ), 
        .INTR_reg_19(
        \CoreGPIO_0.xhdl1.GEN_BITS[19].APB_32.INTR_reg[19] ), 
        .INTR_reg_20(
        \CoreGPIO_0.xhdl1.GEN_BITS[20].APB_32.INTR_reg[20] ), 
        .INTR_reg_21(
        \CoreGPIO_0.xhdl1.GEN_BITS[21].APB_32.INTR_reg[21] ), 
        .INTR_reg_22(
        \CoreGPIO_0.xhdl1.GEN_BITS[22].APB_32.INTR_reg[22] ), 
        .INTR_reg_23(
        \CoreGPIO_0.xhdl1.GEN_BITS[23].APB_32.INTR_reg[23] ), 
        .INTR_reg_24(
        \CoreGPIO_0.xhdl1.GEN_BITS[24].APB_32.INTR_reg[24] ), 
        .INTR_reg_25(
        \CoreGPIO_0.xhdl1.GEN_BITS[25].APB_32.INTR_reg[25] ), 
        .INTR_reg_26(
        \CoreGPIO_0.xhdl1.GEN_BITS[26].APB_32.INTR_reg[26] ), 
        .INTR_reg_27(
        \CoreGPIO_0.xhdl1.GEN_BITS[27].APB_32.INTR_reg[27] ), 
        .INTR_reg_28(
        \CoreGPIO_0.xhdl1.GEN_BITS[28].APB_32.INTR_reg[28] ), 
        .INTR_reg_29(
        \CoreGPIO_0.xhdl1.GEN_BITS[29].APB_32.INTR_reg[29] ), 
        .INTR_reg_30(
        \CoreGPIO_0.xhdl1.GEN_BITS[30].APB_32.INTR_reg[30] ), 
        .INTR_reg_31(
        \CoreGPIO_0.xhdl1.GEN_BITS[31].APB_32.INTR_reg[31] ), 
        .FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_0(
        \FIC_MSS_0_FIC_0_APB_MASTER_PRDATA[3] ), 
        .FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_5(
        \FIC_MSS_0_FIC_0_APB_MASTER_PRDATA[8] ), 
        .FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_10(
        \FIC_MSS_0_FIC_0_APB_MASTER_PRDATA[13] ), 
        .FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_19(
        \FIC_MSS_0_FIC_0_APB_MASTER_PRDATA[22] ), 
        .FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_20(
        \FIC_MSS_0_FIC_0_APB_MASTER_PRDATA[23] ), 
        .FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_6(
        \FIC_MSS_0_FIC_0_APB_MASTER_PRDATA[9] ), 
        .FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_17(
        \FIC_MSS_0_FIC_0_APB_MASTER_PRDATA[20] ), 
        .FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_18(
        \FIC_MSS_0_FIC_0_APB_MASTER_PRDATA[21] ), 
        .FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_7(
        \FIC_MSS_0_FIC_0_APB_MASTER_PRDATA[10] ), 
        .FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_15(
        \FIC_MSS_0_FIC_0_APB_MASTER_PRDATA[18] ), 
        .FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_16(
        \FIC_MSS_0_FIC_0_APB_MASTER_PRDATA[19] ), 
        .FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_8(
        \FIC_MSS_0_FIC_0_APB_MASTER_PRDATA[11] ), 
        .FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_13(
        \FIC_MSS_0_FIC_0_APB_MASTER_PRDATA[16] ), 
        .FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_14(
        \FIC_MSS_0_FIC_0_APB_MASTER_PRDATA[17] ), 
        .FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_9(
        \FIC_MSS_0_FIC_0_APB_MASTER_PRDATA[12] ), 
        .FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_11(
        \FIC_MSS_0_FIC_0_APB_MASTER_PRDATA[14] ), 
        .FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_12(
        \FIC_MSS_0_FIC_0_APB_MASTER_PRDATA[15] ), 
        .FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_21(
        \FIC_MSS_0_FIC_0_APB_MASTER_PRDATA[24] ), 
        .FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_22(
        \FIC_MSS_0_FIC_0_APB_MASTER_PRDATA[25] ), 
        .FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_23(
        \FIC_MSS_0_FIC_0_APB_MASTER_PRDATA[26] ), 
        .FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_24(
        \FIC_MSS_0_FIC_0_APB_MASTER_PRDATA[27] ), 
        .FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_25(
        \FIC_MSS_0_FIC_0_APB_MASTER_PRDATA[28] ), 
        .FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_26(
        \FIC_MSS_0_FIC_0_APB_MASTER_PRDATA[29] ), 
        .FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_27(
        \FIC_MSS_0_FIC_0_APB_MASTER_PRDATA[30] ), 
        .FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_28(
        \FIC_MSS_0_FIC_0_APB_MASTER_PRDATA[31] ), 
        .FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_1(
        \FIC_MSS_0_FIC_0_APB_MASTER_PRDATA[4] ), 
        .FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_4(
        \FIC_MSS_0_FIC_0_APB_MASTER_PRDATA[7] ), .iPRDATA29(
        \CoreAPB3_0.u_mux_p_to_b3.iPRDATA29 ), 
        .FIC_MSS_0_FIC_0_APB_MASTER_PSELx(
        FIC_MSS_0_FIC_0_APB_MASTER_PSELx), 
        .CoreAPB3_0_APBmslave5_PSELx(CoreAPB3_0_APBmslave5_PSELx), 
        .N_245(\CoreGPIO_0.N_245 ), .N_603(\CoreGPIO_0.N_603 ), 
        .PRDATA_N_3_0(\CoreGPIO_0.PRDATA_N_3_0 ), 
        .CoreAPB3_0_APBmslave3_PSELx(CoreAPB3_0_APBmslave3_PSELx), 
        .CoreAPB3_N_8_3_i_0(\CoreAPB3_0.CoreAPB3_N_8_3_i_0 ), .N_247(
        \CoreGPIO_0.N_247 ), .CoreAPB3_N_8_2_i_0(
        \CoreAPB3_0.CoreAPB3_N_8_2_i_0 ), .CoreAPB3_N_8_1_i_0(
        \CoreAPB3_0.CoreAPB3_N_8_1_i_0 ), .CoreAPB3_N_8_i_0(
        \CoreAPB3_0.CoreAPB3_N_8_i_0 ), .N_4755(\CoreGPIO_0.N_4755 ), 
        .N_4731(\CoreGPIO_0.N_4731 ), .N_4699(\CoreGPIO_0.N_4699 ), 
        .N_4675(\CoreGPIO_0.N_4675 ), .N_4875(\CoreGPIO_0.N_4875 ), 
        .N_4851(\CoreGPIO_0.N_4851 ), .N_4819(\CoreGPIO_0.N_4819 ), 
        .N_4795(\CoreGPIO_0.N_4795 ), .N_4761(\CoreGPIO_0.N_4761 ), 
        .N_4737(\CoreGPIO_0.N_4737 ), .N_4705(\CoreGPIO_0.N_4705 ), 
        .N_4681(\CoreGPIO_0.N_4681 ), .N_4881(\CoreGPIO_0.N_4881 ), 
        .N_4857(\CoreGPIO_0.N_4857 ), .N_4825(\CoreGPIO_0.N_4825 ), 
        .N_4801(\CoreGPIO_0.N_4801 ), .N_4760(\CoreGPIO_0.N_4760 ), 
        .N_4736(\CoreGPIO_0.N_4736 ), .N_4704(\CoreGPIO_0.N_4704 ), 
        .N_4680(\CoreGPIO_0.N_4680 ), .N_4880(\CoreGPIO_0.N_4880 ), 
        .N_4856(\CoreGPIO_0.N_4856 ), .N_4824(\CoreGPIO_0.N_4824 ), 
        .N_4800(\CoreGPIO_0.N_4800 ), .N_4756(\CoreGPIO_0.N_4756 ), 
        .N_4732(\CoreGPIO_0.N_4732 ), .N_4700(\CoreGPIO_0.N_4700 ), 
        .N_4676(\CoreGPIO_0.N_4676 ), .N_4876(\CoreGPIO_0.N_4876 ), 
        .N_4852(\CoreGPIO_0.N_4852 ), .N_4820(\CoreGPIO_0.N_4820 ), 
        .N_4796(\CoreGPIO_0.N_4796 ), .N_4757(\CoreGPIO_0.N_4757 ), 
        .N_4733(\CoreGPIO_0.N_4733 ), .N_4701(\CoreGPIO_0.N_4701 ), 
        .N_4677(\CoreGPIO_0.N_4677 ), .N_4877(\CoreGPIO_0.N_4877 ), 
        .N_4853(\CoreGPIO_0.N_4853 ), .N_4821(\CoreGPIO_0.N_4821 ), 
        .N_4797(\CoreGPIO_0.N_4797 ), .N_4759(\CoreGPIO_0.N_4759 ), 
        .N_4735(\CoreGPIO_0.N_4735 ), .N_4703(\CoreGPIO_0.N_4703 ), 
        .N_4679(\CoreGPIO_0.N_4679 ), .N_4879(\CoreGPIO_0.N_4879 ), 
        .N_4855(\CoreGPIO_0.N_4855 ), .N_4823(\CoreGPIO_0.N_4823 ), 
        .N_4799(\CoreGPIO_0.N_4799 ), .N_4758(\CoreGPIO_0.N_4758 ), 
        .N_4734(\CoreGPIO_0.N_4734 ), .N_4702(\CoreGPIO_0.N_4702 ), 
        .N_4678(\CoreGPIO_0.N_4678 ), .N_4878(\CoreGPIO_0.N_4878 ), 
        .N_4854(\CoreGPIO_0.N_4854 ), .N_4822(\CoreGPIO_0.N_4822 ), 
        .N_4798(\CoreGPIO_0.N_4798 ), .CoreAPB3_0_APBmslave2_PENABLE(
        CoreAPB3_0_APBmslave2_PENABLE), .CoreAPB3_0_APBmslave2_PWRITE(
        CoreAPB3_0_APBmslave2_PWRITE), .N_610(\CoreGPIO_0.N_610 ), 
        .PRDATA4_out(\COREAPBLSRAM_0.PRDATA4_out ), 
        .CoreAPB3_N_8_0_i_0(\CoreAPB3_0.CoreAPB3_N_8_0_i_0 ), .N_4762(
        \CoreGPIO_0.N_4762 ), .N_4738(\CoreGPIO_0.N_4738 ), .N_4706(
        \CoreGPIO_0.N_4706 ), .N_4682(\CoreGPIO_0.N_4682 ), .N_4882(
        \CoreGPIO_0.N_4882 ), .N_4858(\CoreGPIO_0.N_4858 ), .N_4826(
        \CoreGPIO_0.N_4826 ), .N_4802(\CoreGPIO_0.N_4802 ), 
        .PRDATA_m1_e_1(\CoreGPIO_0.PRDATA_m1_e_1 ), 
        .CoreAPB3_0_APBmslave3_PREADY(CoreAPB3_0_APBmslave3_PREADY), 
        .CoreAPB3_0_APBmslave2_PREADY(CoreAPB3_0_APBmslave2_PREADY), 
        .PREADY_0_iv_i_0(\CoreAPB3_0.u_mux_p_to_b3.PREADY_0_iv_i_0 ), 
        .\CONFIG_reg[4]2_0_a4_0_a2_0_RNIBB9M2 (
        \xhdl1.GEN_BITS[4].REG_GEN.CONFIG_reg[4]2_0_a4_0_a2_0_RNIBB9M2 )
        , .N_452(\CoreGPIO_0.N_452 ));
    INBUF \GPIO_IN_ibuf[2]  (.PAD(GPIO_IN[2]), .Y(\GPIO_IN_c[2] ));
    OUTBUF \GPIO_OUT_obuf[6]  (.D(\GPIO_OUT_net_2[6] ), .PAD(
        GPIO_OUT[6]));
    OUTBUF \GPIO_OUT_obuf[5]  (.D(\GPIO_OUT_net_2[5] ), .PAD(
        GPIO_OUT[5]));
    OUTBUF \GPIO_OUT_obuf[0]  (.D(\GPIO_OUT_net_2[0] ), .PAD(
        GPIO_OUT[0]));
    INBUF \GPIO_IN_ibuf[1]  (.PAD(GPIO_IN[1]), .Y(\GPIO_IN_c[1] ));
    INBUF \GPIO_IN_ibuf[0]  (.PAD(GPIO_IN[0]), .Y(\GPIO_IN_c[0] ));
    GND GND (.Y(GND_net_1));
    FIC_OSC_0_OSC OSC_0 (
        .OSC_0_RCOSC_25_50MHZ_CCC_OUT_RCOSC_25_50MHZ_CCC(
        OSC_0_RCOSC_25_50MHZ_CCC_OUT_RCOSC_25_50MHZ_CCC));
    INBUF \GPIO_IN_ibuf[6]  (.PAD(GPIO_IN[6]), .Y(\GPIO_IN_c[6] ));
    CLKINT MSS_RESET_N_F2M_ibuf_RNIBBDD (.A(MSS_RESET_N_F2M_ibuf_net_1)
        , .Y(MSS_RESET_N_F2M_c));
    OUTBUF \GPIO_OUT_obuf[2]  (.D(\GPIO_OUT_net_2[2] ), .PAD(
        GPIO_OUT[2]));
    OUTBUF \GPIO_OUT_obuf[1]  (.D(\GPIO_OUT_net_2[1] ), .PAD(
        GPIO_OUT[1]));
    OUTBUF \GPIO_OUT_obuf[4]  (.D(\GPIO_OUT_net_2[4] ), .PAD(
        GPIO_OUT[4]));
    INBUF \GPIO_IN_ibuf[4]  (.PAD(GPIO_IN[4]), .Y(\GPIO_IN_c[4] ));
    FIC_FCCC_0_FCCC FCCC_0 (.FCCC_0_GL1(FCCC_0_GL1), .FCCC_0_LOCK(
        FCCC_0_LOCK), .OSC_0_RCOSC_25_50MHZ_CCC_OUT_RCOSC_25_50MHZ_CCC(
        OSC_0_RCOSC_25_50MHZ_CCC_OUT_RCOSC_25_50MHZ_CCC));
    reg_apb_wrp reg_apb_wrp_0 (.CoreAPB3_0_APBmslave3_PRDATA({
        \CoreAPB3_0_APBmslave3_PRDATA[7] , 
        \CoreAPB3_0_APBmslave3_PRDATA[6] , 
        \CoreAPB3_0_APBmslave3_PRDATA[5] , 
        \CoreAPB3_0_APBmslave3_PRDATA[4] , 
        \CoreAPB3_0_APBmslave3_PRDATA[3] , 
        \CoreAPB3_0_APBmslave3_PRDATA[2] , 
        \CoreAPB3_0_APBmslave3_PRDATA[1] , 
        \CoreAPB3_0_APBmslave3_PRDATA[0] }), 
        .CoreAPB3_0_APBmslave2_PWDATA({
        \CoreAPB3_0_APBmslave2_PWDATA[7] , 
        \CoreAPB3_0_APBmslave2_PWDATA[6] , 
        \CoreAPB3_0_APBmslave2_PWDATA[5] , 
        \CoreAPB3_0_APBmslave2_PWDATA[4] , 
        \CoreAPB3_0_APBmslave2_PWDATA[3] , 
        \CoreAPB3_0_APBmslave2_PWDATA[2] , 
        \CoreAPB3_0_APBmslave2_PWDATA[1] , 
        \CoreAPB3_0_APBmslave2_PWDATA[0] }), 
        .CoreAPB3_0_APBmslave2_PADDR({\CoreAPB3_0_APBmslave2_PADDR[3] , 
        \CoreAPB3_0_APBmslave2_PADDR[2] , 
        \CoreAPB3_0_APBmslave2_PADDR[1] , 
        \CoreAPB3_0_APBmslave2_PADDR[0] }), 
        .CoreAPB3_0_APBmslave3_PREADY(CoreAPB3_0_APBmslave3_PREADY), 
        .MSS_RESET_N_F2M_c(MSS_RESET_N_F2M_c), .FCCC_0_GL1(FCCC_0_GL1), 
        .CoreAPB3_0_APBmslave2_PWRITE(CoreAPB3_0_APBmslave2_PWRITE), 
        .CoreAPB3_0_APBmslave3_PSELx(CoreAPB3_0_APBmslave3_PSELx));
    OUTBUF \GPIO_OUT_obuf[3]  (.D(\GPIO_OUT_net_2[3] ), .PAD(
        GPIO_OUT[3]));
    FIC_MSS FIC_MSS_0 (.CoreAPB3_0_APBmslave2_PADDR({
        \CoreAPB3_0_APBmslave2_PADDR[8] , 
        \CoreAPB3_0_APBmslave2_PADDR[7] , 
        \CoreAPB3_0_APBmslave2_PADDR[6] , 
        \CoreAPB3_0_APBmslave2_PADDR[5] , 
        \CoreAPB3_0_APBmslave2_PADDR[4] , 
        \CoreAPB3_0_APBmslave2_PADDR[3] , 
        \CoreAPB3_0_APBmslave2_PADDR[2] , 
        \CoreAPB3_0_APBmslave2_PADDR[1] , 
        \CoreAPB3_0_APBmslave2_PADDR[0] }), 
        .FIC_MSS_0_FIC_0_APB_MASTER_PADDR({
        \FIC_MSS_0_FIC_0_APB_MASTER_PADDR[31] , 
        \FIC_MSS_0_FIC_0_APB_MASTER_PADDR[30] , 
        \FIC_MSS_0_FIC_0_APB_MASTER_PADDR[29] , 
        \FIC_MSS_0_FIC_0_APB_MASTER_PADDR[28] }), 
        .CoreAPB3_0_APBmslave2_PWDATA({
        \CoreAPB3_0_APBmslave2_PWDATA[31] , 
        \CoreAPB3_0_APBmslave2_PWDATA[30] , 
        \CoreAPB3_0_APBmslave2_PWDATA[29] , 
        \CoreAPB3_0_APBmslave2_PWDATA[28] , 
        \CoreAPB3_0_APBmslave2_PWDATA[27] , 
        \CoreAPB3_0_APBmslave2_PWDATA[26] , 
        \CoreAPB3_0_APBmslave2_PWDATA[25] , 
        \CoreAPB3_0_APBmslave2_PWDATA[24] , 
        \CoreAPB3_0_APBmslave2_PWDATA[23] , 
        \CoreAPB3_0_APBmslave2_PWDATA[22] , 
        \CoreAPB3_0_APBmslave2_PWDATA[21] , 
        \CoreAPB3_0_APBmslave2_PWDATA[20] , 
        \CoreAPB3_0_APBmslave2_PWDATA[19] , 
        \CoreAPB3_0_APBmslave2_PWDATA[18] , 
        \CoreAPB3_0_APBmslave2_PWDATA[17] , 
        \CoreAPB3_0_APBmslave2_PWDATA[16] , 
        \CoreAPB3_0_APBmslave2_PWDATA[15] , 
        \CoreAPB3_0_APBmslave2_PWDATA[14] , 
        \CoreAPB3_0_APBmslave2_PWDATA[13] , 
        \CoreAPB3_0_APBmslave2_PWDATA[12] , 
        \CoreAPB3_0_APBmslave2_PWDATA[11] , 
        \CoreAPB3_0_APBmslave2_PWDATA[10] , 
        \CoreAPB3_0_APBmslave2_PWDATA[9] , 
        \CoreAPB3_0_APBmslave2_PWDATA[8] , 
        \CoreAPB3_0_APBmslave2_PWDATA[7] , 
        \CoreAPB3_0_APBmslave2_PWDATA[6] , 
        \CoreAPB3_0_APBmslave2_PWDATA[5] , 
        \CoreAPB3_0_APBmslave2_PWDATA[4] , 
        \CoreAPB3_0_APBmslave2_PWDATA[3] , 
        \CoreAPB3_0_APBmslave2_PWDATA[2] , 
        \CoreAPB3_0_APBmslave2_PWDATA[1] , 
        \CoreAPB3_0_APBmslave2_PWDATA[0] }), 
        .FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_0(
        \FIC_MSS_0_FIC_0_APB_MASTER_PRDATA[3] ), 
        .FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_1(
        \FIC_MSS_0_FIC_0_APB_MASTER_PRDATA[4] ), 
        .FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_4(
        \FIC_MSS_0_FIC_0_APB_MASTER_PRDATA[7] ), 
        .FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_5(
        \FIC_MSS_0_FIC_0_APB_MASTER_PRDATA[8] ), 
        .FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_6(
        \FIC_MSS_0_FIC_0_APB_MASTER_PRDATA[9] ), 
        .FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_7(
        \FIC_MSS_0_FIC_0_APB_MASTER_PRDATA[10] ), 
        .FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_8(
        \FIC_MSS_0_FIC_0_APB_MASTER_PRDATA[11] ), 
        .FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_9(
        \FIC_MSS_0_FIC_0_APB_MASTER_PRDATA[12] ), 
        .FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_10(
        \FIC_MSS_0_FIC_0_APB_MASTER_PRDATA[13] ), 
        .FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_11(
        \FIC_MSS_0_FIC_0_APB_MASTER_PRDATA[14] ), 
        .FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_12(
        \FIC_MSS_0_FIC_0_APB_MASTER_PRDATA[15] ), 
        .FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_13(
        \FIC_MSS_0_FIC_0_APB_MASTER_PRDATA[16] ), 
        .FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_14(
        \FIC_MSS_0_FIC_0_APB_MASTER_PRDATA[17] ), 
        .FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_15(
        \FIC_MSS_0_FIC_0_APB_MASTER_PRDATA[18] ), 
        .FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_16(
        \FIC_MSS_0_FIC_0_APB_MASTER_PRDATA[19] ), 
        .FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_17(
        \FIC_MSS_0_FIC_0_APB_MASTER_PRDATA[20] ), 
        .FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_18(
        \FIC_MSS_0_FIC_0_APB_MASTER_PRDATA[21] ), 
        .FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_19(
        \FIC_MSS_0_FIC_0_APB_MASTER_PRDATA[22] ), 
        .FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_20(
        \FIC_MSS_0_FIC_0_APB_MASTER_PRDATA[23] ), 
        .FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_21(
        \FIC_MSS_0_FIC_0_APB_MASTER_PRDATA[24] ), 
        .FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_22(
        \FIC_MSS_0_FIC_0_APB_MASTER_PRDATA[25] ), 
        .FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_23(
        \FIC_MSS_0_FIC_0_APB_MASTER_PRDATA[26] ), 
        .FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_24(
        \FIC_MSS_0_FIC_0_APB_MASTER_PRDATA[27] ), 
        .FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_25(
        \FIC_MSS_0_FIC_0_APB_MASTER_PRDATA[28] ), 
        .FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_26(
        \FIC_MSS_0_FIC_0_APB_MASTER_PRDATA[29] ), 
        .FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_27(
        \FIC_MSS_0_FIC_0_APB_MASTER_PRDATA[30] ), 
        .FIC_MSS_0_FIC_0_APB_MASTER_PRDATA_28(
        \FIC_MSS_0_FIC_0_APB_MASTER_PRDATA[31] ), .MMUART_0_TXD(
        MMUART_0_TXD), .MMUART_0_RXD(MMUART_0_RXD), 
        .CoreAPB3_0_APBmslave2_PENABLE(CoreAPB3_0_APBmslave2_PENABLE), 
        .FIC_MSS_0_FIC_0_APB_MASTER_PSELx(
        FIC_MSS_0_FIC_0_APB_MASTER_PSELx), 
        .CoreAPB3_0_APBmslave2_PWRITE(CoreAPB3_0_APBmslave2_PWRITE), 
        .CoreAPB3_N_8_i_0(\CoreAPB3_0.CoreAPB3_N_8_i_0 ), 
        .CoreAPB3_N_8_2_i_0(\CoreAPB3_0.CoreAPB3_N_8_2_i_0 ), 
        .CoreAPB3_N_8_3_i_0(\CoreAPB3_0.CoreAPB3_N_8_3_i_0 ), 
        .CoreAPB3_N_8_1_i_0(\CoreAPB3_0.CoreAPB3_N_8_1_i_0 ), 
        .CoreAPB3_N_8_0_i_0(\CoreAPB3_0.CoreAPB3_N_8_0_i_0 ), 
        .PREADY_0_iv_i_0(\CoreAPB3_0.u_mux_p_to_b3.PREADY_0_iv_i_0 ), 
        .FCCC_0_LOCK(FCCC_0_LOCK), .MSS_RESET_N_F2M_c(
        MSS_RESET_N_F2M_c), .FCCC_0_GL1(FCCC_0_GL1));
    VCC VCC (.Y(VCC_net_1));
    INBUF \GPIO_IN_ibuf[3]  (.PAD(GPIO_IN[3]), .Y(\GPIO_IN_c[3] ));
    INBUF \GPIO_IN_ibuf[5]  (.PAD(GPIO_IN[5]), .Y(\GPIO_IN_c[5] ));
    CoreGPIO_Z3 CoreGPIO_0 (.CoreAPB3_0_APBmslave2_PWDATA({
        \CoreAPB3_0_APBmslave2_PWDATA[31] , 
        \CoreAPB3_0_APBmslave2_PWDATA[30] , 
        \CoreAPB3_0_APBmslave2_PWDATA[29] , 
        \CoreAPB3_0_APBmslave2_PWDATA[28] , 
        \CoreAPB3_0_APBmslave2_PWDATA[27] , 
        \CoreAPB3_0_APBmslave2_PWDATA[26] , 
        \CoreAPB3_0_APBmslave2_PWDATA[25] , 
        \CoreAPB3_0_APBmslave2_PWDATA[24] , 
        \CoreAPB3_0_APBmslave2_PWDATA[23] , 
        \CoreAPB3_0_APBmslave2_PWDATA[22] , 
        \CoreAPB3_0_APBmslave2_PWDATA[21] , 
        \CoreAPB3_0_APBmslave2_PWDATA[20] , 
        \CoreAPB3_0_APBmslave2_PWDATA[19] , 
        \CoreAPB3_0_APBmslave2_PWDATA[18] , 
        \CoreAPB3_0_APBmslave2_PWDATA[17] , 
        \CoreAPB3_0_APBmslave2_PWDATA[16] , 
        \CoreAPB3_0_APBmslave2_PWDATA[15] , 
        \CoreAPB3_0_APBmslave2_PWDATA[14] , 
        \CoreAPB3_0_APBmslave2_PWDATA[13] , 
        \CoreAPB3_0_APBmslave2_PWDATA[12] , 
        \CoreAPB3_0_APBmslave2_PWDATA[11] , 
        \CoreAPB3_0_APBmslave2_PWDATA[10] , 
        \CoreAPB3_0_APBmslave2_PWDATA[9] , 
        \CoreAPB3_0_APBmslave2_PWDATA[8] , 
        \CoreAPB3_0_APBmslave2_PWDATA[7] , 
        \CoreAPB3_0_APBmslave2_PWDATA[6] , 
        \CoreAPB3_0_APBmslave2_PWDATA[5] , 
        \CoreAPB3_0_APBmslave2_PWDATA[4] , 
        \CoreAPB3_0_APBmslave2_PWDATA[3] , 
        \CoreAPB3_0_APBmslave2_PWDATA[2] , 
        \CoreAPB3_0_APBmslave2_PWDATA[1] , 
        \CoreAPB3_0_APBmslave2_PWDATA[0] }), .GPIO_IN_c({
        \GPIO_IN_c[6] , \GPIO_IN_c[5] , \GPIO_IN_c[4] , \GPIO_IN_c[3] , 
        \GPIO_IN_c[2] , \GPIO_IN_c[1] , \GPIO_IN_c[0] }), 
        .GPIO_OUT_net_2({\GPIO_OUT_net_2[6] , \GPIO_OUT_net_2[5] , 
        \GPIO_OUT_net_2[4] , \GPIO_OUT_net_2[3] , \GPIO_OUT_net_2[2] , 
        \GPIO_OUT_net_2[1] , \GPIO_OUT_net_2[0] }), 
        .CoreAPB3_0_APBmslave2_PADDR({\CoreAPB3_0_APBmslave2_PADDR[7] , 
        \CoreAPB3_0_APBmslave2_PADDR[6] , 
        \CoreAPB3_0_APBmslave2_PADDR[5] , 
        \CoreAPB3_0_APBmslave2_PADDR[4] , 
        \CoreAPB3_0_APBmslave2_PADDR[3] , 
        \CoreAPB3_0_APBmslave2_PADDR[2] , 
        \CoreAPB3_0_APBmslave2_PADDR[1] , 
        \CoreAPB3_0_APBmslave2_PADDR[0] }), .iPSELS_2({
        \CoreAPB3_0.iPSELS_2[5] }), .GPOUT_reg_31(
        \CoreGPIO_0.xhdl1.GEN_BITS[31].APB_32.GPOUT_reg[31] ), 
        .GPOUT_reg_30(
        \CoreGPIO_0.xhdl1.GEN_BITS[30].APB_32.GPOUT_reg[30] ), 
        .GPOUT_reg_29(
        \CoreGPIO_0.xhdl1.GEN_BITS[29].APB_32.GPOUT_reg[29] ), 
        .GPOUT_reg_28(
        \CoreGPIO_0.xhdl1.GEN_BITS[28].APB_32.GPOUT_reg[28] ), 
        .GPOUT_reg_27(
        \CoreGPIO_0.xhdl1.GEN_BITS[27].APB_32.GPOUT_reg[27] ), 
        .GPOUT_reg_26(
        \CoreGPIO_0.xhdl1.GEN_BITS[26].APB_32.GPOUT_reg[26] ), 
        .GPOUT_reg_25(
        \CoreGPIO_0.xhdl1.GEN_BITS[25].APB_32.GPOUT_reg[25] ), 
        .GPOUT_reg_24(
        \CoreGPIO_0.xhdl1.GEN_BITS[24].APB_32.GPOUT_reg[24] ), 
        .GPOUT_reg_23(
        \CoreGPIO_0.xhdl1.GEN_BITS[23].APB_32.GPOUT_reg[23] ), 
        .GPOUT_reg_22(
        \CoreGPIO_0.xhdl1.GEN_BITS[22].APB_32.GPOUT_reg[22] ), 
        .GPOUT_reg_21(
        \CoreGPIO_0.xhdl1.GEN_BITS[21].APB_32.GPOUT_reg[21] ), 
        .GPOUT_reg_20(
        \CoreGPIO_0.xhdl1.GEN_BITS[20].APB_32.GPOUT_reg[20] ), 
        .GPOUT_reg_19(
        \CoreGPIO_0.xhdl1.GEN_BITS[19].APB_32.GPOUT_reg[19] ), 
        .GPOUT_reg_18(
        \CoreGPIO_0.xhdl1.GEN_BITS[18].APB_32.GPOUT_reg[18] ), 
        .GPOUT_reg_17(
        \CoreGPIO_0.xhdl1.GEN_BITS[17].APB_32.GPOUT_reg[17] ), 
        .GPOUT_reg_16(
        \CoreGPIO_0.xhdl1.GEN_BITS[16].APB_32.GPOUT_reg[16] ), 
        .GPOUT_reg_15(
        \CoreGPIO_0.xhdl1.GEN_BITS[15].APB_32.GPOUT_reg[15] ), 
        .GPOUT_reg_14(
        \CoreGPIO_0.xhdl1.GEN_BITS[14].APB_32.GPOUT_reg[14] ), 
        .GPOUT_reg_13(
        \CoreGPIO_0.xhdl1.GEN_BITS[13].APB_32.GPOUT_reg[13] ), 
        .GPOUT_reg_12(
        \CoreGPIO_0.xhdl1.GEN_BITS[12].APB_32.GPOUT_reg[12] ), 
        .GPOUT_reg_11(
        \CoreGPIO_0.xhdl1.GEN_BITS[11].APB_32.GPOUT_reg[11] ), 
        .GPOUT_reg_10(
        \CoreGPIO_0.xhdl1.GEN_BITS[10].APB_32.GPOUT_reg[10] ), 
        .GPOUT_reg_9(
        \CoreGPIO_0.xhdl1.GEN_BITS[9].APB_32.GPOUT_reg[9] ), 
        .GPOUT_reg_8(
        \CoreGPIO_0.xhdl1.GEN_BITS[8].APB_32.GPOUT_reg[8] ), 
        .GPOUT_reg_6(
        \CoreGPIO_0.xhdl1.GEN_BITS[6].APB_32.GPOUT_reg[6] ), 
        .GPOUT_reg_5(
        \CoreGPIO_0.xhdl1.GEN_BITS[5].APB_32.GPOUT_reg[5] ), 
        .GPOUT_reg_4(
        \CoreGPIO_0.xhdl1.GEN_BITS[4].APB_32.GPOUT_reg[4] ), 
        .GPOUT_reg_2(
        \CoreGPIO_0.xhdl1.GEN_BITS[2].APB_32.GPOUT_reg[2] ), 
        .GPOUT_reg_1(
        \CoreGPIO_0.xhdl1.GEN_BITS[1].APB_32.GPOUT_reg[1] ), 
        .GPOUT_reg_0(
        \CoreGPIO_0.xhdl1.GEN_BITS[0].APB_32.GPOUT_reg[0] ), 
        .\CONFIG_reg[6]_1 (
        \CoreGPIO_0.xhdl1.GEN_BITS[6].REG_GEN.CONFIG_reg[6][1] ), 
        .\CONFIG_reg[5]_1 (
        \CoreGPIO_0.xhdl1.GEN_BITS[5].REG_GEN.CONFIG_reg[5][1] ), 
        .\CONFIG_reg[3]_1 (
        \CoreGPIO_0.xhdl1.GEN_BITS[3].REG_GEN.CONFIG_reg[3][1] ), 
        .\CONFIG_reg[2]_1 (
        \CoreGPIO_0.xhdl1.GEN_BITS[2].REG_GEN.CONFIG_reg[2][1] ), 
        .\CONFIG_reg[1]_1 (
        \CoreGPIO_0.xhdl1.GEN_BITS[1].REG_GEN.CONFIG_reg[1][1] ), 
        .\CONFIG_reg[0]_1 (
        \CoreGPIO_0.xhdl1.GEN_BITS[0].REG_GEN.CONFIG_reg[0][1] ), 
        .INTR_reg_23(
        \CoreGPIO_0.xhdl1.GEN_BITS[23].APB_32.INTR_reg[23] ), 
        .INTR_reg_24(
        \CoreGPIO_0.xhdl1.GEN_BITS[24].APB_32.INTR_reg[24] ), 
        .INTR_reg_25(
        \CoreGPIO_0.xhdl1.GEN_BITS[25].APB_32.INTR_reg[25] ), 
        .INTR_reg_26(
        \CoreGPIO_0.xhdl1.GEN_BITS[26].APB_32.INTR_reg[26] ), 
        .INTR_reg_27(
        \CoreGPIO_0.xhdl1.GEN_BITS[27].APB_32.INTR_reg[27] ), 
        .INTR_reg_28(
        \CoreGPIO_0.xhdl1.GEN_BITS[28].APB_32.INTR_reg[28] ), 
        .INTR_reg_29(
        \CoreGPIO_0.xhdl1.GEN_BITS[29].APB_32.INTR_reg[29] ), 
        .INTR_reg_30(
        \CoreGPIO_0.xhdl1.GEN_BITS[30].APB_32.INTR_reg[30] ), 
        .INTR_reg_31(
        \CoreGPIO_0.xhdl1.GEN_BITS[31].APB_32.INTR_reg[31] ), 
        .INTR_reg_8(\CoreGPIO_0.xhdl1.GEN_BITS[8].APB_32.INTR_reg[8] ), 
        .INTR_reg_9(\CoreGPIO_0.xhdl1.GEN_BITS[9].APB_32.INTR_reg[9] ), 
        .INTR_reg_10(
        \CoreGPIO_0.xhdl1.GEN_BITS[10].APB_32.INTR_reg[10] ), 
        .INTR_reg_11(
        \CoreGPIO_0.xhdl1.GEN_BITS[11].APB_32.INTR_reg[11] ), 
        .INTR_reg_12(
        \CoreGPIO_0.xhdl1.GEN_BITS[12].APB_32.INTR_reg[12] ), 
        .INTR_reg_13(
        \CoreGPIO_0.xhdl1.GEN_BITS[13].APB_32.INTR_reg[13] ), 
        .INTR_reg_14(
        \CoreGPIO_0.xhdl1.GEN_BITS[14].APB_32.INTR_reg[14] ), 
        .INTR_reg_15(
        \CoreGPIO_0.xhdl1.GEN_BITS[15].APB_32.INTR_reg[15] ), 
        .INTR_reg_16(
        \CoreGPIO_0.xhdl1.GEN_BITS[16].APB_32.INTR_reg[16] ), 
        .INTR_reg_17(
        \CoreGPIO_0.xhdl1.GEN_BITS[17].APB_32.INTR_reg[17] ), 
        .INTR_reg_18(
        \CoreGPIO_0.xhdl1.GEN_BITS[18].APB_32.INTR_reg[18] ), 
        .INTR_reg_19(
        \CoreGPIO_0.xhdl1.GEN_BITS[19].APB_32.INTR_reg[19] ), 
        .INTR_reg_20(
        \CoreGPIO_0.xhdl1.GEN_BITS[20].APB_32.INTR_reg[20] ), 
        .INTR_reg_21(
        \CoreGPIO_0.xhdl1.GEN_BITS[21].APB_32.INTR_reg[21] ), 
        .INTR_reg_22(
        \CoreGPIO_0.xhdl1.GEN_BITS[22].APB_32.INTR_reg[22] ), 
        .INTR_reg_0(\CoreGPIO_0.xhdl1.GEN_BITS[0].APB_32.INTR_reg[0] ), 
        .INTR_reg_1(\CoreGPIO_0.xhdl1.GEN_BITS[1].APB_32.INTR_reg[1] ), 
        .INTR_reg_2(\CoreGPIO_0.xhdl1.GEN_BITS[2].APB_32.INTR_reg[2] ), 
        .INTR_reg_4(\CoreGPIO_0.xhdl1.GEN_BITS[4].APB_32.INTR_reg[4] ), 
        .INTR_reg_5(\CoreGPIO_0.xhdl1.GEN_BITS[5].APB_32.INTR_reg[5] ), 
        .INTR_reg_6(\CoreGPIO_0.xhdl1.GEN_BITS[6].APB_32.INTR_reg[6] ), 
        .INTR_reg_7(\CoreGPIO_0.xhdl1.GEN_BITS[7].APB_32.INTR_reg[7] ), 
        .gpin3_5(\CoreGPIO_0.xhdl1.GEN_BITS[5].gpin3[5] ), .gpin3_6(
        \CoreGPIO_0.xhdl1.GEN_BITS[6].gpin3[6] ), .gpin3_0(
        \CoreGPIO_0.xhdl1.GEN_BITS[0].gpin3[0] ), .gpin3_1(
        \CoreGPIO_0.xhdl1.GEN_BITS[1].gpin3[1] ), .gpin3_2(
        \CoreGPIO_0.xhdl1.GEN_BITS[2].gpin3[2] ), .gpin3_3(
        \CoreGPIO_0.xhdl1.GEN_BITS[3].gpin3[3] ), 
        .FIC_MSS_0_FIC_0_APB_MASTER_PADDR_2(
        \FIC_MSS_0_FIC_0_APB_MASTER_PADDR[31] ), 
        .FIC_MSS_0_FIC_0_APB_MASTER_PADDR_0(
        \FIC_MSS_0_FIC_0_APB_MASTER_PADDR[29] ), .MSS_RESET_N_F2M_c(
        MSS_RESET_N_F2M_c), .FCCC_0_GL1(FCCC_0_GL1), .PRDATA_N_3_0(
        \CoreGPIO_0.PRDATA_N_3_0 ), .N_4801(\CoreGPIO_0.N_4801 ), 
        .N_4762(\CoreGPIO_0.N_4762 ), .N_4706(\CoreGPIO_0.N_4706 ), 
        .N_4682(\CoreGPIO_0.N_4682 ), .N_4852(\CoreGPIO_0.N_4852 ), 
        .N_4857(\CoreGPIO_0.N_4857 ), .N_4825(\CoreGPIO_0.N_4825 ), 
        .N_4736(\CoreGPIO_0.N_4736 ), .N_4705(\CoreGPIO_0.N_4705 ), 
        .N_4858(\CoreGPIO_0.N_4858 ), .N_4819(\CoreGPIO_0.N_4819 ), 
        .N_4851(\CoreGPIO_0.N_4851 ), .N_4761(\CoreGPIO_0.N_4761 ), 
        .N_4802(\CoreGPIO_0.N_4802 ), .N_4738(\CoreGPIO_0.N_4738 ), 
        .N_4880(\CoreGPIO_0.N_4880 ), .N_4879(\CoreGPIO_0.N_4879 ), 
        .N_4877(\CoreGPIO_0.N_4877 ), .N_4735(\CoreGPIO_0.N_4735 ), 
        .N_4881(\CoreGPIO_0.N_4881 ), .N_4798(\CoreGPIO_0.N_4798 ), 
        .N_4797(\CoreGPIO_0.N_4797 ), .N_4796(\CoreGPIO_0.N_4796 ), 
        .N_4758(\CoreGPIO_0.N_4758 ), .N_4757(\CoreGPIO_0.N_4757 ), 
        .N_4756(\CoreGPIO_0.N_4756 ), .N_4878(\CoreGPIO_0.N_4878 ), 
        .N_4823(\CoreGPIO_0.N_4823 ), .N_4876(\CoreGPIO_0.N_4876 ), 
        .N_4734(\CoreGPIO_0.N_4734 ), .N_4733(\CoreGPIO_0.N_4733 ), 
        .N_4732(\CoreGPIO_0.N_4732 ), .N_4731(\CoreGPIO_0.N_4731 ), 
        .N_4676(\CoreGPIO_0.N_4676 ), .N_4675(\CoreGPIO_0.N_4675 ), 
        .N_4795(\CoreGPIO_0.N_4795 ), .N_4826(\CoreGPIO_0.N_4826 ), 
        .N_4701(\CoreGPIO_0.N_4701 ), .N_4882(\CoreGPIO_0.N_4882 ), 
        .N_4755(\CoreGPIO_0.N_4755 ), .N_4702(\CoreGPIO_0.N_4702 ), 
        .N_4853(\CoreGPIO_0.N_4853 ), .N_4677(\CoreGPIO_0.N_4677 ), 
        .N_4820(\CoreGPIO_0.N_4820 ), .N_4854(\CoreGPIO_0.N_4854 ), 
        .N_4759(\CoreGPIO_0.N_4759 ), .N_4678(\CoreGPIO_0.N_4678 ), 
        .N_4760(\CoreGPIO_0.N_4760 ), .N_4681(\CoreGPIO_0.N_4681 ), 
        .N_4824(\CoreGPIO_0.N_4824 ), .N_4703(\CoreGPIO_0.N_4703 ), 
        .N_4737(\CoreGPIO_0.N_4737 ), .N_4704(\CoreGPIO_0.N_4704 ), 
        .N_4679(\CoreGPIO_0.N_4679 ), .N_4699(\CoreGPIO_0.N_4699 ), 
        .N_4799(\CoreGPIO_0.N_4799 ), .N_4855(\CoreGPIO_0.N_4855 ), 
        .N_4680(\CoreGPIO_0.N_4680 ), .N_4875(\CoreGPIO_0.N_4875 ), 
        .N_4800(\CoreGPIO_0.N_4800 ), .N_4822(\CoreGPIO_0.N_4822 ), 
        .N_4821(\CoreGPIO_0.N_4821 ), .N_4700(\CoreGPIO_0.N_4700 ), 
        .N_4856(\CoreGPIO_0.N_4856 ), .N_610(\CoreGPIO_0.N_610 ), 
        .N_603(\CoreGPIO_0.N_603 ), .PRDATA_m1_e_1(
        \CoreGPIO_0.PRDATA_m1_e_1 ), .N_245(\CoreGPIO_0.N_245 ), 
        .N_452(\CoreGPIO_0.N_452 ), .N_247(\CoreGPIO_0.N_247 ), 
        .CoreAPB3_0_APBmslave5_PSELx(CoreAPB3_0_APBmslave5_PSELx), 
        .wen_0(\COREAPBLSRAM_0.wen_0 ), 
        .\CONFIG_reg[4]2_0_a4_0_a2_0_RNIBB9M2 (
        \xhdl1.GEN_BITS[4].REG_GEN.CONFIG_reg[4]2_0_a4_0_a2_0_RNIBB9M2 )
        );
    FIC_COREAPBLSRAM_0_COREAPBLSRAM_Z2 COREAPBLSRAM_0 (.PRDATA_reg({
        \COREAPBLSRAM_0.PRDATA_reg[31] , 
        \COREAPBLSRAM_0.PRDATA_reg[30] , 
        \COREAPBLSRAM_0.PRDATA_reg[29] , 
        \COREAPBLSRAM_0.PRDATA_reg[28] , 
        \COREAPBLSRAM_0.PRDATA_reg[27] , 
        \COREAPBLSRAM_0.PRDATA_reg[26] , 
        \COREAPBLSRAM_0.PRDATA_reg[25] , 
        \COREAPBLSRAM_0.PRDATA_reg[24] , 
        \COREAPBLSRAM_0.PRDATA_reg[23] , 
        \COREAPBLSRAM_0.PRDATA_reg[22] , 
        \COREAPBLSRAM_0.PRDATA_reg[21] , 
        \COREAPBLSRAM_0.PRDATA_reg[20] , 
        \COREAPBLSRAM_0.PRDATA_reg[19] , 
        \COREAPBLSRAM_0.PRDATA_reg[18] , 
        \COREAPBLSRAM_0.PRDATA_reg[17] , 
        \COREAPBLSRAM_0.PRDATA_reg[16] , 
        \COREAPBLSRAM_0.PRDATA_reg[15] , 
        \COREAPBLSRAM_0.PRDATA_reg[14] , 
        \COREAPBLSRAM_0.PRDATA_reg[13] , 
        \COREAPBLSRAM_0.PRDATA_reg[12] , 
        \COREAPBLSRAM_0.PRDATA_reg[11] , 
        \COREAPBLSRAM_0.PRDATA_reg[10] , 
        \COREAPBLSRAM_0.PRDATA_reg[9] , \COREAPBLSRAM_0.PRDATA_reg[8] , 
        \COREAPBLSRAM_0.PRDATA_reg[7] , \COREAPBLSRAM_0.PRDATA_reg[6] , 
        \COREAPBLSRAM_0.PRDATA_reg[5] , \COREAPBLSRAM_0.PRDATA_reg[4] , 
        \COREAPBLSRAM_0.PRDATA_reg[3] , \COREAPBLSRAM_0.PRDATA_reg[2] , 
        \COREAPBLSRAM_0.PRDATA_reg[1] , \COREAPBLSRAM_0.PRDATA_reg[0] })
        , .lsram_width32_PRDATA({
        \COREAPBLSRAM_0.lsram_width32_PRDATA[31] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[30] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[29] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[28] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[27] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[26] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[25] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[24] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[23] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[22] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[21] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[20] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[19] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[18] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[17] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[16] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[15] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[14] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[13] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[12] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[11] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[10] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[9] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[8] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[7] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[6] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[5] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[4] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[3] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[2] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[1] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[0] }), 
        .CoreAPB3_0_APBmslave2_PADDR({\CoreAPB3_0_APBmslave2_PADDR[8] , 
        \CoreAPB3_0_APBmslave2_PADDR[7] , 
        \CoreAPB3_0_APBmslave2_PADDR[6] , 
        \CoreAPB3_0_APBmslave2_PADDR[5] , 
        \CoreAPB3_0_APBmslave2_PADDR[4] , 
        \CoreAPB3_0_APBmslave2_PADDR[3] , 
        \CoreAPB3_0_APBmslave2_PADDR[2] , 
        \CoreAPB3_0_APBmslave2_PADDR[1] , 
        \CoreAPB3_0_APBmslave2_PADDR[0] }), 
        .CoreAPB3_0_APBmslave2_PWDATA({
        \CoreAPB3_0_APBmslave2_PWDATA[31] , 
        \CoreAPB3_0_APBmslave2_PWDATA[30] , 
        \CoreAPB3_0_APBmslave2_PWDATA[29] , 
        \CoreAPB3_0_APBmslave2_PWDATA[28] , 
        \CoreAPB3_0_APBmslave2_PWDATA[27] , 
        \CoreAPB3_0_APBmslave2_PWDATA[26] , 
        \CoreAPB3_0_APBmslave2_PWDATA[25] , 
        \CoreAPB3_0_APBmslave2_PWDATA[24] , 
        \CoreAPB3_0_APBmslave2_PWDATA[23] , 
        \CoreAPB3_0_APBmslave2_PWDATA[22] , 
        \CoreAPB3_0_APBmslave2_PWDATA[21] , 
        \CoreAPB3_0_APBmslave2_PWDATA[20] , 
        \CoreAPB3_0_APBmslave2_PWDATA[19] , 
        \CoreAPB3_0_APBmslave2_PWDATA[18] , 
        \CoreAPB3_0_APBmslave2_PWDATA[17] , 
        \CoreAPB3_0_APBmslave2_PWDATA[16] , 
        \CoreAPB3_0_APBmslave2_PWDATA[15] , 
        \CoreAPB3_0_APBmslave2_PWDATA[14] , 
        \CoreAPB3_0_APBmslave2_PWDATA[13] , 
        \CoreAPB3_0_APBmslave2_PWDATA[12] , 
        \CoreAPB3_0_APBmslave2_PWDATA[11] , 
        \CoreAPB3_0_APBmslave2_PWDATA[10] , 
        \CoreAPB3_0_APBmslave2_PWDATA[9] , 
        \CoreAPB3_0_APBmslave2_PWDATA[8] , 
        \CoreAPB3_0_APBmslave2_PWDATA[7] , 
        \CoreAPB3_0_APBmslave2_PWDATA[6] , 
        \CoreAPB3_0_APBmslave2_PWDATA[5] , 
        \CoreAPB3_0_APBmslave2_PWDATA[4] , 
        \CoreAPB3_0_APBmslave2_PWDATA[3] , 
        \CoreAPB3_0_APBmslave2_PWDATA[2] , 
        \CoreAPB3_0_APBmslave2_PWDATA[1] , 
        \CoreAPB3_0_APBmslave2_PWDATA[0] }), .MSS_RESET_N_F2M_c(
        MSS_RESET_N_F2M_c), .FCCC_0_GL1(FCCC_0_GL1), 
        .CoreAPB3_0_APBmslave2_PREADY(CoreAPB3_0_APBmslave2_PREADY), 
        .CoreAPB3_0_APBmslave2_PENABLE(CoreAPB3_0_APBmslave2_PENABLE), 
        .CoreAPB3_0_APBmslave2_PWRITE(CoreAPB3_0_APBmslave2_PWRITE), 
        .wen_0(\COREAPBLSRAM_0.wen_0 ), .PRDATA4_out(
        \COREAPBLSRAM_0.PRDATA4_out ), .iPRDATA29(
        \CoreAPB3_0.u_mux_p_to_b3.iPRDATA29 ));
    
endmodule
