`timescale 1 ns/100 ps
// Version: 
// File used only for Simulation


module sdf_IOPAD_BI(
       PAD,
       D,
       E,
       Y
    );
inout  PAD;
input  D;
input  E;
output Y;

    wire NET_IOUT_VDD, NET_IOUT_IN, NET_OIN_VDD, NET_EIN_VDD;
    
    IOPAD_BI_VDDI U_VCCI (.OIN_VDD(NET_OIN_VDD), .EIN_VDD(NET_EIN_VDD), 
        .IOUT_VDD(NET_IOUT_VDD), .PAD_P(PAD));
    IOPAD_DELAY U_DELAY (.IOUT_IN(NET_IOUT_IN), .IOUT_P(Y));
    IOPAD_VDD U_VCCA (.OIN_P(D), .EIN_P(E), .IOUT_VDD(NET_IOUT_VDD), 
        .OIN_VDD(NET_OIN_VDD), .EIN_VDD(NET_EIN_VDD), .IOUT_IN(
        NET_IOUT_IN));
    
endmodule


module sdf_IOPAD_TRI(
       PAD,
       D,
       E
    );
output PAD;
input  D;
input  E;

    wire NET_OIN_VDD, NET_EIN_VDD;
    
    IOPAD_TRI_VDDI U_VCCI (.OIN_VDD(NET_OIN_VDD), .EIN_VDD(NET_EIN_VDD)
        , .PAD_P(PAD));
    IOPAD_VDD U_VCCA (.OIN_P(D), .EIN_P(E), .IOUT_VDD(), .OIN_VDD(
        NET_OIN_VDD), .EIN_VDD(NET_EIN_VDD), .IOUT_IN());
    
endmodule


module sdf_IOPADP_TRI(
       PAD_P,
       OIN_P,
       EIN_P
    );
output PAD_P;
input  OIN_P;
input  EIN_P;

    wire NET_OIN_VDD, NET_EIN_VDD;
    
    IOPADP_TRI_VDDI U_VCCI (.OIN_VDD(NET_OIN_VDD), .EIN_VDD(
        NET_EIN_VDD), .PAD_P(PAD_P));
    IOPADP_VDD U_VCCA (.OIN_P(OIN_P), .EIN_P(EIN_P), .IOUT_VDD(), 
        .OIN_VDD(NET_OIN_VDD), .EIN_VDD(NET_EIN_VDD), .IOUT_IN());
    
endmodule


module sdf_IOPADN_BI(
       PAD_P,
       OIN_P,
       EIN_P,
       N2POUT_P
    );
inout  PAD_P;
input  OIN_P;
input  EIN_P;
output N2POUT_P;

    wire NET_IOUT_VDD, NET_IOUT_IN, NET_OIN_VDD, NET_EIN_VDD;
    
    IOPADN_BI_VDDI U_VCCI (.OIN_VDD(NET_OIN_VDD), .EIN_VDD(NET_EIN_VDD)
        , .IOUT_VDD(NET_IOUT_VDD), .PAD_P(PAD_P));
    IOPADN_DELAY U_DELAY (.IOUT_IN(NET_IOUT_IN), .N2POUT_P(N2POUT_P));
    IOPADN_VDD U_VCCA (.OIN_P(OIN_P), .EIN_P(EIN_P), .IOUT_VDD(
        NET_IOUT_VDD), .OIN_VDD(NET_OIN_VDD), .EIN_VDD(NET_EIN_VDD), 
        .IOUT_IN(NET_IOUT_IN));
    
endmodule


module sdf_IOPAD_IN(
       PAD,
       Y
    );
input  PAD;
output Y;

    wire NET_IOUT_VDD, NET_IOUT_IN, ADLIB_GND;
    wire GND_power_net1;
    assign ADLIB_GND = GND_power_net1;
    
    IOPAD_IN_VDDI U_VCCI (.PAD_P(PAD), .IOUT_VDD(NET_IOUT_VDD));
    IOPAD_DELAY U_DELAY (.IOUT_IN(NET_IOUT_IN), .IOUT_P(Y));
    IOPAD_VDD U_VCCA (.OIN_P(ADLIB_GND), .EIN_P(ADLIB_GND), .IOUT_VDD(
        NET_IOUT_VDD), .OIN_VDD(), .EIN_VDD(), .IOUT_IN(NET_IOUT_IN));
    GND GND_power_inst1 (.Y(GND_power_net1));
    
endmodule


module sdf_IOPADP_BI(
       PAD_P,
       N2PIN_P,
       OIN_P,
       EIN_P,
       IOUT_P
    );
inout  PAD_P;
input  N2PIN_P;
input  OIN_P;
input  EIN_P;
output IOUT_P;

    wire NET_IOUT_VDD, NET_IOUT_IN, NET_OIN_VDD, NET_EIN_VDD;
    
    IOPADP_BI_VDDI U_VCCI (.OIN_VDD(NET_OIN_VDD), .EIN_VDD(NET_EIN_VDD)
        , .N2PIN_P(N2PIN_P), .IOUT_VDD(NET_IOUT_VDD), .PAD_P(PAD_P));
    IOPADP_DELAY U_DELAY (.IOUT_IN(NET_IOUT_IN), .IOUT_P(IOUT_P));
    IOPADP_VDD U_VCCA (.OIN_P(OIN_P), .EIN_P(EIN_P), .IOUT_VDD(
        NET_IOUT_VDD), .OIN_VDD(NET_OIN_VDD), .EIN_VDD(NET_EIN_VDD), 
        .IOUT_IN(NET_IOUT_IN));
    
endmodule


module sdf_IOPADN_TRI(
       PAD_P,
       OIN_P,
       EIN_P
    );
output PAD_P;
input  OIN_P;
input  EIN_P;

    wire NET_OIN_VDD, NET_EIN_VDD;
    
    IOPADN_TRI_VDDI U_VCCI (.OIN_VDD(NET_OIN_VDD), .EIN_VDD(
        NET_EIN_VDD), .PAD_P(PAD_P));
    IOPADN_VDD U_VCCA (.OIN_P(OIN_P), .EIN_P(EIN_P), .IOUT_VDD(), 
        .OIN_VDD(NET_OIN_VDD), .EIN_VDD(NET_EIN_VDD), .IOUT_IN());
    
endmodule


module FIC(
       GPIO_IN,
       GPIO_OUT,
       MDDR_ADDR,
       MDDR_BA,
       MDDR_DM_RDQS,
       MDDR_DQ,
       MDDR_DQS,
       MDDR_DQS_N,
       MDDR_DQS_TMATCH_0_IN,
       MMUART_0_RXD,
       MSS_RESET_N_F2M,
       MDDR_CAS_N,
       MDDR_CKE,
       MDDR_CLK,
       MDDR_CLK_N,
       MDDR_CS_N,
       MDDR_DQS_TMATCH_0_OUT,
       MDDR_ODT,
       MDDR_RAS_N,
       MDDR_RESET_N,
       MDDR_WE_N,
       MMUART_0_TXD
    );
input  [0:6] GPIO_IN;
output [0:6] GPIO_OUT;
output [15:0] MDDR_ADDR;
output [2:0] MDDR_BA;
inout  [1:0] MDDR_DM_RDQS;
inout  [15:0] MDDR_DQ;
inout  [1:0] MDDR_DQS;
inout  [1:0] MDDR_DQS_N;
input  MDDR_DQS_TMATCH_0_IN;
input  MMUART_0_RXD;
input  MSS_RESET_N_F2M;
output MDDR_CAS_N;
output MDDR_CKE;
output MDDR_CLK;
output MDDR_CLK_N;
output MDDR_CS_N;
output MDDR_DQS_TMATCH_0_OUT;
output MDDR_ODT;
output MDDR_RAS_N;
output MDDR_RESET_N;
output MDDR_WE_N;
output MMUART_0_TXD;

    wire \GPIO_OUT_net_2[6] , \GPIO_OUT_net_2[5] , \GPIO_OUT_net_2[4] , 
        \GPIO_OUT_net_2[3] , \GPIO_OUT_net_2[2] , \GPIO_OUT_net_2[1] , 
        \GPIO_OUT_net_2[0] , \CoreAPB3_0_APBmslave3_PADDR[0] , 
        \CoreAPB3_0_APBmslave3_PADDR[1] , 
        \CoreAPB3_0_APBmslave3_PADDR[2] , 
        \CoreAPB3_0_APBmslave3_PADDR[3] , 
        \CoreAPB3_0_APBmslave3_PADDR[4] , 
        \CoreAPB3_0_APBmslave3_PADDR[5] , 
        \CoreAPB3_0_APBmslave3_PADDR[6] , 
        \CoreAPB3_0_APBmslave3_PADDR[7] , 
        \FIC_MSS_0_FIC_0_APB_MASTER_PADDR[28] , 
        \FIC_MSS_0_FIC_0_APB_MASTER_PADDR[29] , 
        \FIC_MSS_0_FIC_0_APB_MASTER_PADDR[30] , 
        \FIC_MSS_0_FIC_0_APB_MASTER_PADDR[31] , 
        CoreAPB3_0_APBmslave3_PWRITE, CoreAPB3_0_APBmslave3_PENABLE, 
        FIC_MSS_0_FIC_0_APB_MASTER_PSELx, 
        \CoreAPB3_0_APBmslave3_PWDATA[0] , 
        \CoreAPB3_0_APBmslave3_PWDATA[1] , 
        \CoreAPB3_0_APBmslave3_PWDATA[2] , 
        \CoreAPB3_0_APBmslave3_PWDATA[3] , 
        \CoreAPB3_0_APBmslave3_PWDATA[4] , 
        \CoreAPB3_0_APBmslave3_PWDATA[5] , 
        \CoreAPB3_0_APBmslave3_PWDATA[6] , 
        \CoreAPB3_0_APBmslave3_PWDATA[7] , 
        \CoreAPB3_0_APBmslave3_PWDATA[8] , 
        \CoreAPB3_0_APBmslave3_PWDATA[9] , 
        \CoreAPB3_0_APBmslave3_PWDATA[10] , 
        \CoreAPB3_0_APBmslave3_PWDATA[11] , 
        \CoreAPB3_0_APBmslave3_PWDATA[12] , 
        \CoreAPB3_0_APBmslave3_PWDATA[13] , 
        \CoreAPB3_0_APBmslave3_PWDATA[14] , 
        \CoreAPB3_0_APBmslave3_PWDATA[15] , 
        \CoreAPB3_0_APBmslave3_PWDATA[16] , 
        \CoreAPB3_0_APBmslave3_PWDATA[17] , 
        \CoreAPB3_0_APBmslave3_PWDATA[18] , 
        \CoreAPB3_0_APBmslave3_PWDATA[19] , 
        \CoreAPB3_0_APBmslave3_PWDATA[20] , 
        \CoreAPB3_0_APBmslave3_PWDATA[21] , 
        \CoreAPB3_0_APBmslave3_PWDATA[22] , 
        \CoreAPB3_0_APBmslave3_PWDATA[23] , 
        \CoreAPB3_0_APBmslave3_PWDATA[24] , 
        \CoreAPB3_0_APBmslave3_PWDATA[25] , 
        \CoreAPB3_0_APBmslave3_PWDATA[26] , 
        \CoreAPB3_0_APBmslave3_PWDATA[27] , 
        \CoreAPB3_0_APBmslave3_PWDATA[28] , 
        \CoreAPB3_0_APBmslave3_PWDATA[29] , 
        \CoreAPB3_0_APBmslave3_PWDATA[30] , 
        \CoreAPB3_0_APBmslave3_PWDATA[31] , 
        \FIC_MSS_0_FIC_0_APB_MASTER_PRDATA[7] , 
        \FIC_MSS_0_FIC_0_APB_MASTER_PRDATA[8] , 
        \FIC_MSS_0_FIC_0_APB_MASTER_PRDATA[9] , 
        \FIC_MSS_0_FIC_0_APB_MASTER_PRDATA[10] , 
        \FIC_MSS_0_FIC_0_APB_MASTER_PRDATA[11] , 
        \FIC_MSS_0_FIC_0_APB_MASTER_PRDATA[12] , 
        \FIC_MSS_0_FIC_0_APB_MASTER_PRDATA[13] , 
        \FIC_MSS_0_FIC_0_APB_MASTER_PRDATA[14] , 
        \FIC_MSS_0_FIC_0_APB_MASTER_PRDATA[15] , 
        \FIC_MSS_0_FIC_0_APB_MASTER_PRDATA[16] , 
        \FIC_MSS_0_FIC_0_APB_MASTER_PRDATA[17] , 
        \FIC_MSS_0_FIC_0_APB_MASTER_PRDATA[18] , 
        \FIC_MSS_0_FIC_0_APB_MASTER_PRDATA[19] , 
        \FIC_MSS_0_FIC_0_APB_MASTER_PRDATA[20] , 
        \FIC_MSS_0_FIC_0_APB_MASTER_PRDATA[21] , 
        \FIC_MSS_0_FIC_0_APB_MASTER_PRDATA[22] , 
        \FIC_MSS_0_FIC_0_APB_MASTER_PRDATA[23] , 
        \FIC_MSS_0_FIC_0_APB_MASTER_PRDATA[24] , 
        \FIC_MSS_0_FIC_0_APB_MASTER_PRDATA[25] , 
        \FIC_MSS_0_FIC_0_APB_MASTER_PRDATA[26] , 
        \FIC_MSS_0_FIC_0_APB_MASTER_PRDATA[27] , 
        \FIC_MSS_0_FIC_0_APB_MASTER_PRDATA[28] , 
        \FIC_MSS_0_FIC_0_APB_MASTER_PRDATA[29] , 
        \FIC_MSS_0_FIC_0_APB_MASTER_PRDATA[30] , 
        \FIC_MSS_0_FIC_0_APB_MASTER_PRDATA[31] , 
        \CoreAPB3_0_APBmslave3_PRDATA[0] , 
        \CoreAPB3_0_APBmslave3_PRDATA[1] , 
        \CoreAPB3_0_APBmslave3_PRDATA[2] , 
        \CoreAPB3_0_APBmslave3_PRDATA[3] , 
        \CoreAPB3_0_APBmslave3_PRDATA[4] , 
        \CoreAPB3_0_APBmslave3_PRDATA[5] , 
        \CoreAPB3_0_APBmslave3_PRDATA[6] , 
        \CoreAPB3_0_APBmslave3_PRDATA[7] , 
        CoreAPB3_0_APBmslave3_PREADY, \FCCC_0/GL1_INST/U0_YNn , 
        OSC_0_RCOSC_25_50MHZ_CCC_OUT_RCOSC_25_50MHZ_CCC, FCCC_0_LOCK, 
        CoreAPB3_0_APBmslave5_PSELx, CoreAPB3_0_APBmslave3_PSELx, 
        \CoreAPB3_0.iPSELS_raw23 , 
        \CoreGPIO_0.xhdl1.GEN_BITS[0].gpin3[0] , 
        \CoreGPIO_0.xhdl1.GEN_BITS[1].gpin3[1] , 
        \CoreGPIO_0.xhdl1.GEN_BITS[2].gpin3[2] , 
        \CoreGPIO_0.xhdl1.GEN_BITS[3].gpin3[3] , 
        \CoreGPIO_0.xhdl1.GEN_BITS[4].gpin3[4] , 
        \CoreGPIO_0.xhdl1.GEN_BITS[5].gpin3[5] , 
        \CoreGPIO_0.xhdl1.GEN_BITS[6].gpin3[6] , 
        \CoreGPIO_0.xhdl1.GEN_BITS[1].APB_32.INTR_reg[1] , 
        \CoreGPIO_0.xhdl1.GEN_BITS[3].APB_32.INTR_reg[3] , 
        \CoreGPIO_0.xhdl1.GEN_BITS[4].APB_32.INTR_reg[4] , 
        \CoreGPIO_0.xhdl1.GEN_BITS[5].APB_32.INTR_reg[5] , 
        \CoreGPIO_0.xhdl1.GEN_BITS[6].APB_32.INTR_reg[6] , 
        \CoreGPIO_0.xhdl1.GEN_BITS[10].APB_32.INTR_reg[10] , 
        \CoreGPIO_0.xhdl1.GEN_BITS[18].APB_32.INTR_reg[18] , 
        \CoreGPIO_0.xhdl1.GEN_BITS[26].APB_32.INTR_reg[26] , 
        \CoreGPIO_0.xhdl1.GEN_BITS[0].REG_GEN.CONFIG_reg[0][1] , 
        \CoreGPIO_0.xhdl1.GEN_BITS[1].REG_GEN.CONFIG_reg[1][1] , 
        \CoreGPIO_0.xhdl1.GEN_BITS[2].REG_GEN.CONFIG_reg[2][1] , 
        \CoreGPIO_0.xhdl1.GEN_BITS[3].REG_GEN.CONFIG_reg[3][1] , 
        \CoreGPIO_0.xhdl1.GEN_BITS[4].REG_GEN.CONFIG_reg[4][1] , 
        \CoreGPIO_0.xhdl1.GEN_BITS[5].REG_GEN.CONFIG_reg[5][1] , 
        \CoreGPIO_0.xhdl1.GEN_BITS[6].REG_GEN.CONFIG_reg[6][1] , 
        \CoreGPIO_0.xhdl1.GEN_BITS[1].APB_32.GPOUT_reg[1] , 
        \CoreGPIO_0.xhdl1.GEN_BITS[4].APB_32.GPOUT_reg[4] , 
        \CoreGPIO_0.xhdl1.GEN_BITS[5].APB_32.GPOUT_reg[5] , 
        \CoreGPIO_0.xhdl1.GEN_BITS[6].APB_32.GPOUT_reg[6] , 
        \CoreGPIO_0.xhdl1.GEN_BITS[8].APB_32.GPOUT_reg[8] , 
        \CoreGPIO_0.xhdl1.GEN_BITS[9].APB_32.GPOUT_reg[9] , 
        \CoreGPIO_0.xhdl1.GEN_BITS[11].APB_32.GPOUT_reg[11] , 
        \CoreGPIO_0.xhdl1.GEN_BITS[12].APB_32.GPOUT_reg[12] , 
        \CoreGPIO_0.xhdl1.GEN_BITS[13].APB_32.GPOUT_reg[13] , 
        \CoreGPIO_0.xhdl1.GEN_BITS[14].APB_32.GPOUT_reg[14] , 
        \CoreGPIO_0.xhdl1.GEN_BITS[15].APB_32.GPOUT_reg[15] , 
        \CoreGPIO_0.xhdl1.GEN_BITS[16].APB_32.GPOUT_reg[16] , 
        \CoreGPIO_0.xhdl1.GEN_BITS[17].APB_32.GPOUT_reg[17] , 
        \CoreGPIO_0.xhdl1.GEN_BITS[19].APB_32.GPOUT_reg[19] , 
        \CoreGPIO_0.xhdl1.GEN_BITS[20].APB_32.GPOUT_reg[20] , 
        \CoreGPIO_0.xhdl1.GEN_BITS[21].APB_32.GPOUT_reg[21] , 
        \CoreGPIO_0.xhdl1.GEN_BITS[22].APB_32.GPOUT_reg[22] , 
        \CoreGPIO_0.xhdl1.GEN_BITS[23].APB_32.GPOUT_reg[23] , 
        \CoreGPIO_0.xhdl1.GEN_BITS[24].APB_32.GPOUT_reg[24] , 
        \CoreGPIO_0.xhdl1.GEN_BITS[25].APB_32.GPOUT_reg[25] , 
        \CoreGPIO_0.xhdl1.GEN_BITS[27].APB_32.GPOUT_reg[27] , 
        \CoreGPIO_0.xhdl1.GEN_BITS[28].APB_32.GPOUT_reg[28] , 
        \CoreGPIO_0.xhdl1.GEN_BITS[29].APB_32.GPOUT_reg[29] , 
        \CoreGPIO_0.xhdl1.GEN_BITS[30].APB_32.GPOUT_reg[30] , 
        \CoreGPIO_0.xhdl1.GEN_BITS[31].APB_32.GPOUT_reg[31] , 
        \CoreGPIO_0.xhdl1.GEN_BITS[0].APB_32.GPOUT_reg9 , 
        \CoreGPIO_0.RDATA_32.un12_PRDATA_o , 
        \CoreGPIO_0.CONFIG_reg_o_2[7] , \CoreGPIO_0.N_246 , 
        \CoreGPIO_0.N_247 , \CoreGPIO_0.N_496 , \CoreGPIO_0.N_524 , 
        \CoreGPIO_0.N_526 , \CoreGPIO_0.N_528 , \CoreGPIO_0.N_530 , 
        \CoreGPIO_0.N_532 , \CoreGPIO_0.N_533 , \CoreGPIO_0.N_536 , 
        \CoreGPIO_0.N_538 , \CoreGPIO_0.N_540 , \CoreGPIO_0.N_542 , 
        \CoreGPIO_0.N_544 , \CoreGPIO_0.N_546 , \CoreGPIO_0.N_548 , 
        \CoreGPIO_0.N_549 , \CoreGPIO_0.N_552 , \CoreGPIO_0.N_554 , 
        \CoreGPIO_0.N_556 , \CoreGPIO_0.N_558 , \CoreGPIO_0.N_560 , 
        \CoreGPIO_0.N_562 , \CoreGPIO_0.N_564 , \CoreGPIO_0.N_565 , 
        \CoreGPIO_0.N_568 , \CoreGPIO_0.N_570 , \GPIO_IN_c[6] , 
        \GPIO_IN_c[5] , \GPIO_IN_c[4] , \GPIO_IN_c[3] , \GPIO_IN_c[2] , 
        \GPIO_IN_c[1] , \GPIO_IN_c[0] , 
        \CoreGPIO_0.RDATA_32.un12_PRDATA_o_0_o2_1 , 
        \CoreGPIO_0.PRDATA_iv_0_0_1[2] , 
        \CoreGPIO_0.PRDATA_iv_0_0_1[0] , 
        \CoreGPIO_0.PRDATA_0_iv_0_0_0[7] , \CONFIG_reg_o_2_31_am[3] , 
        \CONFIG_reg_o_2_31_bm[3] , \CoreGPIO_0.PRDATA_iv_0_0_0_0[0] , 
        \CoreGPIO_0.PRDATA_iv_0_0_1[5] , 
        \CoreGPIO_0.PRDATA_iv_0_0_0_0[1] , 
        \CoreGPIO_0.PRDATA_iv_0_0_1[4] , 
        \CoreGPIO_0.PRDATA_iv_0_0_0_0[6] , 
        \CoreGPIO_0.PRDATA_iv_0_0_0_0[2] , 
        \xhdl1.GEN_BITS[0].APB_32.un5_PRDATA_o_0_a2_0_o2_x , 
        MSS_RESET_N_F2M_ibuf, \CoreAPB3_0/iPSELS_1[5] , 
        \CoreAPB3_0/u_mux_p_to_b3/PRDATA_0_iv_1[7]_net_1 , 
        \FCCC_0/GL1_net , VCC, GND, \reg_apb_wrp_0/N_64_i_0 , 
        \reg_apb_wrp_0/N_44_i_0 , \reg_apb_wrp_0/wr_enable_net_1 , 
        \reg_apb_wrp_0/N_70 , \reg_apb_wrp_0/N_45_i_0 , 
        \reg_apb_wrp_0/rd_enable_net_1 , \reg_apb_wrp_0/N_76 , 
        \reg_apb_wrp_0/fsm[0]_net_1 , \reg_apb_wrp_0/fsm_ns[0] , 
        \reg_apb_wrp_0/fsm[1]_net_1 , \reg_apb_wrp_0/fsm_ns[1] , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_122_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_26_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_10_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_80_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_28_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_12_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_81_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_57_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_112_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_104_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_16_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_88_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_97_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_72_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_7_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_125_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_29_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_13_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_14_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_82_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_59_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_113_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_105_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_17_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_89_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_98_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_73_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_5_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_127_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_31_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_15_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_2_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_124_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_84_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_56_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_114_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_106_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_18_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_90_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_99_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_74_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_64_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_49_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_33_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_40_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_4_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_126_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_30_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_61_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_115_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_107_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_19_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_91_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_96_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_75_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_66_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_51_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_35_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_42_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_6_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_48_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_32_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_43_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_116_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_108_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_20_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_92_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_101_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_76_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_68_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_53_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_37_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_44_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_65_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_50_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_34_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_41_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_85_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_109_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_21_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_93_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_102_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_77_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_69_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_54_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_39_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_46_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_67_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_52_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_36_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_47_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_86_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_58_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_22_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_94_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_103_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_78_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_70_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_3_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_121_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_25_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_9_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_83_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_38_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_45_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_87_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_62_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_117_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_95_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_100_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_79_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_71_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_1_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_123_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_27_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_11_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_55_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_120_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_24_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_8_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_63_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_118_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_110_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_60_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_119_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_111_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_23_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/temp_data[0]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/N_5_i_0 , 
        \reg_apb_wrp_0/reg16x8_0/temp_data[1]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/N_7_i_0 , 
        \reg_apb_wrp_0/reg16x8_0/temp_data[2]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/N_9_i_0 , 
        \reg_apb_wrp_0/reg16x8_0/temp_data[3]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/N_11_i_0 , 
        \reg_apb_wrp_0/reg16x8_0/temp_data[4]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/N_19_i_0 , 
        \reg_apb_wrp_0/reg16x8_0/temp_data[5]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/N_25_i_0 , 
        \reg_apb_wrp_0/reg16x8_0/temp_data[6]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/N_52_i_0 , 
        \reg_apb_wrp_0/reg16x8_0/temp_data[7]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/N_86_i_0 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_23_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_231_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_12_rs[7] , 
        \reg_apb_wrp_0/reg16x8_0/mem_12_[7]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_231_i , 
        \reg_apb_wrp_0/reg16x8_0/mem_12__1_sqmuxa , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_111_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_239_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_13_rs[7] , 
        \reg_apb_wrp_0/reg16x8_0/mem_13_[7]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_239_i , 
        \reg_apb_wrp_0/reg16x8_0/mem_13__1_sqmuxa , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_119_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_247_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_14_rs[7] , 
        \reg_apb_wrp_0/reg16x8_0/mem_14_[7]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_247_i , 
        \reg_apb_wrp_0/reg16x8_0/mem_14__1_sqmuxa , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_60_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_252_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_15_rs[7] , 
        \reg_apb_wrp_0/reg16x8_0/mem_15_[7]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_252_i , 
        \reg_apb_wrp_0/reg16x8_0/mem_15__1_sqmuxa , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_110_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_238_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_13_rs[6] , 
        \reg_apb_wrp_0/reg16x8_0/mem_13_[6]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_238_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_118_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_246_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_14_rs[6] , 
        \reg_apb_wrp_0/reg16x8_0/mem_14_[6]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_246_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_63_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_255_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_15_rs[6] , 
        \reg_apb_wrp_0/reg16x8_0/mem_15_[6]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_255_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_8_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_135_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_0_rs[7] , 
        \reg_apb_wrp_0/reg16x8_0/mem_0_[7]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_135_i , 
        \reg_apb_wrp_0/reg16x8_0/mem_0__1_sqmuxa , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_24_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_143_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_1_rs[7] , 
        \reg_apb_wrp_0/reg16x8_0/mem_1_[7]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_143_i , 
        \reg_apb_wrp_0/reg16x8_0/mem_1__1_sqmuxa , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_120_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_151_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_2_rs[7] , 
        \reg_apb_wrp_0/reg16x8_0/mem_2_[7]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_151_i , 
        \reg_apb_wrp_0/reg16x8_0/mem_2__1_sqmuxa , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_55_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_160_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_3_rs[7] , 
        \reg_apb_wrp_0/reg16x8_0/mem_3_[7]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_160_i , 
        \reg_apb_wrp_0/reg16x8_0/mem_3__1_sqmuxa , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_11_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_170_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_4_rs[7] , 
        \reg_apb_wrp_0/reg16x8_0/mem_4_[7]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_170_i , 
        \reg_apb_wrp_0/reg16x8_0/mem_4__1_sqmuxa , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_27_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_186_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_5_rs[7] , 
        \reg_apb_wrp_0/reg16x8_0/mem_5_[7]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_186_i , 
        \reg_apb_wrp_0/reg16x8_0/mem_5__1_sqmuxa , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_123_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_202_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_6_rs[7] , 
        \reg_apb_wrp_0/reg16x8_0/mem_6_[7]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_202_i , 
        \reg_apb_wrp_0/reg16x8_0/mem_6__1_sqmuxa , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_1_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_217_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_7_rs[7] , 
        \reg_apb_wrp_0/reg16x8_0/mem_7_[7]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_217_i , 
        \reg_apb_wrp_0/reg16x8_0/mem_7__1_sqmuxa , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_71_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_173_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_8_rs[7] , 
        \reg_apb_wrp_0/reg16x8_0/mem_8_[7]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_173_i , 
        \reg_apb_wrp_0/reg16x8_0/mem_8__1_sqmuxa , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_79_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_189_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_9_rs[7] , 
        \reg_apb_wrp_0/reg16x8_0/mem_9_[7]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_189_i , 
        \reg_apb_wrp_0/reg16x8_0/mem_9__1_sqmuxa , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_100_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_205_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_10_rs[7] , 
        \reg_apb_wrp_0/reg16x8_0/mem_10_[7]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_205_i , 
        \reg_apb_wrp_0/reg16x8_0/mem_10__1_sqmuxa , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_95_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_220_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_11_rs[7] , 
        \reg_apb_wrp_0/reg16x8_0/mem_11_[7]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_220_i , 
        \reg_apb_wrp_0/reg16x8_0/mem_11__1_sqmuxa , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_117_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_245_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_14_rs[5] , 
        \reg_apb_wrp_0/reg16x8_0/mem_14_[5]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_245_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_62_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_254_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_15_rs[5] , 
        \reg_apb_wrp_0/reg16x8_0/mem_15_[5]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_254_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_87_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_134_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_0_rs[6] , 
        \reg_apb_wrp_0/reg16x8_0/mem_0_[6]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_134_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_45_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_142_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_1_rs[6] , 
        \reg_apb_wrp_0/reg16x8_0/mem_1_[6]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_142_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_38_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_150_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_2_rs[6] , 
        \reg_apb_wrp_0/reg16x8_0/mem_2_[6]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_150_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_83_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_159_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_3_rs[6] , 
        \reg_apb_wrp_0/reg16x8_0/mem_3_[6]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_159_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_9_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_168_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_4_rs[6] , 
        \reg_apb_wrp_0/reg16x8_0/mem_4_[6]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_168_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_25_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_184_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_5_rs[6] , 
        \reg_apb_wrp_0/reg16x8_0/mem_5_[6]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_184_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_121_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_200_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_6_rs[6] , 
        \reg_apb_wrp_0/reg16x8_0/mem_6_[6]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_200_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_3_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_215_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_7_rs[6] , 
        \reg_apb_wrp_0/reg16x8_0/mem_7_[6]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_215_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_70_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_171_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_8_rs[6] , 
        \reg_apb_wrp_0/reg16x8_0/mem_8_[6]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_171_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_78_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_187_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_9_rs[6] , 
        \reg_apb_wrp_0/reg16x8_0/mem_9_[6]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_187_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_103_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_203_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_10_rs[6] , 
        \reg_apb_wrp_0/reg16x8_0/mem_10_[6]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_203_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_94_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_218_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_11_rs[6] , 
        \reg_apb_wrp_0/reg16x8_0/mem_11_[6]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_218_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_22_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_230_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_12_rs[6] , 
        \reg_apb_wrp_0/reg16x8_0/mem_12_[6]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_230_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_58_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_253_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_15_rs[4] , 
        \reg_apb_wrp_0/reg16x8_0/mem_15_[4]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_253_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_86_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_133_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_0_rs[5] , 
        \reg_apb_wrp_0/reg16x8_0/mem_0_[5]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_133_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_47_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_141_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_1_rs[5] , 
        \reg_apb_wrp_0/reg16x8_0/mem_1_[5]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_141_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_36_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_149_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_2_rs[5] , 
        \reg_apb_wrp_0/reg16x8_0/mem_2_[5]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_149_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_52_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_157_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_3_rs[5] , 
        \reg_apb_wrp_0/reg16x8_0/mem_3_[5]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_157_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_67_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_166_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_4_rs[5] , 
        \reg_apb_wrp_0/reg16x8_0/mem_4_[5]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_166_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_46_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_182_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_5_rs[5] , 
        \reg_apb_wrp_0/reg16x8_0/mem_5_[5]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_182_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_39_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_198_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_6_rs[5] , 
        \reg_apb_wrp_0/reg16x8_0/mem_6_[5]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_198_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_54_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_213_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_7_rs[5] , 
        \reg_apb_wrp_0/reg16x8_0/mem_7_[5]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_213_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_69_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_169_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_8_rs[5] , 
        \reg_apb_wrp_0/reg16x8_0/mem_8_[5]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_169_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_77_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_185_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_9_rs[5] , 
        \reg_apb_wrp_0/reg16x8_0/mem_9_[5]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_185_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_102_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_201_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_10_rs[5] , 
        \reg_apb_wrp_0/reg16x8_0/mem_10_[5]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_201_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_93_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_216_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_11_rs[5] , 
        \reg_apb_wrp_0/reg16x8_0/mem_11_[5]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_216_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_21_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_229_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_12_rs[5] , 
        \reg_apb_wrp_0/reg16x8_0/mem_12_[5]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_229_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_109_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_237_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_13_rs[5] , 
        \reg_apb_wrp_0/reg16x8_0/mem_13_[5]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_237_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_85_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_132_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_0_rs[4] , 
        \reg_apb_wrp_0/reg16x8_0/mem_0_[4]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_132_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_41_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_140_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_1_rs[4] , 
        \reg_apb_wrp_0/reg16x8_0/mem_1_[4]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_140_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_34_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_148_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_2_rs[4] , 
        \reg_apb_wrp_0/reg16x8_0/mem_2_[4]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_148_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_50_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_156_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_3_rs[4] , 
        \reg_apb_wrp_0/reg16x8_0/mem_3_[4]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_156_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_65_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_165_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_4_rs[4] , 
        \reg_apb_wrp_0/reg16x8_0/mem_4_[4]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_165_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_44_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_180_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_5_rs[4] , 
        \reg_apb_wrp_0/reg16x8_0/mem_5_[4]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_180_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_37_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_196_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_6_rs[4] , 
        \reg_apb_wrp_0/reg16x8_0/mem_6_[4]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_196_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_53_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_158_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_7_rs[4] , 
        \reg_apb_wrp_0/reg16x8_0/mem_7_[4]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_158_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_68_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_167_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_8_rs[4] , 
        \reg_apb_wrp_0/reg16x8_0/mem_8_[4]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_167_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_76_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_183_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_9_rs[4] , 
        \reg_apb_wrp_0/reg16x8_0/mem_9_[4]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_183_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_101_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_199_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_10_rs[4] , 
        \reg_apb_wrp_0/reg16x8_0/mem_10_[4]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_199_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_92_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_214_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_11_rs[4] , 
        \reg_apb_wrp_0/reg16x8_0/mem_11_[4]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_214_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_20_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_228_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_12_rs[4] , 
        \reg_apb_wrp_0/reg16x8_0/mem_12_[4]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_228_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_108_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_236_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_13_rs[4] , 
        \reg_apb_wrp_0/reg16x8_0/mem_13_[4]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_236_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_116_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_244_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_14_rs[4] , 
        \reg_apb_wrp_0/reg16x8_0/mem_14_[4]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_244_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_43_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_139_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_1_rs[3] , 
        \reg_apb_wrp_0/reg16x8_0/mem_1_[3]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_139_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_32_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_147_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_2_rs[3] , 
        \reg_apb_wrp_0/reg16x8_0/mem_2_[3]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_147_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_48_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_155_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_3_rs[3] , 
        \reg_apb_wrp_0/reg16x8_0/mem_3_[3]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_155_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_6_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_164_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_4_rs[3] , 
        \reg_apb_wrp_0/reg16x8_0/mem_4_[3]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_164_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_42_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_178_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_5_rs[3] , 
        \reg_apb_wrp_0/reg16x8_0/mem_5_[3]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_178_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_35_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_194_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_6_rs[3] , 
        \reg_apb_wrp_0/reg16x8_0/mem_6_[3]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_194_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_51_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_210_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_7_rs[3] , 
        \reg_apb_wrp_0/reg16x8_0/mem_7_[3]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_210_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_66_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_225_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_8_rs[3] , 
        \reg_apb_wrp_0/reg16x8_0/mem_8_[3]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_225_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_75_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_181_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_9_rs[3] , 
        \reg_apb_wrp_0/reg16x8_0/mem_9_[3]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_181_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_96_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_197_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_10_rs[3] , 
        \reg_apb_wrp_0/reg16x8_0/mem_10_[3]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_197_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_91_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_212_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_11_rs[3] , 
        \reg_apb_wrp_0/reg16x8_0/mem_11_[3]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_212_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_19_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_227_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_12_rs[3] , 
        \reg_apb_wrp_0/reg16x8_0/mem_12_[3]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_227_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_107_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_235_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_13_rs[3] , 
        \reg_apb_wrp_0/reg16x8_0/mem_13_[3]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_235_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_115_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_243_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_14_rs[3] , 
        \reg_apb_wrp_0/reg16x8_0/mem_14_[3]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_243_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_61_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_251_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_15_rs[3] , 
        \reg_apb_wrp_0/reg16x8_0/mem_15_[3]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_251_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_30_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_146_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_2_rs[2] , 
        \reg_apb_wrp_0/reg16x8_0/mem_2_[2]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_146_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_126_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_154_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_3_rs[2] , 
        \reg_apb_wrp_0/reg16x8_0/mem_3_[2]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_154_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_4_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_163_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_4_rs[2] , 
        \reg_apb_wrp_0/reg16x8_0/mem_4_[2]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_163_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_40_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_176_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_5_rs[2] , 
        \reg_apb_wrp_0/reg16x8_0/mem_5_[2]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_176_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_33_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_192_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_6_rs[2] , 
        \reg_apb_wrp_0/reg16x8_0/mem_6_[2]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_192_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_49_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_208_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_7_rs[2] , 
        \reg_apb_wrp_0/reg16x8_0/mem_7_[2]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_208_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_64_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_223_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_8_rs[2] , 
        \reg_apb_wrp_0/reg16x8_0/mem_8_[2]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_223_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_74_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_179_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_9_rs[2] , 
        \reg_apb_wrp_0/reg16x8_0/mem_9_[2]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_179_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_99_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_195_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_10_rs[2] , 
        \reg_apb_wrp_0/reg16x8_0/mem_10_[2]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_195_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_90_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_211_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_11_rs[2] , 
        \reg_apb_wrp_0/reg16x8_0/mem_11_[2]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_211_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_18_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_226_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_12_rs[2] , 
        \reg_apb_wrp_0/reg16x8_0/mem_12_[2]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_226_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_106_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_234_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_13_rs[2] , 
        \reg_apb_wrp_0/reg16x8_0/mem_13_[2]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_234_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_114_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_242_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_14_rs[2] , 
        \reg_apb_wrp_0/reg16x8_0/mem_14_[2]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_242_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_56_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_250_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_15_rs[2] , 
        \reg_apb_wrp_0/reg16x8_0/mem_15_[2]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_250_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_84_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_130_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_0_rs[3] , 
        \reg_apb_wrp_0/reg16x8_0/mem_0_[3]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_130_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_124_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_153_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_3_rs[1] , 
        \reg_apb_wrp_0/reg16x8_0/mem_3_[1]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_153_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_2_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_162_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_4_rs[1] , 
        \reg_apb_wrp_0/reg16x8_0/mem_4_[1]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_162_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_15_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_174_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_5_rs[1] , 
        \reg_apb_wrp_0/reg16x8_0/mem_5_[1]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_174_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_31_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_190_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_6_rs[1] , 
        \reg_apb_wrp_0/reg16x8_0/mem_6_[1]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_190_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_127_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_206_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_7_rs[1] , 
        \reg_apb_wrp_0/reg16x8_0/mem_7_[1]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_206_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_5_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_221_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_8_rs[1] , 
        \reg_apb_wrp_0/reg16x8_0/mem_8_[1]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_221_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_73_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_177_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_9_rs[1] , 
        \reg_apb_wrp_0/reg16x8_0/mem_9_[1]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_177_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_98_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_193_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_10_rs[1] , 
        \reg_apb_wrp_0/reg16x8_0/mem_10_[1]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_193_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_89_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_209_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_11_rs[1] , 
        \reg_apb_wrp_0/reg16x8_0/mem_11_[1]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_209_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_17_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_224_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_12_rs[1] , 
        \reg_apb_wrp_0/reg16x8_0/mem_12_[1]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_224_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_105_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_233_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_13_rs[1] , 
        \reg_apb_wrp_0/reg16x8_0/mem_13_[1]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_233_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_113_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_241_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_14_rs[1] , 
        \reg_apb_wrp_0/reg16x8_0/mem_14_[1]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_241_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_59_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_249_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_15_rs[1] , 
        \reg_apb_wrp_0/reg16x8_0/mem_15_[1]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_249_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_82_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_129_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_0_rs[2] , 
        \reg_apb_wrp_0/reg16x8_0/mem_0_[2]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_129_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_14_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_138_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_1_rs[2] , 
        \reg_apb_wrp_0/reg16x8_0/mem_1_[2]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_138_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_161_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_4_rs[0] , 
        \reg_apb_wrp_0/reg16x8_0/mem_4_[0]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_161_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_13_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_172_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_5_rs[0] , 
        \reg_apb_wrp_0/reg16x8_0/mem_5_[0]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_172_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_29_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_188_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_6_rs[0] , 
        \reg_apb_wrp_0/reg16x8_0/mem_6_[0]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_188_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_125_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_204_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_7_rs[0] , 
        \reg_apb_wrp_0/reg16x8_0/mem_7_[0]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_204_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_7_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_219_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_8_rs[0] , 
        \reg_apb_wrp_0/reg16x8_0/mem_8_[0]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_219_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_72_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_175_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_9_rs[0] , 
        \reg_apb_wrp_0/reg16x8_0/mem_9_[0]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_175_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_97_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_191_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_10_rs[0] , 
        \reg_apb_wrp_0/reg16x8_0/mem_10_[0]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_191_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_88_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_207_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_11_rs[0] , 
        \reg_apb_wrp_0/reg16x8_0/mem_11_[0]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_207_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_16_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_222_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_12_rs[0] , 
        \reg_apb_wrp_0/reg16x8_0/mem_12_[0]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_222_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_104_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_232_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_13_rs[0] , 
        \reg_apb_wrp_0/reg16x8_0/mem_13_[0]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_232_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_112_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_240_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_14_rs[0] , 
        \reg_apb_wrp_0/reg16x8_0/mem_14_[0]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_240_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_57_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_248_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_15_rs[0] , 
        \reg_apb_wrp_0/reg16x8_0/mem_15_[0]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_248_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_81_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_128_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_0_rs[1] , 
        \reg_apb_wrp_0/reg16x8_0/mem_0_[1]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_128_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_12_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_137_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_1_rs[1] , 
        \reg_apb_wrp_0/reg16x8_0/mem_1_[1]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_137_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_28_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_145_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_2_rs[1] , 
        \reg_apb_wrp_0/reg16x8_0/mem_2_[1]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_145_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_80_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_131_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_0_rs[0] , 
        \reg_apb_wrp_0/reg16x8_0/mem_0_[0]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_131_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_10_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_136_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_1_rs[0] , 
        \reg_apb_wrp_0/reg16x8_0/mem_1_[0]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_136_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_26_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_144_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_2_rs[0] , 
        \reg_apb_wrp_0/reg16x8_0/mem_2_[0]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_144_i , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_122_set_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_152_rs_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/mem_3_rs[0] , 
        \reg_apb_wrp_0/reg16x8_0/mem_3_[0]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_152_i , 
        \reg_apb_wrp_0/reg16x8_0/N_505 , 
        \reg_apb_wrp_0/reg16x8_0/N_504 , 
        \reg_apb_wrp_0/reg16x8_0/N_503 , 
        \reg_apb_wrp_0/reg16x8_0/N_502 , 
        \reg_apb_wrp_0/reg16x8_0/N_501 , 
        \reg_apb_wrp_0/reg16x8_0/N_500 , 
        \reg_apb_wrp_0/reg16x8_0/N_499 , 
        \reg_apb_wrp_0/reg16x8_0/N_498 , 
        \reg_apb_wrp_0/reg16x8_0/N_497 , 
        \reg_apb_wrp_0/reg16x8_0/N_496 , 
        \reg_apb_wrp_0/reg16x8_0/N_495 , 
        \reg_apb_wrp_0/reg16x8_0/N_494 , 
        \reg_apb_wrp_0/reg16x8_0/N_493 , 
        \reg_apb_wrp_0/reg16x8_0/N_492 , 
        \reg_apb_wrp_0/reg16x8_0/N_491 , 
        \reg_apb_wrp_0/reg16x8_0/N_490 , 
        \reg_apb_wrp_0/reg16x8_0/N_478 , 
        \reg_apb_wrp_0/reg16x8_0/N_470 , 
        \reg_apb_wrp_0/reg16x8_0/N_460 , 
        \reg_apb_wrp_0/reg16x8_0/N_458 , 
        \reg_apb_wrp_0/reg16x8_0/N_452 , 
        \reg_apb_wrp_0/reg16x8_0/N_450 , 
        \reg_apb_wrp_0/reg16x8_0/N_432 , 
        \reg_apb_wrp_0/reg16x8_0/N_414 , 
        \reg_apb_wrp_0/reg16x8_0/N_406 , 
        \reg_apb_wrp_0/reg16x8_0/N_400 , 
        \reg_apb_wrp_0/reg16x8_0/N_398 , 
        \reg_apb_wrp_0/reg16x8_0/N_392 , 
        \reg_apb_wrp_0/reg16x8_0/N_390 , 
        \reg_apb_wrp_0/reg16x8_0/N_382 , 
        \reg_apb_wrp_0/reg16x8_0/N_374 , 
        \reg_apb_wrp_0/reg16x8_0/N_368 , 
        \reg_apb_wrp_0/reg16x8_0/N_366 , 
        \reg_apb_wrp_0/reg16x8_0/N_360 , 
        \reg_apb_wrp_0/reg16x8_0/N_358 , 
        \reg_apb_wrp_0/reg16x8_0/N_350 , 
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_7[2]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_5[2]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_3[2]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_1[2]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_7[3]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_6[3]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_5[3]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_4[3]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_3[3]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_1[3]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_7[4]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_6[4]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_5[4]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_4[4]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_3[4]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_1[4]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_0[4]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_0_7[5]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_0_6[5]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_0_5[5]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_0_4[5]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_0_3[5]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_0_1[5]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_0_0[5]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_7[6]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_5[6]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_3[6]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_1[6]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_7[1]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_6[1]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_5[1]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_4[1]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_3[1]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_1[1]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_7[0]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_5[0]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_3[0]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_1[0]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_7[7]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_6[7]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_5[7]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_4[7]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_3[7]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_1[7]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_11[2]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_10[2]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_9[2]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_8[2]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_9[3]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_8[3]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_9[4]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_0_9[5]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_11[6]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_10[6]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_9[6]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_8[6]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_9[1]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_8[1]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_11[0]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_10[0]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_9[0]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_8[0]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_9[7]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_8[7]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_13[3]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_13[4]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_0_13[5]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_13[1]_net_1 , 
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_13[7]_net_1 , 
        \FIC_MSS_0/MSS_ADLIB_INST_MMUART0_TXD_USBC_DIR_MGPIO27B_OUT , 
        \FIC_MSS_0/MSS_ADLIB_INST_MMUART0_TXD_USBC_DIR_MGPIO27B_OE , 
        \FIC_MSS_0/MMUART_0_RXD_PAD_Y , 
        \FIC_MSS_0/MSS_ADLIB_INST_DRAM_WEN , 
        \FIC_MSS_0/MSS_ADLIB_INST_DRAM_RSTN , 
        \FIC_MSS_0/MSS_ADLIB_INST_DRAM_RASN , 
        \FIC_MSS_0/MSS_ADLIB_INST_DRAM_ODT , 
        \FIC_MSS_0/DRAM_FIFO_WE_OUT_net_0[0] , 
        \FIC_MSS_0/MDDR_DQS_TMATCH_0_IN_PAD_Y , 
        \FIC_MSS_0/MDDR_DQ_15_PAD_Y , 
        \FIC_MSS_0/DRAM_DQ_OUT_net_0[15] , 
        \FIC_MSS_0/DRAM_DQ_OE_net_0[15] , \FIC_MSS_0/MDDR_DQ_14_PAD_Y , 
        \FIC_MSS_0/DRAM_DQ_OUT_net_0[14] , 
        \FIC_MSS_0/DRAM_DQ_OE_net_0[14] , \FIC_MSS_0/MDDR_DQ_13_PAD_Y , 
        \FIC_MSS_0/DRAM_DQ_OUT_net_0[13] , 
        \FIC_MSS_0/DRAM_DQ_OE_net_0[13] , \FIC_MSS_0/MDDR_DQ_12_PAD_Y , 
        \FIC_MSS_0/DRAM_DQ_OUT_net_0[12] , 
        \FIC_MSS_0/DRAM_DQ_OE_net_0[12] , \FIC_MSS_0/MDDR_DQ_11_PAD_Y , 
        \FIC_MSS_0/DRAM_DQ_OUT_net_0[11] , 
        \FIC_MSS_0/DRAM_DQ_OE_net_0[11] , \FIC_MSS_0/MDDR_DQ_10_PAD_Y , 
        \FIC_MSS_0/DRAM_DQ_OUT_net_0[10] , 
        \FIC_MSS_0/DRAM_DQ_OE_net_0[10] , \FIC_MSS_0/MDDR_DQ_9_PAD_Y , 
        \FIC_MSS_0/DRAM_DQ_OUT_net_0[9] , 
        \FIC_MSS_0/DRAM_DQ_OE_net_0[9] , \FIC_MSS_0/MDDR_DQ_8_PAD_Y , 
        \FIC_MSS_0/DRAM_DQ_OUT_net_0[8] , 
        \FIC_MSS_0/DRAM_DQ_OE_net_0[8] , \FIC_MSS_0/MDDR_DQ_7_PAD_Y , 
        \FIC_MSS_0/DRAM_DQ_OUT_net_0[7] , 
        \FIC_MSS_0/DRAM_DQ_OE_net_0[7] , \FIC_MSS_0/MDDR_DQ_6_PAD_Y , 
        \FIC_MSS_0/DRAM_DQ_OUT_net_0[6] , 
        \FIC_MSS_0/DRAM_DQ_OE_net_0[6] , \FIC_MSS_0/MDDR_DQ_5_PAD_Y , 
        \FIC_MSS_0/DRAM_DQ_OUT_net_0[5] , 
        \FIC_MSS_0/DRAM_DQ_OE_net_0[5] , \FIC_MSS_0/MDDR_DQ_4_PAD_Y , 
        \FIC_MSS_0/DRAM_DQ_OUT_net_0[4] , 
        \FIC_MSS_0/DRAM_DQ_OE_net_0[4] , \FIC_MSS_0/MDDR_DQ_3_PAD_Y , 
        \FIC_MSS_0/DRAM_DQ_OUT_net_0[3] , 
        \FIC_MSS_0/DRAM_DQ_OE_net_0[3] , \FIC_MSS_0/MDDR_DQ_2_PAD_Y , 
        \FIC_MSS_0/DRAM_DQ_OUT_net_0[2] , 
        \FIC_MSS_0/DRAM_DQ_OE_net_0[2] , \FIC_MSS_0/MDDR_DQ_1_PAD_Y , 
        \FIC_MSS_0/DRAM_DQ_OUT_net_0[1] , 
        \FIC_MSS_0/DRAM_DQ_OE_net_0[1] , \FIC_MSS_0/MDDR_DQ_0_PAD_Y , 
        \FIC_MSS_0/DRAM_DQ_OUT_net_0[0] , 
        \FIC_MSS_0/DRAM_DQ_OE_net_0[0] , 
        \FIC_MSS_0/MDDR_DM_RDQS_1_PAD_Y , 
        \FIC_MSS_0/DRAM_DM_RDQS_OUT_net_0[1] , 
        \FIC_MSS_0/DM_OE_net_0[1] , \FIC_MSS_0/MDDR_DM_RDQS_0_PAD_Y , 
        \FIC_MSS_0/DRAM_DM_RDQS_OUT_net_0[0] , 
        \FIC_MSS_0/DM_OE_net_0[0] , 
        \FIC_MSS_0/MSS_ADLIB_INST_DRAM_CSN , 
        \FIC_MSS_0/MSS_ADLIB_INST_DRAM_CKE , 
        \FIC_MSS_0/MSS_ADLIB_INST_DRAM_CASN , 
        \FIC_MSS_0/DRAM_BA_net_0[2] , \FIC_MSS_0/DRAM_BA_net_0[1] , 
        \FIC_MSS_0/DRAM_BA_net_0[0] , \FIC_MSS_0/DRAM_ADDR_net_0[15] , 
        \FIC_MSS_0/DRAM_ADDR_net_0[14] , 
        \FIC_MSS_0/DRAM_ADDR_net_0[13] , 
        \FIC_MSS_0/DRAM_ADDR_net_0[12] , 
        \FIC_MSS_0/DRAM_ADDR_net_0[11] , 
        \FIC_MSS_0/DRAM_ADDR_net_0[10] , 
        \FIC_MSS_0/DRAM_ADDR_net_0[9] , \FIC_MSS_0/DRAM_ADDR_net_0[8] , 
        \FIC_MSS_0/DRAM_ADDR_net_0[7] , \FIC_MSS_0/DRAM_ADDR_net_0[6] , 
        \FIC_MSS_0/DRAM_ADDR_net_0[5] , \FIC_MSS_0/DRAM_ADDR_net_0[4] , 
        \FIC_MSS_0/DRAM_ADDR_net_0[3] , \FIC_MSS_0/DRAM_ADDR_net_0[2] , 
        \FIC_MSS_0/DRAM_ADDR_net_0[1] , \FIC_MSS_0/DRAM_ADDR_net_0[0] , 
        \FIC_MSS_0/CoreAPB3_0_APBmslave5_PRDATA_m_c_d[4] , 
        \FIC_MSS_0/CoreAPB3_0_APBmslave5_PRDATA_m_0_0[1] , 
        \FIC_MSS_0/CoreAPB3_0_APBmslave5_PRDATA_m_0_1_1[1] , 
        \FIC_MSS_0/FIC_MSS_0_FIC_0_APB_MASTER_PRDATA[1] , 
        \FIC_MSS_0/CoreAPB3_0_APBmslave5_PRDATA_m_0_1_0[1] , 
        \FIC_MSS_0/CoreAPB3_0_APBmslave5_PRDATA_m_0_0[5] , 
        \FIC_MSS_0/CoreAPB3_0_APBmslave5_PRDATA_m_0_1_1[5] , 
        \FIC_MSS_0/FIC_MSS_0_FIC_0_APB_MASTER_PRDATA[5] , 
        \FIC_MSS_0/CoreAPB3_0_APBmslave5_PRDATA_m_0_1_0[5] , 
        \FIC_MSS_0/CoreAPB3_0_APBmslave5_PRDATA_m_0_0[6] , 
        \FIC_MSS_0/CoreAPB3_0_APBmslave5_PRDATA_m_0_1_1[6] , 
        \FIC_MSS_0/FIC_MSS_0_FIC_0_APB_MASTER_PRDATA[6] , 
        \FIC_MSS_0/CoreAPB3_0_APBmslave5_PRDATA_m_0_1_0[6] , 
        \FIC_MSS_0/CoreAPB3_0_APBmslave5_PRDATA_m_0_0[2] , 
        \FIC_MSS_0/CoreAPB3_0_APBmslave5_PRDATA_m_0_1[2] , 
        \FIC_MSS_0/FIC_MSS_0_FIC_0_APB_MASTER_PRDATA[2] , 
        \FIC_MSS_0/CoreAPB3_0_APBmslave5_PRDATA_m_0_0[0] , 
        \FIC_MSS_0/CoreAPB3_0_APBmslave5_PRDATA_m_0_1[0] , 
        \FIC_MSS_0/FIC_MSS_0_FIC_0_APB_MASTER_PRDATA[0] , 
        \FIC_MSS_0/CoreAPB3_0_APBmslave5_PRDATA_m_0_1[4] , 
        \FIC_MSS_0/CoreAPB3_0_APBmslave5_PRDATA_m_0_1_0[4] , 
        \FIC_MSS_0/FIC_MSS_0_FIC_0_APB_MASTER_PRDATA[4] , 
        \FIC_MSS_0/CoreAPB3_0_APBmslave5_PRDATA_m_0_0[3] , 
        \FIC_MSS_0/CoreAPB3_0_APBmslave5_PRDATA_m_0_1[3] , 
        \FIC_MSS_0/CoreAPB3_0_APBmslave5_PRDATA_m_d[3] , 
        \FIC_MSS_0/FIC_MSS_0_FIC_0_APB_MASTER_PRDATA[3] , 
        \FIC_MSS_0/CoreAPB3_0_APBmslave5_PRDATA_m_c_c_0[5] , 
        \FIC_MSS_0/CoreAPB3_0_APBmslave5_PRDATA_m_c_c_0[1] , 
        \FIC_MSS_0/CoreAPB3_0_APBmslave5_PRDATA_m_c_c_0[6] , 
        \FIC_MSS_0/CoreAPB3_0_APBmslave5_PRDATA_m_c_c_1[3] , 
        \FIC_MSS_0/FIC_MSS_0_FIC_0_APB_MASTER_PREADY1_i_m_i_0 , 
        \FIC_MSS_0/CoreAPB3_0_APBmslave5_PRDATA_m_c_c[4] , 
        \FIC_MSS_0/MDDR_DQS_0_PAD_Y , \FIC_MSS_0/MDDR_DQS_1_PAD_Y , 
        \FIC_MSS_0/MSS_ADLIB_INST_DRAM_CLK , 
        \FIC_MSS_0/DRAM_DQS_OUT_net_0[0] , 
        \FIC_MSS_0/DRAM_DQS_OUT_net_0[1] , 
        \FIC_MSS_0/DRAM_DQS_OE_net_0[0] , 
        \FIC_MSS_0/DRAM_DQS_OE_net_0[1] , \CoreGPIO_0/edge_pos[31] , 
        \CoreGPIO_0/edge_neg_443[31] , 
        \CoreGPIO_0/edge_pos_2_sqmuxa_19_i_1 , 
        \CoreGPIO_0/edge_pos[30] , \CoreGPIO_0/edge_neg_429[30] , 
        \CoreGPIO_0/edge_neg_2_sqmuxa_6_i_1 , 
        \CoreGPIO_0/edge_pos[29] , \CoreGPIO_0/edge_neg_415[29] , 
        \CoreGPIO_0/N_190 , \CoreGPIO_0/edge_pos[28] , 
        \CoreGPIO_0/N_87_i_0 , \CoreGPIO_0/N_163 , 
        \CoreGPIO_0/edge_neg[27] , \CoreGPIO_0/N_5912_i_0 , 
        \CoreGPIO_0/N_161 , \CoreGPIO_0/edge_pos[26] , 
        \CoreGPIO_0/N_106_i_0 , \CoreGPIO_0/N_159 , 
        \CoreGPIO_0/edge_neg[25] , \CoreGPIO_0/N_5911_i_0 , 
        \CoreGPIO_0/N_157 , \CoreGPIO_0/edge_pos[24] , 
        \CoreGPIO_0/N_100_i_0 , \CoreGPIO_0/N_155 , 
        \CoreGPIO_0/edge_neg[23] , \CoreGPIO_0/N_96_i_0 , 
        \CoreGPIO_0/edge_pos_2_sqmuxa_26_i_1 , 
        \CoreGPIO_0/edge_neg[22] , \CoreGPIO_0/edge_neg_317[22] , 
        \CoreGPIO_0/N_200 , \CoreGPIO_0/edge_neg[21] , 
        \CoreGPIO_0/edge_neg_303[21] , \CoreGPIO_0/N_198 , 
        \CoreGPIO_0/edge_neg[20] , \CoreGPIO_0/edge_neg_289[20] , 
        \CoreGPIO_0/N_196 , \CoreGPIO_0/edge_neg[19] , 
        \CoreGPIO_0/edge_neg_275[19] , \CoreGPIO_0/N_194 , 
        \CoreGPIO_0/edge_neg[18] , \CoreGPIO_0/edge_neg_261[18] , 
        \CoreGPIO_0/N_192 , \CoreGPIO_0/edge_neg[17] , 
        \CoreGPIO_0/edge_neg_247[17] , 
        \CoreGPIO_0/edge_pos_2_sqmuxa_30_i_1 , 
        \CoreGPIO_0/edge_neg[16] , \CoreGPIO_0/edge_neg_233[16] , 
        \CoreGPIO_0/edge_pos_2_sqmuxa_29_i_1 , 
        \CoreGPIO_0/edge_neg[14] , \CoreGPIO_0/edge_neg_205[14] , 
        \CoreGPIO_0/edge_pos_2_sqmuxa_8_i_1 , 
        \CoreGPIO_0/edge_neg[13] , \CoreGPIO_0/edge_neg_191[13] , 
        \CoreGPIO_0/edge_pos_2_sqmuxa_9_i_1 , 
        \CoreGPIO_0/edge_neg[12] , \CoreGPIO_0/edge_neg_177[12] , 
        \CoreGPIO_0/N_188 , \CoreGPIO_0/edge_neg[11] , 
        \CoreGPIO_0/edge_neg_163[11] , \CoreGPIO_0/N_186 , 
        \CoreGPIO_0/edge_pos[10] , \CoreGPIO_0/edge_neg_149[10] , 
        \CoreGPIO_0/N_184 , \CoreGPIO_0/edge_neg[9] , 
        \CoreGPIO_0/edge_neg_135[9] , \CoreGPIO_0/N_182 , 
        \CoreGPIO_0/edge_pos[8] , \CoreGPIO_0/edge_neg_121[8] , 
        \CoreGPIO_0/edge_neg_2_sqmuxa_4_i_1 , \CoreGPIO_0/edge_pos[7] , 
        \CoreGPIO_0/N_83_i_0 , \CoreGPIO_0/edge_pos_2_sqmuxa_1_i_1 , 
        \CoreGPIO_0/edge_both[6] , \CoreGPIO_0/N_22_i_0 , 
        \CoreGPIO_0/N_78 , \CoreGPIO_0/edge_both[5] , 
        \CoreGPIO_0/N_89 , \CoreGPIO_0/N_76 , 
        \CoreGPIO_0/edge_both[4] , \CoreGPIO_0/N_91 , 
        \CoreGPIO_0/N_84 , \CoreGPIO_0/edge_both[3] , 
        \CoreGPIO_0/edge_both_51_iv_i_0[3] , 
        \CoreGPIO_0/edge_both_2_sqmuxa_12_i_1 , 
        \CoreGPIO_0/edge_both[2] , \CoreGPIO_0/N_93 , 
        \CoreGPIO_0/N_86 , \CoreGPIO_0/edge_both[1] , 
        \CoreGPIO_0/N_95 , \CoreGPIO_0/N_82 , 
        \CoreGPIO_0/edge_both[0] , \CoreGPIO_0/N_97 , 
        \CoreGPIO_0/N_80 , \CoreGPIO_0/edge_neg[6] , 
        \CoreGPIO_0/N_113 , \CoreGPIO_0/N_62 , 
        \CoreGPIO_0/edge_neg[5] , \CoreGPIO_0/N_115 , 
        \CoreGPIO_0/N_60 , \CoreGPIO_0/edge_neg[4] , 
        \CoreGPIO_0/N_117 , \CoreGPIO_0/N_58 , 
        \CoreGPIO_0/edge_neg[3] , \CoreGPIO_0/edge_neg_51_iv_i_1[3] , 
        \CoreGPIO_0/N_81 , \CoreGPIO_0/edge_neg[2] , 
        \CoreGPIO_0/N_119 , \CoreGPIO_0/N_56 , 
        \CoreGPIO_0/edge_neg[1] , \CoreGPIO_0/N_121 , 
        \CoreGPIO_0/N_54 , \CoreGPIO_0/edge_neg[0] , 
        \CoreGPIO_0/N_123 , \CoreGPIO_0/N_52 , 
        \CoreGPIO_0/edge_neg[15] , \CoreGPIO_0/edge_pos_219[15] , 
        \CoreGPIO_0/edge_pos_2_sqmuxa_7_i_1 , \CoreGPIO_0/edge_pos[6] , 
        \CoreGPIO_0/N_99 , \CoreGPIO_0/N_72 , \CoreGPIO_0/edge_pos[5] , 
        \CoreGPIO_0/N_101 , \CoreGPIO_0/N_70 , 
        \CoreGPIO_0/edge_pos[4] , \CoreGPIO_0/N_103 , 
        \CoreGPIO_0/N_68 , \CoreGPIO_0/edge_pos[3] , \CoreGPIO_0/N_73 , 
        \CoreGPIO_0/N_79 , \CoreGPIO_0/edge_pos[2] , 
        \CoreGPIO_0/N_105 , \CoreGPIO_0/N_64 , 
        \CoreGPIO_0/edge_pos[1] , \CoreGPIO_0/N_107 , 
        \CoreGPIO_0/N_66 , \CoreGPIO_0/edge_pos[0] , 
        \CoreGPIO_0/N_109 , \CoreGPIO_0/N_74 , 
        \CoreGPIO_0/GPOUT_reg_0_sqmuxa , \CoreGPIO_0/GPOUT_reg[26] , 
        \CoreGPIO_0/GPOUT_reg[18] , \CoreGPIO_0/GPOUT_reg[10] , 
        \CoreGPIO_0/GPOUT_reg[7] , \CoreGPIO_0/GPOUT_reg[3] , 
        \CoreGPIO_0/GPOUT_reg[2] , \CoreGPIO_0/GPOUT_reg[0] , 
        \CoreGPIO_0/CONFIG_reg[31][0] , \CoreGPIO_0/CONFIG_reg[31]2 , 
        \CoreGPIO_0/CONFIG_reg[31][1] , \CoreGPIO_0/CONFIG_reg[31][2] , 
        \CoreGPIO_0/CONFIG_reg[31][3] , \CoreGPIO_0/CONFIG_reg[31][4] , 
        \CoreGPIO_0/CONFIG_reg[31][5] , \CoreGPIO_0/CONFIG_reg[31][6] , 
        \CoreGPIO_0/CONFIG_reg[31][7] , \CoreGPIO_0/CONFIG_reg[30][0] , 
        \CoreGPIO_0/CONFIG_reg[30]2 , \CoreGPIO_0/CONFIG_reg[30][1] , 
        \CoreGPIO_0/CONFIG_reg[30][2] , \CoreGPIO_0/CONFIG_reg[30][3] , 
        \CoreGPIO_0/CONFIG_reg[30][4] , \CoreGPIO_0/CONFIG_reg[30][5] , 
        \CoreGPIO_0/CONFIG_reg[30][6] , \CoreGPIO_0/CONFIG_reg[30][7] , 
        \CoreGPIO_0/CONFIG_reg[29][0] , \CoreGPIO_0/CONFIG_reg[29]2 , 
        \CoreGPIO_0/CONFIG_reg[29][1] , \CoreGPIO_0/CONFIG_reg[29][2] , 
        \CoreGPIO_0/CONFIG_reg[29][3] , \CoreGPIO_0/CONFIG_reg[29][4] , 
        \CoreGPIO_0/CONFIG_reg[29][5] , \CoreGPIO_0/CONFIG_reg[29][6] , 
        \CoreGPIO_0/CONFIG_reg[29][7] , \CoreGPIO_0/CONFIG_reg[28][0] , 
        \CoreGPIO_0/CONFIG_reg[28]2 , \CoreGPIO_0/CONFIG_reg[28][1] , 
        \CoreGPIO_0/CONFIG_reg[28][2] , \CoreGPIO_0/CONFIG_reg[28][3] , 
        \CoreGPIO_0/CONFIG_reg[28][4] , \CoreGPIO_0/CONFIG_reg[28][5] , 
        \CoreGPIO_0/CONFIG_reg[28][6] , \CoreGPIO_0/CONFIG_reg[28][7] , 
        \CoreGPIO_0/CONFIG_reg[27][0] , \CoreGPIO_0/CONFIG_reg[27]2 , 
        \CoreGPIO_0/CONFIG_reg[27][1] , \CoreGPIO_0/CONFIG_reg[27][2] , 
        \CoreGPIO_0/CONFIG_reg[27][3] , \CoreGPIO_0/CONFIG_reg[27][4] , 
        \CoreGPIO_0/CONFIG_reg[27][5] , \CoreGPIO_0/CONFIG_reg[27][6] , 
        \CoreGPIO_0/CONFIG_reg[27][7] , \CoreGPIO_0/CONFIG_reg[26][0] , 
        \CoreGPIO_0/CONFIG_reg[26]2 , \CoreGPIO_0/CONFIG_reg[26][1] , 
        \CoreGPIO_0/CONFIG_reg[26][2] , \CoreGPIO_0/CONFIG_reg[26][3] , 
        \CoreGPIO_0/CONFIG_reg[26][4] , \CoreGPIO_0/CONFIG_reg[26][5] , 
        \CoreGPIO_0/CONFIG_reg[26][6] , \CoreGPIO_0/CONFIG_reg[26][7] , 
        \CoreGPIO_0/CONFIG_reg[25][0] , \CoreGPIO_0/CONFIG_reg[25]2 , 
        \CoreGPIO_0/CONFIG_reg[25][1] , \CoreGPIO_0/CONFIG_reg[25][2] , 
        \CoreGPIO_0/CONFIG_reg[25][3] , \CoreGPIO_0/CONFIG_reg[25][4] , 
        \CoreGPIO_0/CONFIG_reg[25][5] , \CoreGPIO_0/CONFIG_reg[25][6] , 
        \CoreGPIO_0/CONFIG_reg[25][7] , \CoreGPIO_0/CONFIG_reg[24][0] , 
        \CoreGPIO_0/CONFIG_reg[24]2 , \CoreGPIO_0/CONFIG_reg[24][1] , 
        \CoreGPIO_0/CONFIG_reg[24][2] , \CoreGPIO_0/CONFIG_reg[24][3] , 
        \CoreGPIO_0/CONFIG_reg[24][4] , \CoreGPIO_0/CONFIG_reg[24][5] , 
        \CoreGPIO_0/CONFIG_reg[24][6] , \CoreGPIO_0/CONFIG_reg[24][7] , 
        \CoreGPIO_0/CONFIG_reg[23][0] , \CoreGPIO_0/CONFIG_reg[23]2 , 
        \CoreGPIO_0/CONFIG_reg[23][1] , \CoreGPIO_0/CONFIG_reg[23][2] , 
        \CoreGPIO_0/CONFIG_reg[23][3] , \CoreGPIO_0/CONFIG_reg[23][4] , 
        \CoreGPIO_0/CONFIG_reg[23][5] , \CoreGPIO_0/CONFIG_reg[23][6] , 
        \CoreGPIO_0/CONFIG_reg[23][7] , \CoreGPIO_0/CONFIG_reg[22][0] , 
        \CoreGPIO_0/CONFIG_reg[22]2 , \CoreGPIO_0/CONFIG_reg[22][1] , 
        \CoreGPIO_0/CONFIG_reg[22][2] , \CoreGPIO_0/CONFIG_reg[22][3] , 
        \CoreGPIO_0/CONFIG_reg[22][4] , \CoreGPIO_0/CONFIG_reg[22][5] , 
        \CoreGPIO_0/CONFIG_reg[22][6] , \CoreGPIO_0/CONFIG_reg[22][7] , 
        \CoreGPIO_0/CONFIG_reg[21][0] , \CoreGPIO_0/CONFIG_reg[21]2 , 
        \CoreGPIO_0/CONFIG_reg[21][1] , \CoreGPIO_0/CONFIG_reg[21][2] , 
        \CoreGPIO_0/CONFIG_reg[21][3] , \CoreGPIO_0/CONFIG_reg[21][4] , 
        \CoreGPIO_0/CONFIG_reg[21][5] , \CoreGPIO_0/CONFIG_reg[21][6] , 
        \CoreGPIO_0/CONFIG_reg[21][7] , \CoreGPIO_0/CONFIG_reg[20][0] , 
        \CoreGPIO_0/CONFIG_reg[20]2 , \CoreGPIO_0/CONFIG_reg[20][1] , 
        \CoreGPIO_0/CONFIG_reg[20][2] , \CoreGPIO_0/CONFIG_reg[20][3] , 
        \CoreGPIO_0/CONFIG_reg[20][4] , \CoreGPIO_0/CONFIG_reg[20][5] , 
        \CoreGPIO_0/CONFIG_reg[20][6] , \CoreGPIO_0/CONFIG_reg[20][7] , 
        \CoreGPIO_0/CONFIG_reg[19][0] , \CoreGPIO_0/CONFIG_reg[19]2 , 
        \CoreGPIO_0/CONFIG_reg[19][1] , \CoreGPIO_0/CONFIG_reg[19][2] , 
        \CoreGPIO_0/CONFIG_reg[19][3] , \CoreGPIO_0/CONFIG_reg[19][4] , 
        \CoreGPIO_0/CONFIG_reg[19][5] , \CoreGPIO_0/CONFIG_reg[19][6] , 
        \CoreGPIO_0/CONFIG_reg[19][7] , \CoreGPIO_0/CONFIG_reg[18][0] , 
        \CoreGPIO_0/CONFIG_reg[18]2 , \CoreGPIO_0/CONFIG_reg[18][1] , 
        \CoreGPIO_0/CONFIG_reg[18][2] , \CoreGPIO_0/CONFIG_reg[18][3] , 
        \CoreGPIO_0/CONFIG_reg[18][4] , \CoreGPIO_0/CONFIG_reg[18][5] , 
        \CoreGPIO_0/CONFIG_reg[18][6] , \CoreGPIO_0/CONFIG_reg[18][7] , 
        \CoreGPIO_0/CONFIG_reg[17][0] , \CoreGPIO_0/CONFIG_reg[17]2 , 
        \CoreGPIO_0/CONFIG_reg[17][1] , \CoreGPIO_0/CONFIG_reg[17][2] , 
        \CoreGPIO_0/CONFIG_reg[17][3] , \CoreGPIO_0/CONFIG_reg[17][4] , 
        \CoreGPIO_0/CONFIG_reg[17][5] , \CoreGPIO_0/CONFIG_reg[17][6] , 
        \CoreGPIO_0/CONFIG_reg[17][7] , \CoreGPIO_0/CONFIG_reg[16][0] , 
        \CoreGPIO_0/CONFIG_reg[16]2 , \CoreGPIO_0/CONFIG_reg[16][1] , 
        \CoreGPIO_0/CONFIG_reg[16][2] , \CoreGPIO_0/CONFIG_reg[16][3] , 
        \CoreGPIO_0/CONFIG_reg[16][4] , \CoreGPIO_0/CONFIG_reg[16][5] , 
        \CoreGPIO_0/CONFIG_reg[16][6] , \CoreGPIO_0/CONFIG_reg[16][7] , 
        \CoreGPIO_0/CONFIG_reg[15][0] , \CoreGPIO_0/CONFIG_reg[15]2 , 
        \CoreGPIO_0/CONFIG_reg[15][1] , \CoreGPIO_0/CONFIG_reg[15][2] , 
        \CoreGPIO_0/CONFIG_reg[15][3] , \CoreGPIO_0/CONFIG_reg[15][4] , 
        \CoreGPIO_0/CONFIG_reg[15][5] , \CoreGPIO_0/CONFIG_reg[15][6] , 
        \CoreGPIO_0/CONFIG_reg[15][7] , \CoreGPIO_0/CONFIG_reg[14][0] , 
        \CoreGPIO_0/CONFIG_reg[14]2 , \CoreGPIO_0/CONFIG_reg[14][1] , 
        \CoreGPIO_0/CONFIG_reg[14][2] , \CoreGPIO_0/CONFIG_reg[14][3] , 
        \CoreGPIO_0/CONFIG_reg[14][4] , \CoreGPIO_0/CONFIG_reg[14][5] , 
        \CoreGPIO_0/CONFIG_reg[14][6] , \CoreGPIO_0/CONFIG_reg[14][7] , 
        \CoreGPIO_0/CONFIG_reg[13][0] , \CoreGPIO_0/CONFIG_reg[13]2 , 
        \CoreGPIO_0/CONFIG_reg[13][1] , \CoreGPIO_0/CONFIG_reg[13][2] , 
        \CoreGPIO_0/CONFIG_reg[13][3] , \CoreGPIO_0/CONFIG_reg[13][4] , 
        \CoreGPIO_0/CONFIG_reg[13][5] , \CoreGPIO_0/CONFIG_reg[13][6] , 
        \CoreGPIO_0/CONFIG_reg[13][7] , \CoreGPIO_0/CONFIG_reg[12][0] , 
        \CoreGPIO_0/CONFIG_reg[12]2 , \CoreGPIO_0/CONFIG_reg[12][1] , 
        \CoreGPIO_0/CONFIG_reg[12][2] , \CoreGPIO_0/CONFIG_reg[12][3] , 
        \CoreGPIO_0/CONFIG_reg[12][4] , \CoreGPIO_0/CONFIG_reg[12][5] , 
        \CoreGPIO_0/CONFIG_reg[12][6] , \CoreGPIO_0/CONFIG_reg[12][7] , 
        \CoreGPIO_0/CONFIG_reg[11][0] , \CoreGPIO_0/CONFIG_reg[11]2 , 
        \CoreGPIO_0/CONFIG_reg[11][1] , \CoreGPIO_0/CONFIG_reg[11][2] , 
        \CoreGPIO_0/CONFIG_reg[11][3] , \CoreGPIO_0/CONFIG_reg[11][4] , 
        \CoreGPIO_0/CONFIG_reg[11][5] , \CoreGPIO_0/CONFIG_reg[11][6] , 
        \CoreGPIO_0/CONFIG_reg[11][7] , \CoreGPIO_0/CONFIG_reg[10][0] , 
        \CoreGPIO_0/CONFIG_reg[10]2 , \CoreGPIO_0/CONFIG_reg[10][1] , 
        \CoreGPIO_0/CONFIG_reg[10][2] , \CoreGPIO_0/CONFIG_reg[10][3] , 
        \CoreGPIO_0/CONFIG_reg[10][4] , \CoreGPIO_0/CONFIG_reg[10][5] , 
        \CoreGPIO_0/CONFIG_reg[10][6] , \CoreGPIO_0/CONFIG_reg[10][7] , 
        \CoreGPIO_0/CONFIG_reg[9][0] , \CoreGPIO_0/CONFIG_reg[9]2 , 
        \CoreGPIO_0/CONFIG_reg[9][1] , \CoreGPIO_0/CONFIG_reg[9][2] , 
        \CoreGPIO_0/CONFIG_reg[9][3] , \CoreGPIO_0/CONFIG_reg[9][4] , 
        \CoreGPIO_0/CONFIG_reg[9][5] , \CoreGPIO_0/CONFIG_reg[9][6] , 
        \CoreGPIO_0/CONFIG_reg[9][7] , \CoreGPIO_0/CONFIG_reg[8][0] , 
        \CoreGPIO_0/CONFIG_reg[8]2 , \CoreGPIO_0/CONFIG_reg[8][1] , 
        \CoreGPIO_0/CONFIG_reg[8][2] , \CoreGPIO_0/CONFIG_reg[8][3] , 
        \CoreGPIO_0/CONFIG_reg[8][4] , \CoreGPIO_0/CONFIG_reg[8][5] , 
        \CoreGPIO_0/CONFIG_reg[8][6] , \CoreGPIO_0/CONFIG_reg[8][7] , 
        \CoreGPIO_0/CONFIG_reg[7][0] , \CoreGPIO_0/CONFIG_reg[7]2 , 
        \CoreGPIO_0/CONFIG_reg[7][1] , \CoreGPIO_0/CONFIG_reg[7][2] , 
        \CoreGPIO_0/CONFIG_reg[7][3] , \CoreGPIO_0/CONFIG_reg[7][4] , 
        \CoreGPIO_0/CONFIG_reg[7][5] , \CoreGPIO_0/CONFIG_reg[7][6] , 
        \CoreGPIO_0/CONFIG_reg[7][7] , \CoreGPIO_0/CONFIG_reg[6][0] , 
        \CoreGPIO_0/CONFIG_reg[6]2 , \CoreGPIO_0/CONFIG_reg[6][2] , 
        \CoreGPIO_0/CONFIG_reg[6][3] , \CoreGPIO_0/CONFIG_reg[6][4] , 
        \CoreGPIO_0/CONFIG_reg[6][5] , \CoreGPIO_0/CONFIG_reg[6][6] , 
        \CoreGPIO_0/CONFIG_reg[6][7] , \CoreGPIO_0/CONFIG_reg[5][0] , 
        \CoreGPIO_0/CONFIG_reg[5]2 , \CoreGPIO_0/CONFIG_reg[5][2] , 
        \CoreGPIO_0/CONFIG_reg[5][3] , \CoreGPIO_0/CONFIG_reg[5][4] , 
        \CoreGPIO_0/CONFIG_reg[5][5] , \CoreGPIO_0/CONFIG_reg[5][6] , 
        \CoreGPIO_0/CONFIG_reg[5][7] , \CoreGPIO_0/CONFIG_reg[4][0] , 
        \CoreGPIO_0/CONFIG_reg[4]2 , \CoreGPIO_0/CONFIG_reg[4][2] , 
        \CoreGPIO_0/CONFIG_reg[4][3] , \CoreGPIO_0/CONFIG_reg[4][4] , 
        \CoreGPIO_0/CONFIG_reg[4][5] , \CoreGPIO_0/CONFIG_reg[4][6] , 
        \CoreGPIO_0/CONFIG_reg[4][7] , \CoreGPIO_0/CONFIG_reg[3][0] , 
        \CoreGPIO_0/CONFIG_reg[3]2 , \CoreGPIO_0/CONFIG_reg[3][2] , 
        \CoreGPIO_0/CONFIG_reg[3][3] , \CoreGPIO_0/CONFIG_reg[3][4] , 
        \CoreGPIO_0/CONFIG_reg[3][5] , \CoreGPIO_0/CONFIG_reg[3][6] , 
        \CoreGPIO_0/CONFIG_reg[3][7] , \CoreGPIO_0/CONFIG_reg[2][0] , 
        \CoreGPIO_0/CONFIG_reg[2]2 , \CoreGPIO_0/CONFIG_reg[2][2] , 
        \CoreGPIO_0/CONFIG_reg[2][3] , \CoreGPIO_0/CONFIG_reg[2][4] , 
        \CoreGPIO_0/CONFIG_reg[2][5] , \CoreGPIO_0/CONFIG_reg[2][6] , 
        \CoreGPIO_0/CONFIG_reg[2][7] , \CoreGPIO_0/CONFIG_reg[1][0] , 
        \CoreGPIO_0/CONFIG_reg[1]2 , \CoreGPIO_0/CONFIG_reg[1][2] , 
        \CoreGPIO_0/CONFIG_reg[1][3] , \CoreGPIO_0/CONFIG_reg[1][4] , 
        \CoreGPIO_0/CONFIG_reg[1][5] , \CoreGPIO_0/CONFIG_reg[1][6] , 
        \CoreGPIO_0/CONFIG_reg[1][7] , \CoreGPIO_0/CONFIG_reg[0][0] , 
        \CoreGPIO_0/CONFIG_reg[0]2 , \CoreGPIO_0/CONFIG_reg[0][2] , 
        \CoreGPIO_0/CONFIG_reg[0][3] , \CoreGPIO_0/CONFIG_reg[0][4] , 
        \CoreGPIO_0/CONFIG_reg[0][5] , \CoreGPIO_0/CONFIG_reg[0][6] , 
        \CoreGPIO_0/CONFIG_reg[0][7] , \CoreGPIO_0/INTR_reg[23] , 
        \CoreGPIO_0/INTR_reg_308[23] , \CoreGPIO_0/INTR_reg[24] , 
        \CoreGPIO_0/INTR_reg_321[24] , \CoreGPIO_0/INTR_reg[25] , 
        \CoreGPIO_0/INTR_reg_334[25] , \CoreGPIO_0/INTR_reg_347[26] , 
        \CoreGPIO_0/INTR_reg[27] , \CoreGPIO_0/INTR_reg_360[27] , 
        \CoreGPIO_0/INTR_reg[28] , \CoreGPIO_0/INTR_reg_373[28] , 
        \CoreGPIO_0/INTR_reg[29] , \CoreGPIO_0/INTR_reg_386[29] , 
        \CoreGPIO_0/INTR_reg[30] , \CoreGPIO_0/INTR_reg_399[30] , 
        \CoreGPIO_0/INTR_reg[31] , \CoreGPIO_0/INTR_reg_412[31] , 
        \CoreGPIO_0/INTR_reg[8] , \CoreGPIO_0/INTR_reg_113[8] , 
        \CoreGPIO_0/INTR_reg[9] , \CoreGPIO_0/INTR_reg_126[9] , 
        \CoreGPIO_0/INTR_reg_139[10] , \CoreGPIO_0/INTR_reg[11] , 
        \CoreGPIO_0/INTR_reg_152[11] , \CoreGPIO_0/INTR_reg[12] , 
        \CoreGPIO_0/INTR_reg_165[12] , \CoreGPIO_0/INTR_reg[13] , 
        \CoreGPIO_0/INTR_reg_178[13] , \CoreGPIO_0/INTR_reg[14] , 
        \CoreGPIO_0/INTR_reg_191[14] , \CoreGPIO_0/INTR_reg[15] , 
        \CoreGPIO_0/INTR_reg_204[15] , \CoreGPIO_0/INTR_reg[16] , 
        \CoreGPIO_0/INTR_reg_217[16] , \CoreGPIO_0/INTR_reg[17] , 
        \CoreGPIO_0/INTR_reg_230[17] , \CoreGPIO_0/INTR_reg_243[18] , 
        \CoreGPIO_0/INTR_reg[19] , \CoreGPIO_0/INTR_reg_256[19] , 
        \CoreGPIO_0/INTR_reg[20] , \CoreGPIO_0/INTR_reg_269[20] , 
        \CoreGPIO_0/INTR_reg[21] , \CoreGPIO_0/INTR_reg_282[21] , 
        \CoreGPIO_0/INTR_reg[22] , \CoreGPIO_0/INTR_reg_295[22] , 
        \CoreGPIO_0/INTR_reg[0] , \CoreGPIO_0/INTR_reg_9[0] , 
        \CoreGPIO_0/INTR_reg_22[1] , \CoreGPIO_0/INTR_reg[2] , 
        \CoreGPIO_0/INTR_reg_35[2] , \CoreGPIO_0/INTR_reg_48[3] , 
        \CoreGPIO_0/INTR_reg_61[4] , \CoreGPIO_0/INTR_reg_74[5] , 
        \CoreGPIO_0/INTR_reg_87[6] , \CoreGPIO_0/INTR_reg[7] , 
        \CoreGPIO_0/INTR_reg_100[7] , \CoreGPIO_0/gpin2[4] , 
        \CoreGPIO_0/gpin2[5] , \CoreGPIO_0/gpin2[6] , 
        \CoreGPIO_0/gpin2[0] , \CoreGPIO_0/gpin2[1] , 
        \CoreGPIO_0/gpin2[2] , \CoreGPIO_0/gpin2[3] , 
        \CoreGPIO_0/gpin1[4] , \CoreGPIO_0/gpin1[5] , 
        \CoreGPIO_0/gpin1[6] , \CoreGPIO_0/gpin1[0] , 
        \CoreGPIO_0/gpin1[1] , \CoreGPIO_0/gpin1[2] , 
        \CoreGPIO_0/gpin1[3] , \CoreGPIO_0/un34_intr_u_ns_1 , 
        \CoreGPIO_0/un5_PRDATA_o_0_a2_0_o2_sx , 
        \CoreGPIO_0/CONFIG_reg_o_2_31_am[2]_net_1 , 
        \CoreGPIO_0/CONFIG_reg_o_2_31_bm[2]_net_1 , 
        \CoreGPIO_0/CONFIG_reg_o_2_31_am[6]_net_1 , 
        \CoreGPIO_0/CONFIG_reg_o_2_31_bm[6]_net_1 , 
        \CoreGPIO_0/CONFIG_reg_o_2_31_am[4]_net_1 , 
        \CoreGPIO_0/CONFIG_reg_o_2_31_bm[4]_net_1 , 
        \CoreGPIO_0/CONFIG_reg_o_2_31_am[1]_net_1 , 
        \CoreGPIO_0/CONFIG_reg_o_2_31_bm[1]_net_1 , 
        \CoreGPIO_0/CONFIG_reg_o_2_31_am[5]_net_1 , 
        \CoreGPIO_0/CONFIG_reg_o_2_31_bm[5]_net_1 , 
        \CoreGPIO_0/CONFIG_reg_o_2_31_am[0]_net_1 , 
        \CoreGPIO_0/CONFIG_reg_o_2_31_bm[0]_net_1 , 
        \CoreGPIO_0/CONFIG_reg_o_2_31_am_RNO[0]_net_1 , 
        \CoreGPIO_0/CONFIG_reg_o_2_31_am_1[0] , 
        \CoreGPIO_0/CONFIG_reg_o_2_31_am_RNO_0[0]_net_1 , 
        \CoreGPIO_0/CONFIG_reg_o_2_31_am_1_1_RNO[0]_net_1 , 
        \CoreGPIO_0/CONFIG_reg_o_2_31_am_1_RNO_0[0]_net_1 , 
        \CoreGPIO_0/CONFIG_reg_o_2_31_bm_RNO[0]_net_1 , 
        \CoreGPIO_0/CONFIG_reg_o_2_31_bm_1[0] , 
        \CoreGPIO_0/CONFIG_reg_o_2_31_bm_RNO_0[0]_net_1 , 
        \CoreGPIO_0/CONFIG_reg_o_2_31_bm_1_1_RNO[0]_net_1 , 
        \CoreGPIO_0/CONFIG_reg_o_2_31_bm_1_RNO_0[0]_net_1 , 
        \CoreGPIO_0/CONFIG_reg_o_2_31_am_RNO[1]_net_1 , 
        \CoreGPIO_0/CONFIG_reg_o_2_31_am_1[1] , 
        \CoreGPIO_0/CONFIG_reg_o_2_31_am_RNO_0[1]_net_1 , 
        \CoreGPIO_0/CONFIG_reg_o_2_31_am_1_1_RNO[1]_net_1 , 
        \CoreGPIO_0/CONFIG_reg_o_2_31_am_1_RNO_0[1]_net_1 , 
        \CoreGPIO_0/CONFIG_reg_o_2_31_bm_RNO[1]_net_1 , 
        \CoreGPIO_0/CONFIG_reg_o_2_31_bm_1[1] , 
        \CoreGPIO_0/CONFIG_reg_o_2_31_bm_RNO_0[1]_net_1 , 
        \CoreGPIO_0/CONFIG_reg_o_2_31_bm_1_1_RNO[1]_net_1 , 
        \CoreGPIO_0/CONFIG_reg_o_2_31_bm_1_RNO_0[1]_net_1 , 
        \CoreGPIO_0/CONFIG_reg_o_2_31_am_RNO[2]_net_1 , 
        \CoreGPIO_0/CONFIG_reg_o_2_31_am_1[2] , 
        \CoreGPIO_0/CONFIG_reg_o_2_31_am_RNO_0[2]_net_1 , 
        \CoreGPIO_0/CONFIG_reg_o_2_31_am_1_1_RNO[2]_net_1 , 
        \CoreGPIO_0/CONFIG_reg_o_2_31_am_1_RNO_0[2]_net_1 , 
        \CoreGPIO_0/CONFIG_reg_o_2_31_bm_RNO[2]_net_1 , 
        \CoreGPIO_0/CONFIG_reg_o_2_31_bm_1[2] , 
        \CoreGPIO_0/CONFIG_reg_o_2_31_bm_RNO_0[2]_net_1 , 
        \CoreGPIO_0/CONFIG_reg_o_2_31_bm_1_1_RNO[2]_net_1 , 
        \CoreGPIO_0/CONFIG_reg_o_2_31_bm_1_RNO_0[2]_net_1 , 
        \CoreGPIO_0/CONFIG_reg_o_2_31_am_RNO[3]_net_1 , 
        \CoreGPIO_0/CONFIG_reg_o_2_31_am_1[3] , 
        \CoreGPIO_0/CONFIG_reg_o_2_31_am_RNO_0[3]_net_1 , 
        \CoreGPIO_0/CONFIG_reg_o_2_31_am_1_1_RNO[3]_net_1 , 
        \CoreGPIO_0/CONFIG_reg_o_2_31_am_1_RNO_0[3]_net_1 , 
        \CoreGPIO_0/CONFIG_reg_o_2_31_bm_RNO[3]_net_1 , 
        \CoreGPIO_0/CONFIG_reg_o_2_31_bm_1[3] , 
        \CoreGPIO_0/CONFIG_reg_o_2_31_bm_RNO_0[3]_net_1 , 
        \CoreGPIO_0/CONFIG_reg_o_2_31_bm_1_1_RNO[3]_net_1 , 
        \CoreGPIO_0/CONFIG_reg_o_2_31_bm_1_RNO_0[3]_net_1 , 
        \CoreGPIO_0/CONFIG_reg_o_2_31_am_RNO[4]_net_1 , 
        \CoreGPIO_0/CONFIG_reg_o_2_31_am_1[4] , 
        \CoreGPIO_0/CONFIG_reg_o_2_31_am_RNO_0[4]_net_1 , 
        \CoreGPIO_0/CONFIG_reg_o_2_31_am_1_1_RNO[4]_net_1 , 
        \CoreGPIO_0/CONFIG_reg_o_2_31_am_1_RNO_0[4]_net_1 , 
        \CoreGPIO_0/CONFIG_reg_o_2_31_bm_RNO[4]_net_1 , 
        \CoreGPIO_0/CONFIG_reg_o_2_31_bm_1[4] , 
        \CoreGPIO_0/CONFIG_reg_o_2_31_bm_RNO_0[4]_net_1 , 
        \CoreGPIO_0/CONFIG_reg_o_2_31_bm_1_1_RNO[4]_net_1 , 
        \CoreGPIO_0/CONFIG_reg_o_2_31_bm_1_RNO_0[4]_net_1 , 
        \CoreGPIO_0/CONFIG_reg_o_2_31_am_RNO[5]_net_1 , 
        \CoreGPIO_0/CONFIG_reg_o_2_31_am_1[5] , 
        \CoreGPIO_0/CONFIG_reg_o_2_31_am_RNO_0[5]_net_1 , 
        \CoreGPIO_0/CONFIG_reg_o_2_31_am_1_1_RNO[5]_net_1 , 
        \CoreGPIO_0/CONFIG_reg_o_2_31_am_1_RNO_0[5]_net_1 , 
        \CoreGPIO_0/CONFIG_reg_o_2_31_bm_RNO[5]_net_1 , 
        \CoreGPIO_0/CONFIG_reg_o_2_31_bm_1[5] , 
        \CoreGPIO_0/CONFIG_reg_o_2_31_bm_RNO_0[5]_net_1 , 
        \CoreGPIO_0/CONFIG_reg_o_2_31_bm_1_1_RNO[5]_net_1 , 
        \CoreGPIO_0/CONFIG_reg_o_2_31_bm_1_RNO_0[5]_net_1 , 
        \CoreGPIO_0/CONFIG_reg_o_2_31_am_RNO[6]_net_1 , 
        \CoreGPIO_0/CONFIG_reg_o_2_31_am_1[6] , 
        \CoreGPIO_0/CONFIG_reg_o_2_31_am_RNO_0[6]_net_1 , 
        \CoreGPIO_0/CONFIG_reg_o_2_31_am_1_1_RNO[6]_net_1 , 
        \CoreGPIO_0/CONFIG_reg_o_2_31_am_1_RNO_0[6]_net_1 , 
        \CoreGPIO_0/CONFIG_reg_o_2_31_bm_RNO[6]_net_1 , 
        \CoreGPIO_0/CONFIG_reg_o_2_31_bm_1[6] , 
        \CoreGPIO_0/CONFIG_reg_o_2_31_bm_RNO_0[6]_net_1 , 
        \CoreGPIO_0/CONFIG_reg_o_2_31_bm_1_1_RNO[6]_net_1 , 
        \CoreGPIO_0/CONFIG_reg_o_2_31_bm_1_RNO_0[6]_net_1 , 
        \CoreGPIO_0/CONFIG_reg_o_2_31_am_RNO[7]_net_1 , 
        \CoreGPIO_0/CONFIG_reg_o_2_31_am_1[7] , 
        \CoreGPIO_0/CONFIG_reg_o_2_31_am_RNO_0[7]_net_1 , 
        \CoreGPIO_0/CONFIG_reg_o_2_31_am[7]_net_1 , 
        \CoreGPIO_0/CONFIG_reg_o_2_31_am_1_1_RNO[7]_net_1 , 
        \CoreGPIO_0/CONFIG_reg_o_2_31_am_1_RNO_0[7]_net_1 , 
        \CoreGPIO_0/CONFIG_reg_o_2_31_bm_RNO[7]_net_1 , 
        \CoreGPIO_0/CONFIG_reg_o_2_31_bm_1[7] , 
        \CoreGPIO_0/CONFIG_reg_o_2_31_bm_RNO_0[7]_net_1 , 
        \CoreGPIO_0/CONFIG_reg_o_2_31_bm[7]_net_1 , 
        \CoreGPIO_0/CONFIG_reg_o_2_31_bm_1_1_RNO[7]_net_1 , 
        \CoreGPIO_0/CONFIG_reg_o_2_31_bm_1_RNO_0[7]_net_1 , 
        \CoreGPIO_0/INTR_reg_9_0_0_50_tz_1 , 
        \CoreGPIO_0/INTR_reg_9_0_0_m2[0] , \CoreGPIO_0/N_1575_tz , 
        \CoreGPIO_0/INTR_reg_22_0_0_51_tz_1 , \CoreGPIO_0/N_177 , 
        \CoreGPIO_0/N_1576_tz , \CoreGPIO_0/INTR_reg_35_0_0_52_tz_1 , 
        \CoreGPIO_0/N_178 , \CoreGPIO_0/N_1577_tz , 
        \CoreGPIO_0/INTR_reg_61_0_0_53_tz_1 , \CoreGPIO_0/N_179 , 
        \CoreGPIO_0/N_1578_tz , \CoreGPIO_0/INTR_reg_74_0_0_54_tz_1 , 
        \CoreGPIO_0/INTR_reg_74_0_0_m2[5] , \CoreGPIO_0/N_1579_tz , 
        \CoreGPIO_0/INTR_reg_87_0_0_55_tz_1 , 
        \CoreGPIO_0/INTR_reg_87_0_0_m2[6] , \CoreGPIO_0/N_1580_tz , 
        \CoreGPIO_0/CONFIG_reg_o_2_3_1[1] , 
        \CoreGPIO_0/CONFIG_reg_o_2_3_1[5] , 
        \CoreGPIO_0/CONFIG_reg_o_2_3_1[2] , 
        \CoreGPIO_0/CONFIG_reg_o_2_3_1[0] , 
        \CoreGPIO_0/CONFIG_reg_o_2_6_1[3] , 
        \CoreGPIO_0/CONFIG_reg_o_2_3_1[3] , 
        \CoreGPIO_0/CONFIG_reg_o_2_6_1[6] , 
        \CoreGPIO_0/CONFIG_reg_o_2_6_1[7] , 
        \CoreGPIO_0/CONFIG_reg_o_2_6_1[4] , 
        \CoreGPIO_0/CONFIG_reg_o_2_3_1[4] , 
        \CoreGPIO_0/CONFIG_reg_o_2_6_1[1] , 
        \CoreGPIO_0/CONFIG_reg_o_2_6_1[2] , 
        \CoreGPIO_0/CONFIG_reg_o_2_3_1[6] , 
        \CoreGPIO_0/CONFIG_reg_o_2_6_1[5] , 
        \CoreGPIO_0/CONFIG_reg_o_2_13_1_1[2] , 
        \CoreGPIO_0/CONFIG_reg_o_2_13_1_1[3] , 
        \CoreGPIO_0/CONFIG_reg_o_2_13_1_1[0] , 
        \CoreGPIO_0/CONFIG_reg_o_2_13_1_1[1] , 
        \CoreGPIO_0/CONFIG_reg_o_2_3_1[7] , 
        \CoreGPIO_0/CONFIG_reg_o_2_13_1_1[7] , 
        \CoreGPIO_0/CONFIG_reg_o_2_13_1_1[4] , 
        \CoreGPIO_0/CONFIG_reg_o_2_13_1_1[5] , 
        \CoreGPIO_0/CONFIG_reg_o_2_6_1[0] , 
        \CoreGPIO_0/CONFIG_reg_o_2_21_1[0] , 
        \CoreGPIO_0/CONFIG_reg_o_2_21_1[1] , 
        \CoreGPIO_0/CONFIG_reg_o_2_21_1[2] , 
        \CoreGPIO_0/CONFIG_reg_o_2_21_1[3] , 
        \CoreGPIO_0/CONFIG_reg_o_2_21_1[4] , 
        \CoreGPIO_0/CONFIG_reg_o_2_21_1[5] , 
        \CoreGPIO_0/CONFIG_reg_o_2_21_1[6] , 
        \CoreGPIO_0/CONFIG_reg_o_2_21_1[7] , 
        \CoreGPIO_0/CONFIG_reg_o_2_13_1_1[6] , 
        \CoreGPIO_0/CONFIG_reg_o_2_18_1[7] , 
        \CoreGPIO_0/CONFIG_reg_o_2_10_1_1[5] , 
        \CoreGPIO_0/CONFIG_reg_o_2_10_1_1[6] , 
        \CoreGPIO_0/CONFIG_reg_o_2_10_1_1[7] , 
        \CoreGPIO_0/CONFIG_reg_o_2_25_1_1[7] , 
        \CoreGPIO_0/CONFIG_reg_o_2_18_1[0] , 
        \CoreGPIO_0/CONFIG_reg_o_2_18_1[1] , 
        \CoreGPIO_0/CONFIG_reg_o_2_18_1[2] , 
        \CoreGPIO_0/CONFIG_reg_o_2_18_1[3] , 
        \CoreGPIO_0/CONFIG_reg_o_2_18_1[4] , 
        \CoreGPIO_0/CONFIG_reg_o_2_18_1[5] , 
        \CoreGPIO_0/CONFIG_reg_o_2_18_1[6] , 
        \CoreGPIO_0/CONFIG_reg_o_2_10_1_1[4] , 
        \CoreGPIO_0/CONFIG_reg_o_2_28_1_1[7] , 
        \CoreGPIO_0/CONFIG_reg_o_2_25_1_1[5] , 
        \CoreGPIO_0/CONFIG_reg_o_2_25_1_1[6] , 
        \CoreGPIO_0/CONFIG_reg_o_2_28_1_1[1] , 
        \CoreGPIO_0/CONFIG_reg_o_2_10_1_1[0] , 
        \CoreGPIO_0/CONFIG_reg_o_2_10_1_1[1] , 
        \CoreGPIO_0/CONFIG_reg_o_2_28_1_1[0] , 
        \CoreGPIO_0/CONFIG_reg_o_2_10_1_1[3] , 
        \CoreGPIO_0/CONFIG_reg_o_2_28_1_1[6] , 
        \CoreGPIO_0/CONFIG_reg_o_2_25_1_1[4] , 
        \CoreGPIO_0/CONFIG_reg_o_2_10_1_1[2] , 
        \CoreGPIO_0/CONFIG_reg_o_2_28_1_1[4] , 
        \CoreGPIO_0/CONFIG_reg_o_2_28_1_1[2] , 
        \CoreGPIO_0/CONFIG_reg_o_2_28_1_1[3] , 
        \CoreGPIO_0/CONFIG_reg_o_2_25_1_1[0] , 
        \CoreGPIO_0/CONFIG_reg_o_2_28_1_1[5] , 
        \CoreGPIO_0/CONFIG_reg_o_2_25_1_1[3] , 
        \CoreGPIO_0/CONFIG_reg_o_2_25_1_1[1] , 
        \CoreGPIO_0/CONFIG_reg_o_2_25_1_1[2] , 
        \CoreGPIO_0/un34_intr_u_bm , \CoreGPIO_0/un34_intr , 
        \CoreGPIO_0/PRDATA_iv_0_0_a2_0_0[2]_net_1 , 
        \CoreGPIO_0/PRDATA_iv_0_0_a2_0_0[0]_net_1 , 
        \CoreGPIO_0/PRDATA_0_iv_0_0_a2_0_0[7]_net_1 , 
        \CoreGPIO_0/N_253_i , \CoreGPIO_0/N_252_i , \CoreGPIO_0/N_689 , 
        \CoreGPIO_0/N_688 , \CoreGPIO_0/N_687 , \CoreGPIO_0/N_686 , 
        \CoreGPIO_0/N_610 , \CoreGPIO_0/N_606 , \CoreGPIO_0/N_605 , 
        \CoreGPIO_0/N_603 , \CoreGPIO_0/N_144_i , \CoreGPIO_0/N_143_i , 
        \CoreGPIO_0/N_142_i , \CoreGPIO_0/N_141_i , 
        \CoreGPIO_0/N_139_i , \CoreGPIO_0/N_406 , \CoreGPIO_0/N_405 , 
        \CoreGPIO_0/N_402 , \CoreGPIO_0/N_401 , \CoreGPIO_0/N_400 , 
        \CoreGPIO_0/N_399 , \CoreGPIO_0/N_398 , \CoreGPIO_0/N_397 , 
        \CoreGPIO_0/N_396 , \CoreGPIO_0/N_395 , \CoreGPIO_0/N_171 , 
        \CoreGPIO_0/INTR_reg_87_0_0_m2_0[6] , \CoreGPIO_0/N_175 , 
        \CoreGPIO_0/N_174 , \CoreGPIO_0/N_173 , \CoreGPIO_0/N_172 , 
        \CoreGPIO_0/N_4549 , \CoreGPIO_0/N_243 , 
        \CoreGPIO_0/INTR_reg_269_0_o2_0[20] , 
        \CoreGPIO_0/INTR_reg_399_0_o2_0[30] , 
        \CoreGPIO_0/INTR_reg_217_0_o2_0[16] , 
        \CoreGPIO_0/INTR_reg_243_0_o2_0[18] , 
        \CoreGPIO_0/INTR_reg_191_0_o2_0[14] , 
        \CoreGPIO_0/INTR_reg_126_0_o2_0[9] , 
        \CoreGPIO_0/INTR_reg_139_0_o2_0[10] , 
        \CoreGPIO_0/INTR_reg_256_0_o2_0[19] , 
        \CoreGPIO_0/INTR_reg_100_0_o2_0[7] , 
        \CoreGPIO_0/INTR_reg_360_0_o2_0[27] , 
        \CoreGPIO_0/INTR_reg_178_0_o2_0[13] , 
        \CoreGPIO_0/INTR_reg_204_0_o2_0[15] , 
        \CoreGPIO_0/INTR_reg_230_0_o2_0[17] , 
        \CoreGPIO_0/INTR_reg_373_0_o2_0[28] , 
        \CoreGPIO_0/INTR_reg_386_0_o2_0[29] , 
        \CoreGPIO_0/INTR_reg_412_0_o2_0[31] , 
        \CoreGPIO_0/INTR_reg_282_0_o2_0[21] , 
        \CoreGPIO_0/INTR_reg_308_0_o2_0[23] , 
        \CoreGPIO_0/INTR_reg_321_0_o2_0[24] , 
        \CoreGPIO_0/INTR_reg_347_0_o2_0[26] , 
        \CoreGPIO_0/INTR_reg_295_0_o2_0[22] , 
        \CoreGPIO_0/INTR_reg_334_0_o2_0[25] , 
        \CoreGPIO_0/INTR_reg_113_0_o2_0[8] , 
        \CoreGPIO_0/INTR_reg_152_0_o2_0[11] , 
        \CoreGPIO_0/INTR_reg_165_0_o2_0[12] , 
        \CoreGPIO_0/INTR_reg_269_0_o2_1[20] , 
        \CoreGPIO_0/INTR_reg_399_0_o2_1[30] , 
        \CoreGPIO_0/INTR_reg_217_0_o2_1[16] , 
        \CoreGPIO_0/INTR_reg_243_0_o2_1[18] , 
        \CoreGPIO_0/INTR_reg_191_0_o2_1[14] , 
        \CoreGPIO_0/INTR_reg_126_0_o2_1[9] , 
        \CoreGPIO_0/INTR_reg_139_0_o2_1[10] , 
        \CoreGPIO_0/INTR_reg_256_0_o2_1[19] , 
        \CoreGPIO_0/INTR_reg_100_0_o2_1[7] , 
        \CoreGPIO_0/INTR_reg_360_0_o2_1[27] , 
        \CoreGPIO_0/INTR_reg_178_0_o2_1[13] , 
        \CoreGPIO_0/INTR_reg_204_0_o2_1[15] , 
        \CoreGPIO_0/INTR_reg_230_0_o2_1[17] , 
        \CoreGPIO_0/INTR_reg_373_0_o2_1[28] , 
        \CoreGPIO_0/INTR_reg_386_0_o2_1[29] , 
        \CoreGPIO_0/INTR_reg_412_0_o2_1[31] , 
        \CoreGPIO_0/INTR_reg_282_0_o2_1[21] , 
        \CoreGPIO_0/INTR_reg_308_0_o2_1[23] , 
        \CoreGPIO_0/INTR_reg_321_0_o2_1[24] , 
        \CoreGPIO_0/INTR_reg_347_0_o2_1[26] , 
        \CoreGPIO_0/INTR_reg_295_0_o2_1[22] , 
        \CoreGPIO_0/INTR_reg_334_0_o2_1[25] , 
        \CoreGPIO_0/INTR_reg_113_0_o2_1[8] , 
        \CoreGPIO_0/INTR_reg_152_0_o2_1[11] , 
        \CoreGPIO_0/INTR_reg_165_0_o2_1[12] , \CoreGPIO_0/INTR_reg21 , 
        \CoreGPIO_0/N_248 , \CoreGPIO_0/N_604 , \CoreGPIO_0/N_598 , 
        ff_to_start_net, \GPIO_OUT_obuf[6]/U0/DOUT1 , 
        \GPIO_OUT_obuf[6]/U0/DOUT , \GPIO_OUT_obuf[6]/U0/EOUT1 , 
        \GPIO_OUT_obuf[6]/U0/EOUT , \GPIO_OUT_obuf[5]/U0/DOUT1 , 
        \GPIO_OUT_obuf[5]/U0/DOUT , \GPIO_OUT_obuf[5]/U0/EOUT1 , 
        \GPIO_OUT_obuf[5]/U0/EOUT , \FIC_MSS_0/MDDR_DM_RDQS_1_PAD/YIN , 
        \GPIO_IN_ibuf[6]/U0/YIN1 , \GPIO_IN_ibuf[6]/U0/YIN , 
        \FIC_MSS_0/MDDR_DQ_15_PAD/YIN , \GPIO_OUT_obuf[4]/U0/DOUT1 , 
        \GPIO_OUT_obuf[4]/U0/DOUT , \GPIO_OUT_obuf[4]/U0/EOUT1 , 
        \GPIO_OUT_obuf[4]/U0/EOUT , \FIC_MSS_0/MDDR_ADDR_10_PAD/EOUT , 
        \FIC_MSS_0/MDDR_CAS_N_PAD/EOUT , 
        \FIC_MSS_0/MDDR_DQ_10_PAD/YIN , 
        \FIC_MSS_0/MDDR_ADDR_5_PAD/EOUT , 
        \FIC_MSS_0/MDDR_CS_N_PAD/EOUT , 
        \FIC_MSS_0/MDDR_ADDR_15_PAD/EOUT , 
        \FIC_MSS_0/MDDR_ODT_PAD/EOUT , \FIC_MSS_0/MDDR_DQ_8_PAD/YIN , 
        \FIC_MSS_0/MDDR_RAS_N_PAD/EOUT , \GPIO_IN_ibuf[3]/U0/YIN1 , 
        \GPIO_IN_ibuf[3]/U0/YIN , \FIC_MSS_0/MDDR_ADDR_14_PAD/EOUT , 
        \FIC_MSS_0/MDDR_DQ_5_PAD/YIN , \FIC_MSS_0/MDDR_DQ_14_PAD/YIN , 
        \GPIO_IN_ibuf[2]/U0/YIN1 , \GPIO_IN_ibuf[2]/U0/YIN , 
        \GPIO_IN_ibuf[4]/U0/YIN1 , \GPIO_IN_ibuf[4]/U0/YIN , 
        \FIC_MSS_0/MDDR_CKE_PAD/EOUT , \FIC_MSS_0/MDDR_DQ_2_PAD/YIN , 
        \FIC_MSS_0/MDDR_ADDR_2_PAD/EOUT , \GPIO_IN_ibuf[1]/U0/YIN1 , 
        \GPIO_IN_ibuf[1]/U0/YIN , \FIC_MSS_0/MDDR_DQ_7_PAD/YIN , 
        \FIC_MSS_0/MDDR_ADDR_11_PAD/EOUT , 
        \MSS_RESET_N_F2M_ibuf/U0/YIN1 , \MSS_RESET_N_F2M_ibuf/U0/YIN , 
        \FIC_MSS_0/MDDR_ADDR_4_PAD/EOUT , 
        \FIC_MSS_0/MDDR_ADDR_1_PAD/EOUT , 
        \FIC_MSS_0/MDDR_DQS_TMATCH_0_OUT_PAD/EOUT , 
        \GPIO_OUT_obuf[3]/U0/DOUT1 , \GPIO_OUT_obuf[3]/U0/DOUT , 
        \GPIO_OUT_obuf[3]/U0/EOUT1 , \GPIO_OUT_obuf[3]/U0/EOUT , 
        \GPIO_IN_ibuf[0]/U0/YIN1 , \GPIO_IN_ibuf[0]/U0/YIN , 
        \FIC_MSS_0/MDDR_DQS_0_PAD/U2_N2P , 
        \FIC_MSS_0/MDDR_DQS_0_PAD/YIN , \GPIO_OUT_obuf[1]/U0/DOUT1 , 
        \GPIO_OUT_obuf[1]/U0/DOUT , \GPIO_OUT_obuf[1]/U0/EOUT1 , 
        \GPIO_OUT_obuf[1]/U0/EOUT , \GPIO_IN_ibuf[5]/U0/YIN1 , 
        \GPIO_IN_ibuf[5]/U0/YIN , \FIC_MSS_0/MDDR_ADDR_0_PAD/EOUT , 
        \FCCC_0/CCC_INST/CLK0_net , \FCCC_0/CCC_INST/CLK1_net , 
        \FCCC_0/CCC_INST/CLK2_net , \FCCC_0/CCC_INST/CLK3_net , 
        \FCCC_0/CCC_INST/NGMUX0_SEL_net , 
        \FCCC_0/CCC_INST/NGMUX1_SEL_net , 
        \FCCC_0/CCC_INST/NGMUX2_SEL_net , 
        \FCCC_0/CCC_INST/NGMUX3_SEL_net , 
        \FCCC_0/CCC_INST/NGMUX0_HOLD_N_net , 
        \FCCC_0/CCC_INST/NGMUX1_HOLD_N_net , 
        \FCCC_0/CCC_INST/NGMUX2_HOLD_N_net , 
        \FCCC_0/CCC_INST/NGMUX3_HOLD_N_net , 
        \FCCC_0/CCC_INST/NGMUX0_ARST_N_net , 
        \FCCC_0/CCC_INST/NGMUX1_ARST_N_net , 
        \FCCC_0/CCC_INST/NGMUX2_ARST_N_net , 
        \FCCC_0/CCC_INST/NGMUX3_ARST_N_net , 
        \FCCC_0/CCC_INST/PLL_BYPASS_N_net , 
        \FCCC_0/CCC_INST/PLL_ARST_N_net , 
        \FCCC_0/CCC_INST/PLL_POWERDOWN_N_net , 
        \FCCC_0/CCC_INST/GPD0_ARST_N_net , 
        \FCCC_0/CCC_INST/GPD1_ARST_N_net , 
        \FCCC_0/CCC_INST/GPD2_ARST_N_net , 
        \FCCC_0/CCC_INST/GPD3_ARST_N_net , 
        \FCCC_0/CCC_INST/PRESET_N_net , \FCCC_0/CCC_INST/PCLK_net , 
        \FCCC_0/CCC_INST/PSEL_net , \FCCC_0/CCC_INST/PENABLE_net , 
        \FCCC_0/CCC_INST/PWRITE_net , \FCCC_0/CCC_INST/PADDR_net[7] , 
        \FCCC_0/CCC_INST/PADDR_net[6] , \FCCC_0/CCC_INST/PADDR_net[5] , 
        \FCCC_0/CCC_INST/PADDR_net[4] , \FCCC_0/CCC_INST/PADDR_net[3] , 
        \FCCC_0/CCC_INST/PADDR_net[2] , 
        \FCCC_0/CCC_INST/PWDATA_net[7] , 
        \FCCC_0/CCC_INST/PWDATA_net[6] , 
        \FCCC_0/CCC_INST/PWDATA_net[5] , 
        \FCCC_0/CCC_INST/PWDATA_net[4] , 
        \FCCC_0/CCC_INST/PWDATA_net[3] , 
        \FCCC_0/CCC_INST/PWDATA_net[2] , 
        \FCCC_0/CCC_INST/PWDATA_net[1] , 
        \FCCC_0/CCC_INST/PWDATA_net[0] , \GPIO_OUT_obuf[2]/U0/DOUT1 , 
        \GPIO_OUT_obuf[2]/U0/DOUT , \GPIO_OUT_obuf[2]/U0/EOUT1 , 
        \GPIO_OUT_obuf[2]/U0/EOUT , \FIC_MSS_0/MDDR_DQ_3_PAD/YIN , 
        \FIC_MSS_0/MDDR_DQS_TMATCH_0_IN_PAD/YIN , 
        \FIC_MSS_0/MDDR_WE_N_PAD/EOUT , \FIC_MSS_0/MDDR_DQ_1_PAD/YIN , 
        \GPIO_OUT_obuf[0]/U0/DOUT1 , \GPIO_OUT_obuf[0]/U0/DOUT , 
        \GPIO_OUT_obuf[0]/U0/EOUT1 , \GPIO_OUT_obuf[0]/U0/EOUT , 
        \FIC_MSS_0/MDDR_BA_1_PAD/EOUT , 
        \FIC_MSS_0/MDDR_RESET_N_PAD/EOUT , 
        \FIC_MSS_0/MDDR_DQ_4_PAD/YIN , 
        \FIC_MSS_0/MSS_ADLIB_INST/CAN_RXBUS_F2H_SCP_net , 
        \FIC_MSS_0/MSS_ADLIB_INST/CAN_TX_EBL_F2H_SCP_net , 
        \FIC_MSS_0/MSS_ADLIB_INST/CAN_TXBUS_F2H_SCP_net , 
        \FIC_MSS_0/MSS_ADLIB_INST/COLF_net , 
        \FIC_MSS_0/MSS_ADLIB_INST/CRSF_net , 
        \FIC_MSS_0/MSS_ADLIB_INST/F2_DMAREADY_net[1] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F2_DMAREADY_net[0] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[15] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[14] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[13] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[12] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[11] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[10] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[9] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[8] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[7] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[6] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[5] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[4] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[3] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[2] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[1] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[0] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F2HCALIB_net , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_DMAREADY_net[1] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_DMAREADY_net[0] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[31] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[30] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[29] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[28] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[27] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[26] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[25] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[24] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[23] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[22] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[21] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[20] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[19] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[18] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[17] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[16] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[15] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[14] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[13] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[12] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[11] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[10] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[9] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[8] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[7] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[6] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[5] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[4] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[3] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[2] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[1] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[0] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_ENABLE_net , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_MASTLOCK_net , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_READY_net , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_SEL_net , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_SIZE_net[1] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_SIZE_net[0] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_TRANS1_net , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[31] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[30] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[29] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[28] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[27] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[26] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[25] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[24] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[23] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[22] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[21] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[20] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[19] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[18] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[17] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[16] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[15] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[14] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[13] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[12] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[11] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[10] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[9] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[8] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[7] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[6] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[5] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[4] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[3] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[2] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[1] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[0] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_WRITE_net , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[31] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[30] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[29] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[28] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[27] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[26] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[25] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[24] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[23] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[22] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[21] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[20] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[19] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[18] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[17] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[16] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[15] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[14] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[13] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[12] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[11] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[10] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[9] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[8] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[7] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[6] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[5] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[4] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[3] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[2] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[1] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[0] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_HM0_READY_net , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_HM0_RESP_net , 
        \FIC_MSS_0/MSS_ADLIB_INST/FAB_AVALID_net , 
        \FIC_MSS_0/MSS_ADLIB_INST/FAB_HOSTDISCON_net , 
        \FIC_MSS_0/MSS_ADLIB_INST/FAB_IDDIG_net , 
        \FIC_MSS_0/MSS_ADLIB_INST/FAB_LINESTATE_net[1] , 
        \FIC_MSS_0/MSS_ADLIB_INST/FAB_LINESTATE_net[0] , 
        \FIC_MSS_0/MSS_ADLIB_INST/FAB_M3_RESET_N_net , 
        \FIC_MSS_0/MSS_ADLIB_INST/FAB_PLL_LOCK_net , 
        \FIC_MSS_0/MSS_ADLIB_INST/FAB_RXACTIVE_net , 
        \FIC_MSS_0/MSS_ADLIB_INST/FAB_RXERROR_net , 
        \FIC_MSS_0/MSS_ADLIB_INST/FAB_RXVALID_net , 
        \FIC_MSS_0/MSS_ADLIB_INST/FAB_RXVALIDH_net , 
        \FIC_MSS_0/MSS_ADLIB_INST/FAB_SESSEND_net , 
        \FIC_MSS_0/MSS_ADLIB_INST/FAB_TXREADY_net , 
        \FIC_MSS_0/MSS_ADLIB_INST/FAB_VBUSVALID_net , 
        \FIC_MSS_0/MSS_ADLIB_INST/FAB_VSTATUS_net[7] , 
        \FIC_MSS_0/MSS_ADLIB_INST/FAB_VSTATUS_net[6] , 
        \FIC_MSS_0/MSS_ADLIB_INST/FAB_VSTATUS_net[5] , 
        \FIC_MSS_0/MSS_ADLIB_INST/FAB_VSTATUS_net[4] , 
        \FIC_MSS_0/MSS_ADLIB_INST/FAB_VSTATUS_net[3] , 
        \FIC_MSS_0/MSS_ADLIB_INST/FAB_VSTATUS_net[2] , 
        \FIC_MSS_0/MSS_ADLIB_INST/FAB_VSTATUS_net[1] , 
        \FIC_MSS_0/MSS_ADLIB_INST/FAB_VSTATUS_net[0] , 
        \FIC_MSS_0/MSS_ADLIB_INST/FAB_XDATAIN_net[7] , 
        \FIC_MSS_0/MSS_ADLIB_INST/FAB_XDATAIN_net[6] , 
        \FIC_MSS_0/MSS_ADLIB_INST/FAB_XDATAIN_net[5] , 
        \FIC_MSS_0/MSS_ADLIB_INST/FAB_XDATAIN_net[4] , 
        \FIC_MSS_0/MSS_ADLIB_INST/FAB_XDATAIN_net[3] , 
        \FIC_MSS_0/MSS_ADLIB_INST/FAB_XDATAIN_net[2] , 
        \FIC_MSS_0/MSS_ADLIB_INST/FAB_XDATAIN_net[1] , 
        \FIC_MSS_0/MSS_ADLIB_INST/FAB_XDATAIN_net[0] , 
        \FIC_MSS_0/MSS_ADLIB_INST/GTX_CLKPF_net , 
        \FIC_MSS_0/MSS_ADLIB_INST/I2C0_BCLK_net , 
        \FIC_MSS_0/MSS_ADLIB_INST/I2C0_SCL_F2H_SCP_net , 
        \FIC_MSS_0/MSS_ADLIB_INST/I2C0_SDA_F2H_SCP_net , 
        \FIC_MSS_0/MSS_ADLIB_INST/I2C1_BCLK_net , 
        \FIC_MSS_0/MSS_ADLIB_INST/I2C1_SCL_F2H_SCP_net , 
        \FIC_MSS_0/MSS_ADLIB_INST/I2C1_SDA_F2H_SCP_net , 
        \FIC_MSS_0/MSS_ADLIB_INST/MDIF_net , 
        \FIC_MSS_0/MSS_ADLIB_INST/MGPIO0A_F2H_GPIN_net , 
        \FIC_MSS_0/MSS_ADLIB_INST/MGPIO10A_F2H_GPIN_net , 
        \FIC_MSS_0/MSS_ADLIB_INST/MGPIO11A_F2H_GPIN_net , 
        \FIC_MSS_0/MSS_ADLIB_INST/MGPIO11B_F2H_GPIN_net , 
        \FIC_MSS_0/MSS_ADLIB_INST/MGPIO12A_F2H_GPIN_net , 
        \FIC_MSS_0/MSS_ADLIB_INST/MGPIO13A_F2H_GPIN_net , 
        \FIC_MSS_0/MSS_ADLIB_INST/MGPIO14A_F2H_GPIN_net , 
        \FIC_MSS_0/MSS_ADLIB_INST/MGPIO15A_F2H_GPIN_net , 
        \FIC_MSS_0/MSS_ADLIB_INST/MGPIO16A_F2H_GPIN_net , 
        \FIC_MSS_0/MSS_ADLIB_INST/MGPIO17B_F2H_GPIN_net , 
        \FIC_MSS_0/MSS_ADLIB_INST/MGPIO18B_F2H_GPIN_net , 
        \FIC_MSS_0/MSS_ADLIB_INST/MGPIO19B_F2H_GPIN_net , 
        \FIC_MSS_0/MSS_ADLIB_INST/MGPIO1A_F2H_GPIN_net , 
        \FIC_MSS_0/MSS_ADLIB_INST/MGPIO20B_F2H_GPIN_net , 
        \FIC_MSS_0/MSS_ADLIB_INST/MGPIO21B_F2H_GPIN_net , 
        \FIC_MSS_0/MSS_ADLIB_INST/MGPIO22B_F2H_GPIN_net , 
        \FIC_MSS_0/MSS_ADLIB_INST/MGPIO24B_F2H_GPIN_net , 
        \FIC_MSS_0/MSS_ADLIB_INST/MGPIO25B_F2H_GPIN_net , 
        \FIC_MSS_0/MSS_ADLIB_INST/MGPIO26B_F2H_GPIN_net , 
        \FIC_MSS_0/MSS_ADLIB_INST/MGPIO27B_F2H_GPIN_net , 
        \FIC_MSS_0/MSS_ADLIB_INST/MGPIO28B_F2H_GPIN_net , 
        \FIC_MSS_0/MSS_ADLIB_INST/MGPIO29B_F2H_GPIN_net , 
        \FIC_MSS_0/MSS_ADLIB_INST/MGPIO2A_F2H_GPIN_net , 
        \FIC_MSS_0/MSS_ADLIB_INST/MGPIO30B_F2H_GPIN_net , 
        \FIC_MSS_0/MSS_ADLIB_INST/MGPIO31B_F2H_GPIN_net , 
        \FIC_MSS_0/MSS_ADLIB_INST/MGPIO3A_F2H_GPIN_net , 
        \FIC_MSS_0/MSS_ADLIB_INST/MGPIO4A_F2H_GPIN_net , 
        \FIC_MSS_0/MSS_ADLIB_INST/MGPIO5A_F2H_GPIN_net , 
        \FIC_MSS_0/MSS_ADLIB_INST/MGPIO6A_F2H_GPIN_net , 
        \FIC_MSS_0/MSS_ADLIB_INST/MGPIO7A_F2H_GPIN_net , 
        \FIC_MSS_0/MSS_ADLIB_INST/MGPIO8A_F2H_GPIN_net , 
        \FIC_MSS_0/MSS_ADLIB_INST/MGPIO9A_F2H_GPIN_net , 
        \FIC_MSS_0/MSS_ADLIB_INST/MMUART0_CTS_F2H_SCP_net , 
        \FIC_MSS_0/MSS_ADLIB_INST/MMUART0_DCD_F2H_SCP_net , 
        \FIC_MSS_0/MSS_ADLIB_INST/MMUART0_DSR_F2H_SCP_net , 
        \FIC_MSS_0/MSS_ADLIB_INST/MMUART0_DTR_F2H_SCP_net , 
        \FIC_MSS_0/MSS_ADLIB_INST/MMUART0_RI_F2H_SCP_net , 
        \FIC_MSS_0/MSS_ADLIB_INST/MMUART0_RTS_F2H_SCP_net , 
        \FIC_MSS_0/MSS_ADLIB_INST/MMUART0_RXD_F2H_SCP_net , 
        \FIC_MSS_0/MSS_ADLIB_INST/MMUART0_SCK_F2H_SCP_net , 
        \FIC_MSS_0/MSS_ADLIB_INST/MMUART0_TXD_F2H_SCP_net , 
        \FIC_MSS_0/MSS_ADLIB_INST/MMUART1_CTS_F2H_SCP_net , 
        \FIC_MSS_0/MSS_ADLIB_INST/MMUART1_DCD_F2H_SCP_net , 
        \FIC_MSS_0/MSS_ADLIB_INST/MMUART1_DSR_F2H_SCP_net , 
        \FIC_MSS_0/MSS_ADLIB_INST/MMUART1_RI_F2H_SCP_net , 
        \FIC_MSS_0/MSS_ADLIB_INST/MMUART1_RTS_F2H_SCP_net , 
        \FIC_MSS_0/MSS_ADLIB_INST/MMUART1_RXD_F2H_SCP_net , 
        \FIC_MSS_0/MSS_ADLIB_INST/MMUART1_SCK_F2H_SCP_net , 
        \FIC_MSS_0/MSS_ADLIB_INST/MMUART1_TXD_F2H_SCP_net , 
        \FIC_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[31] , 
        \FIC_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[30] , 
        \FIC_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[29] , 
        \FIC_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[28] , 
        \FIC_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[27] , 
        \FIC_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[26] , 
        \FIC_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[25] , 
        \FIC_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[24] , 
        \FIC_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[23] , 
        \FIC_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[22] , 
        \FIC_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[21] , 
        \FIC_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[20] , 
        \FIC_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[19] , 
        \FIC_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[18] , 
        \FIC_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[17] , 
        \FIC_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[16] , 
        \FIC_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[15] , 
        \FIC_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[14] , 
        \FIC_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[13] , 
        \FIC_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[12] , 
        \FIC_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[11] , 
        \FIC_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[10] , 
        \FIC_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[9] , 
        \FIC_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[8] , 
        \FIC_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[7] , 
        \FIC_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[6] , 
        \FIC_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[5] , 
        \FIC_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[4] , 
        \FIC_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[3] , 
        \FIC_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[2] , 
        \FIC_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[1] , 
        \FIC_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[0] , 
        \FIC_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PREADY_net , 
        \FIC_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PSLVERR_net , 
        \FIC_MSS_0/MSS_ADLIB_INST/RCGF_net[9] , 
        \FIC_MSS_0/MSS_ADLIB_INST/RCGF_net[8] , 
        \FIC_MSS_0/MSS_ADLIB_INST/RCGF_net[7] , 
        \FIC_MSS_0/MSS_ADLIB_INST/RCGF_net[6] , 
        \FIC_MSS_0/MSS_ADLIB_INST/RCGF_net[5] , 
        \FIC_MSS_0/MSS_ADLIB_INST/RCGF_net[4] , 
        \FIC_MSS_0/MSS_ADLIB_INST/RCGF_net[3] , 
        \FIC_MSS_0/MSS_ADLIB_INST/RCGF_net[2] , 
        \FIC_MSS_0/MSS_ADLIB_INST/RCGF_net[1] , 
        \FIC_MSS_0/MSS_ADLIB_INST/RCGF_net[0] , 
        \FIC_MSS_0/MSS_ADLIB_INST/RX_CLKPF_net , 
        \FIC_MSS_0/MSS_ADLIB_INST/RX_DVF_net , 
        \FIC_MSS_0/MSS_ADLIB_INST/RX_ERRF_net , 
        \FIC_MSS_0/MSS_ADLIB_INST/RX_EV_net , 
        \FIC_MSS_0/MSS_ADLIB_INST/RXDF_net[7] , 
        \FIC_MSS_0/MSS_ADLIB_INST/RXDF_net[6] , 
        \FIC_MSS_0/MSS_ADLIB_INST/RXDF_net[5] , 
        \FIC_MSS_0/MSS_ADLIB_INST/RXDF_net[4] , 
        \FIC_MSS_0/MSS_ADLIB_INST/RXDF_net[3] , 
        \FIC_MSS_0/MSS_ADLIB_INST/RXDF_net[2] , 
        \FIC_MSS_0/MSS_ADLIB_INST/RXDF_net[1] , 
        \FIC_MSS_0/MSS_ADLIB_INST/RXDF_net[0] , 
        \FIC_MSS_0/MSS_ADLIB_INST/SLEEPHOLDREQ_net , 
        \FIC_MSS_0/MSS_ADLIB_INST/SMBALERT_NI0_net , 
        \FIC_MSS_0/MSS_ADLIB_INST/SMBALERT_NI1_net , 
        \FIC_MSS_0/MSS_ADLIB_INST/SMBSUS_NI0_net , 
        \FIC_MSS_0/MSS_ADLIB_INST/SMBSUS_NI1_net , 
        \FIC_MSS_0/MSS_ADLIB_INST/SPI0_CLK_IN_net , 
        \FIC_MSS_0/MSS_ADLIB_INST/SPI0_SDI_F2H_SCP_net , 
        \FIC_MSS_0/MSS_ADLIB_INST/SPI0_SDO_F2H_SCP_net , 
        \FIC_MSS_0/MSS_ADLIB_INST/SPI0_SS0_F2H_SCP_net , 
        \FIC_MSS_0/MSS_ADLIB_INST/SPI0_SS1_F2H_SCP_net , 
        \FIC_MSS_0/MSS_ADLIB_INST/SPI0_SS2_F2H_SCP_net , 
        \FIC_MSS_0/MSS_ADLIB_INST/SPI0_SS3_F2H_SCP_net , 
        \FIC_MSS_0/MSS_ADLIB_INST/SPI1_CLK_IN_net , 
        \FIC_MSS_0/MSS_ADLIB_INST/SPI1_SDI_F2H_SCP_net , 
        \FIC_MSS_0/MSS_ADLIB_INST/SPI1_SDO_F2H_SCP_net , 
        \FIC_MSS_0/MSS_ADLIB_INST/SPI1_SS0_F2H_SCP_net , 
        \FIC_MSS_0/MSS_ADLIB_INST/SPI1_SS1_F2H_SCP_net , 
        \FIC_MSS_0/MSS_ADLIB_INST/SPI1_SS2_F2H_SCP_net , 
        \FIC_MSS_0/MSS_ADLIB_INST/SPI1_SS3_F2H_SCP_net , 
        \FIC_MSS_0/MSS_ADLIB_INST/TX_CLKPF_net , 
        \FIC_MSS_0/MSS_ADLIB_INST/USER_MSS_GPIO_RESET_N_net , 
        \FIC_MSS_0/MSS_ADLIB_INST/USER_MSS_RESET_N_net , 
        \FIC_MSS_0/MSS_ADLIB_INST/XCLK_FAB_net , 
        \FIC_MSS_0/MSS_ADLIB_INST/CLK_BASE_net , 
        \FIC_MSS_0/MSS_ADLIB_INST/CLK_MDDR_APB_net , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[31] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[30] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[29] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[28] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[27] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[26] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[25] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[24] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[23] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[22] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[21] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[20] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[19] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[18] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[17] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[16] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[15] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[14] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[13] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[12] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[11] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[10] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[9] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[8] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[7] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[6] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[5] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[4] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[3] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[2] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[1] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[0] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_ARBURST_HTRANS1_net[1] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_ARBURST_HTRANS1_net[0] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_ARID_HSEL1_net[3] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_ARID_HSEL1_net[2] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_ARID_HSEL1_net[1] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_ARID_HSEL1_net[0] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_ARLEN_HBURST1_net[3] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_ARLEN_HBURST1_net[2] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_ARLEN_HBURST1_net[1] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_ARLEN_HBURST1_net[0] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_ARLOCK_HMASTLOCK1_net[1] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_ARLOCK_HMASTLOCK1_net[0] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_ARSIZE_HSIZE1_net[1] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_ARSIZE_HSIZE1_net[0] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_ARVALID_HWRITE1_net , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[31] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[30] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[29] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[28] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[27] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[26] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[25] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[24] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[23] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[22] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[21] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[20] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[19] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[18] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[17] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[16] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[15] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[14] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[13] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[12] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[11] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[10] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[9] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[8] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[7] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[6] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[5] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[4] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[3] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[2] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[1] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[0] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_AWBURST_HTRANS0_net[1] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_AWBURST_HTRANS0_net[0] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_AWID_HSEL0_net[3] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_AWID_HSEL0_net[2] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_AWID_HSEL0_net[1] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_AWID_HSEL0_net[0] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_AWLEN_HBURST0_net[3] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_AWLEN_HBURST0_net[2] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_AWLEN_HBURST0_net[1] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_AWLEN_HBURST0_net[0] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_AWLOCK_HMASTLOCK0_net[1] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_AWLOCK_HMASTLOCK0_net[0] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_AWSIZE_HSIZE0_net[1] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_AWSIZE_HSIZE0_net[0] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_AWVALID_HWRITE0_net , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_BREADY_net , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_RMW_AXI_net , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_RREADY_net , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[63] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[62] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[61] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[60] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[59] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[58] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[57] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[56] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[55] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[54] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[53] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[52] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[51] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[50] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[49] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[48] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[47] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[46] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[45] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[44] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[43] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[42] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[41] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[40] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[39] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[38] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[37] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[36] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[35] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[34] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[33] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[32] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[31] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[30] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[29] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[28] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[27] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[26] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[25] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[24] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[23] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[22] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[21] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[20] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[19] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[18] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[17] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[16] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[15] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[14] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[13] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[12] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[11] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[10] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[9] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[8] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[7] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[6] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[5] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[4] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[3] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[2] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[1] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[0] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_WID_HREADY01_net[3] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_WID_HREADY01_net[2] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_WID_HREADY01_net[1] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_WID_HREADY01_net[0] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_WLAST_net , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_WSTRB_net[7] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_WSTRB_net[6] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_WSTRB_net[5] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_WSTRB_net[4] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_WSTRB_net[3] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_WSTRB_net[2] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_WSTRB_net[1] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_WSTRB_net[0] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_WVALID_net , 
        \FIC_MSS_0/MSS_ADLIB_INST/FPGA_MDDR_ARESET_N_net , 
        \FIC_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PADDR_net[10] , 
        \FIC_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PADDR_net[9] , 
        \FIC_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PADDR_net[8] , 
        \FIC_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PADDR_net[7] , 
        \FIC_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PADDR_net[6] , 
        \FIC_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PADDR_net[5] , 
        \FIC_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PADDR_net[4] , 
        \FIC_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PADDR_net[3] , 
        \FIC_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PADDR_net[2] , 
        \FIC_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PENABLE_net , 
        \FIC_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PSEL_net , 
        \FIC_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[15] , 
        \FIC_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[14] , 
        \FIC_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[13] , 
        \FIC_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[12] , 
        \FIC_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[11] , 
        \FIC_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[10] , 
        \FIC_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[9] , 
        \FIC_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[8] , 
        \FIC_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[7] , 
        \FIC_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[6] , 
        \FIC_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[5] , 
        \FIC_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[4] , 
        \FIC_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[3] , 
        \FIC_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[2] , 
        \FIC_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[1] , 
        \FIC_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[0] , 
        \FIC_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWRITE_net , 
        \FIC_MSS_0/MSS_ADLIB_INST/PRESET_N_net , 
        \FIC_MSS_0/MDDR_DQ_11_PAD/YIN , 
        \FIC_MSS_0/MDDR_DQS_1_PAD/U2_N2P , 
        \FIC_MSS_0/MDDR_DQS_1_PAD/YIN , \FIC_MSS_0/MDDR_BA_0_PAD/EOUT , 
        \FIC_MSS_0/MDDR_ADDR_8_PAD/EOUT , 
        \FIC_MSS_0/MDDR_ADDR_13_PAD/EOUT , 
        \FIC_MSS_0/MDDR_ADDR_9_PAD/EOUT , 
        \FIC_MSS_0/MDDR_ADDR_3_PAD/EOUT , 
        \FIC_MSS_0/MDDR_DQ_13_PAD/YIN , \FIC_MSS_0/MDDR_BA_2_PAD/EOUT , 
        \FIC_MSS_0/MDDR_ADDR_6_PAD/EOUT , 
        \FIC_MSS_0/MMUART_0_RXD_PAD/YIN , 
        \FIC_MSS_0/MDDR_DQ_12_PAD/YIN , \FIC_MSS_0/MDDR_DQ_9_PAD/YIN , 
        \FIC_MSS_0/MDDR_ADDR_7_PAD/EOUT , 
        \FIC_MSS_0/MDDR_ADDR_12_PAD/EOUT , 
        \FIC_MSS_0/MDDR_DQ_0_PAD/YIN , \FIC_MSS_0/MDDR_DQ_6_PAD/YIN , 
        \FIC_MSS_0/MDDR_DM_RDQS_0_PAD/YIN , CFG0_GND_INST_NET, 
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_YR , 
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB0_rgbr_net_1 , 
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB1_rgbr_net_1 , 
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB1_rgbl_net_1 , 
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB2_rgbr_net_1 , 
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB2_rgbl_net_1 , 
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB3_rgbr_net_1 , 
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB4_rgbr_net_1 , 
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB5_rgbr_net_1 , 
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB6_rgbr_net_1 , 
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB7_rgbr_net_1 , 
        \FCCC_0/GL1_INST/U0_RGB1_YR , 
        \FCCC_0/GL1_INST/U0_RGB1_RGB0_rgbl_net_1 , 
        \FCCC_0/GL1_INST/U0_RGB1_RGB1_rgbl_net_1 , 
        \FCCC_0/GL1_INST/U0_RGB1_RGB1_rgbr_net_1 , 
        \FCCC_0/GL1_INST/U0_RGB1_RGB2_rgbl_net_1 , 
        \FCCC_0/GL1_INST/U0_RGB1_RGB2_rgbr_net_1 , 
        \FCCC_0/GL1_INST/U0_RGB1_RGB3_rgbl_net_1 , 
        \FCCC_0/GL1_INST/U0_RGB1_RGB4_rgbr_net_1 , 
        \FCCC_0/GL1_INST/U0_RGB1_RGB4_rgbl_net_1 , 
        \FCCC_0/GL1_INST/U0_RGB1_RGB5_rgbr_net_1 , 
        \FCCC_0/GL1_INST/U0_RGB1_RGB5_rgbl_net_1 , 
        \FCCC_0/GL1_INST/U0_RGB1_RGB6_rgbr_net_1 , 
        \FCCC_0/GL1_INST/U0_RGB1_RGB6_rgbl_net_1 , 
        \FCCC_0/GL1_INST/U0_RGB1_RGB7_rgbr_net_1 , 
        \FCCC_0/GL1_INST/U0_RGB1_RGB7_rgbl_net_1 , 
        \FCCC_0/GL1_INST/U0_RGB1_RGB8_rgbl_net_1 , 
        \FCCC_0/GL1_INST/U0_RGB1_RGB8_rgbr_net_1 , 
        \FCCC_0/GL1_INST/U0_RGB1_RGB9_rgbr_net_1 , 
        \FCCC_0/GL1_INST/U0_RGB1_RGB9_rgbl_net_1 , 
        \FCCC_0/GL1_INST/U0_RGB1_RGB10_rgbr_net_1 , 
        \FCCC_0/GL1_INST/U0_RGB1_RGB10_rgbl_net_1 , 
        \FCCC_0/GL1_INST/U0_RGB1_RGB11_rgbr_net_1 , 
        \FCCC_0/GL1_INST/U0_RGB1_RGB11_rgbl_net_1 , 
        \FCCC_0/GL1_INST/U0_RGB1_RGB12_rgbr_net_1 , 
        \FCCC_0/GL1_INST/U0_RGB1_RGB12_rgbl_net_1 , 
        \FCCC_0/GL1_INST/U0_RGB1_RGB13_rgbr_net_1 , 
        \FCCC_0/GL1_INST/U0_RGB1_RGB13_rgbl_net_1 , 
        \FCCC_0/GL1_INST/U0_RGB1_RGB14_rgbr_net_1 , 
        \FCCC_0/GL1_INST/U0_RGB1_RGB14_rgbl_net_1 , 
        \FCCC_0/GL1_INST/U0_RGB1_RGB15_rgbr_net_1 , 
        \FCCC_0/GL1_INST/U0_RGB1_RGB15_rgbl_net_1 , 
        \FCCC_0/GL1_INST/U0_RGB1_RGB16_rgbr_net_1 , 
        \FCCC_0/GL1_INST/U0_RGB1_RGB16_rgbl_net_1 , 
        \FCCC_0/GL1_INST/U0_RGB1_RGB17_rgbr_net_1 , 
        \FCCC_0/GL1_INST/U0_RGB1_RGB17_rgbl_net_1 , 
        \FCCC_0/GL1_INST/U0_RGB1_RGB18_rgbl_net_1 , 
        \FCCC_0/GL1_INST/U0_RGB1_RGB19_rgbl_net_1 , 
        \FCCC_0/GL1_INST/U0_YNn_GSouth , 
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_YNn_GSouth , AFLSDF_VCC, 
        AFLSDF_GND, AFLSDF_INV_0_net_1, AFLSDF_INV_1_net_1, 
        AFLSDF_INV_2_net_1, AFLSDF_INV_3_net_1, AFLSDF_INV_4_net_1, 
        AFLSDF_INV_5_net_1, AFLSDF_INV_6_net_1, AFLSDF_INV_7_net_1, 
        AFLSDF_INV_8_net_1, AFLSDF_INV_9_net_1, AFLSDF_INV_10_net_1, 
        AFLSDF_INV_11_net_1, AFLSDF_INV_12_net_1, AFLSDF_INV_13_net_1, 
        AFLSDF_INV_14_net_1, AFLSDF_INV_15_net_1, AFLSDF_INV_16_net_1, 
        AFLSDF_INV_17_net_1, AFLSDF_INV_18_net_1, AFLSDF_INV_19_net_1, 
        AFLSDF_INV_20_net_1, AFLSDF_INV_21_net_1, AFLSDF_INV_22_net_1, 
        AFLSDF_INV_23_net_1, AFLSDF_INV_24_net_1, AFLSDF_INV_25_net_1, 
        AFLSDF_INV_26_net_1, AFLSDF_INV_27_net_1, AFLSDF_INV_28_net_1, 
        AFLSDF_INV_29_net_1, AFLSDF_INV_30_net_1, AFLSDF_INV_31_net_1, 
        AFLSDF_INV_32_net_1, AFLSDF_INV_33_net_1, AFLSDF_INV_34_net_1, 
        AFLSDF_INV_35_net_1, AFLSDF_INV_36_net_1, AFLSDF_INV_37_net_1, 
        AFLSDF_INV_38_net_1, AFLSDF_INV_39_net_1, AFLSDF_INV_40_net_1, 
        AFLSDF_INV_41_net_1, AFLSDF_INV_42_net_1, AFLSDF_INV_43_net_1, 
        AFLSDF_INV_44_net_1, AFLSDF_INV_45_net_1, AFLSDF_INV_46_net_1, 
        AFLSDF_INV_47_net_1, AFLSDF_INV_48_net_1, AFLSDF_INV_49_net_1, 
        AFLSDF_INV_50_net_1, AFLSDF_INV_51_net_1, AFLSDF_INV_52_net_1, 
        AFLSDF_INV_53_net_1, AFLSDF_INV_54_net_1, AFLSDF_INV_55_net_1, 
        AFLSDF_INV_56_net_1, AFLSDF_INV_57_net_1, AFLSDF_INV_58_net_1, 
        AFLSDF_INV_59_net_1, AFLSDF_INV_60_net_1, AFLSDF_INV_61_net_1, 
        AFLSDF_INV_62_net_1, AFLSDF_INV_63_net_1, AFLSDF_INV_64_net_1, 
        AFLSDF_INV_65_net_1, AFLSDF_INV_66_net_1, AFLSDF_INV_67_net_1, 
        AFLSDF_INV_68_net_1, AFLSDF_INV_69_net_1, AFLSDF_INV_70_net_1, 
        AFLSDF_INV_71_net_1, AFLSDF_INV_72_net_1, AFLSDF_INV_73_net_1, 
        AFLSDF_INV_74_net_1, AFLSDF_INV_75_net_1, AFLSDF_INV_76_net_1, 
        AFLSDF_INV_77_net_1, AFLSDF_INV_78_net_1, AFLSDF_INV_79_net_1, 
        AFLSDF_INV_80_net_1, AFLSDF_INV_81_net_1, AFLSDF_INV_82_net_1, 
        AFLSDF_INV_83_net_1, AFLSDF_INV_84_net_1, AFLSDF_INV_85_net_1, 
        AFLSDF_INV_86_net_1, AFLSDF_INV_87_net_1, AFLSDF_INV_88_net_1, 
        AFLSDF_INV_89_net_1, AFLSDF_INV_90_net_1, AFLSDF_INV_91_net_1, 
        AFLSDF_INV_92_net_1, AFLSDF_INV_93_net_1, AFLSDF_INV_94_net_1, 
        AFLSDF_INV_95_net_1, AFLSDF_INV_96_net_1, AFLSDF_INV_97_net_1, 
        AFLSDF_INV_98_net_1, AFLSDF_INV_99_net_1, AFLSDF_INV_100_net_1, 
        AFLSDF_INV_101_net_1, AFLSDF_INV_102_net_1, 
        AFLSDF_INV_103_net_1, AFLSDF_INV_104_net_1, 
        AFLSDF_INV_105_net_1, AFLSDF_INV_106_net_1, 
        AFLSDF_INV_107_net_1, AFLSDF_INV_108_net_1, 
        AFLSDF_INV_109_net_1, AFLSDF_INV_110_net_1, 
        AFLSDF_INV_111_net_1, AFLSDF_INV_112_net_1, 
        AFLSDF_INV_113_net_1, AFLSDF_INV_114_net_1, 
        AFLSDF_INV_115_net_1, AFLSDF_INV_116_net_1, 
        AFLSDF_INV_117_net_1, AFLSDF_INV_118_net_1, 
        AFLSDF_INV_119_net_1, AFLSDF_INV_120_net_1, 
        AFLSDF_INV_121_net_1, AFLSDF_INV_122_net_1, 
        AFLSDF_INV_123_net_1, AFLSDF_INV_124_net_1, 
        AFLSDF_INV_125_net_1, AFLSDF_INV_126_net_1, 
        AFLSDF_INV_127_net_1, AFLSDF_INV_128_net_1, 
        AFLSDF_INV_129_net_1;
    wire GND_power_net1;
    wire VCC_power_net1;
    assign GND = GND_power_net1;
    assign AFLSDF_GND = GND_power_net1;
    assign VCC = VCC_power_net1;
    assign AFLSDF_VCC = VCC_power_net1;
    
    CFG4 #( .INIT(16'h0F35) )  
        \CoreGPIO_0/CONFIG_reg_o_2_31_am_1_RNO_2[5]  (.A(
        \CoreGPIO_0/CONFIG_reg[0][5] ), .B(
        \CoreGPIO_0/CONFIG_reg[16][5] ), .C(
        \CoreAPB3_0_APBmslave3_PADDR[6] ), .D(
        \CoreAPB3_0_APBmslave3_PADDR[5] ), .Y(
        \CoreGPIO_0/CONFIG_reg_o_2_3_1[5] ));
    CFG2 #( .INIT(4'h7) )  \CoreGPIO_0/edge_both_2_sqmuxa_30_i  (.A(
        \CoreGPIO_0/N_248 ), .B(\CoreGPIO_0/CONFIG_reg[25][3] ), .Y(
        \CoreGPIO_0/N_157 ));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_7_[0]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[0] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB7_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_7__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_204_i ), .ADn(VCC), .SLn(
        VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_7_rs[0] ));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_6_[7]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[7] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB8_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_6__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_202_i ), .ADn(VCC), .SLn(
        VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_6_rs[7] ));
    CFG4 #( .INIT(16'hA9FF) )  
        \CoreGPIO_0/xhdl1.GEN_BITS[28].APB_32.INTR_reg_373_0_o2_0_0[28]  
        (.A(\CoreGPIO_0/CONFIG_reg[28][7] ), .B(
        \CoreGPIO_0/CONFIG_reg[28][6] ), .C(
        \CoreGPIO_0/CONFIG_reg[28][5] ), .D(
        \CoreGPIO_0/CONFIG_reg[28][3] ), .Y(
        \CoreGPIO_0/INTR_reg_373_0_o2_0[28] ));
    CFG2 #( .INIT(4'h4) )  \CoreGPIO_0/PRDATA_0_iv_0_a2_0[28]  (.A(
        \CoreGPIO_0.N_247 ), .B(\CoreGPIO_0/INTR_reg[28] ), .Y(
        \CoreGPIO_0.N_530 ));
    CFG4 #( .INIT(16'hEC00) )  \CoreAPB3_0/u_mux_p_to_b3/PRDATA[23]  (
        .A(\CoreGPIO_0.xhdl1.GEN_BITS[0].APB_32.GPOUT_reg9 ), .B(
        \CoreGPIO_0.N_540 ), .C(
        \CoreGPIO_0.xhdl1.GEN_BITS[23].APB_32.GPOUT_reg[23] ), .D(
        CoreAPB3_0_APBmslave5_PSELx), .Y(
        \FIC_MSS_0_FIC_0_APB_MASTER_PRDATA[23] ));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_2_[4]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[4] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB11_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_2__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_148_i ), .ADn(VCC), .SLn(
        VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_2_rs[4] ));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_3_[6]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[6] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB18_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_3__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_159_i ), .ADn(VCC), .SLn(
        VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_3_rs[6] ));
    IOTRI_OB_EB \FIC_MSS_0/MDDR_RAS_N_PAD/U_IOOUT  (.D(VCC), .E(VCC), 
        .DOUT(), .EOUT(\FIC_MSS_0/MDDR_RAS_N_PAD/EOUT ));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_238_rs_RNIQOHL  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_110_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_238_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_13_rs[6] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_13_[6]_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_131_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_80_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_131_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_131_rs_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_9_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB18_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_4__1_sqmuxa ), .ALn(
        AFLSDF_INV_0_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(GND), 
        .Q(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_9_set_net_1 ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[6].APB_32.GPOUT_reg[6]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[6] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB13_rgbr_net_1 ), .EN(
        \CoreGPIO_0/GPOUT_reg_0_sqmuxa ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB3_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0.xhdl1.GEN_BITS[6].APB_32.GPOUT_reg[6] ));
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_12  (
        .A(\reg_apb_wrp_0/reg16x8_0/mem_1_[1]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_502 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_12_net_1 ));
    CFG3 #( .INIT(8'hF7) )  \FIC_MSS_0/MSS_ADLIB_INST_RNO_6  (.A(
        FIC_MSS_0_FIC_0_APB_MASTER_PSELx), .B(
        \CoreAPB3_0.iPSELS_raw23 ), .C(CoreAPB3_0_APBmslave3_PREADY), 
        .Y(\FIC_MSS_0/FIC_MSS_0_FIC_0_APB_MASTER_PREADY1_i_m_i_0 ));
    CFG3 #( .INIT(8'hDF) )  \CoreGPIO_0/edge_both_2_sqmuxa_12_i_0  (.A(
        \CoreGPIO_0/CONFIG_reg[3][3] ), .B(\CoreGPIO_0/N_253_i ), .C(
        \CoreGPIO_0/N_248 ), .Y(\CoreGPIO_0/edge_both_2_sqmuxa_12_i_1 )
        );
    INV_BA AFLSDF_INV_36 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_70_net_1 ), .Y(
        AFLSDF_INV_36_net_1));
    sdf_IOPAD_BI \FIC_MSS_0/MDDR_DQ_1_PAD/U_IOPAD  (.PAD(MDDR_DQ[1]), 
        .D(\FIC_MSS_0/DRAM_DQ_OUT_net_0[1] ), .E(
        \FIC_MSS_0/DRAM_DQ_OE_net_0[1] ), .Y(
        \FIC_MSS_0/MDDR_DQ_1_PAD_Y ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[25].REG_GEN.CONFIG_reg[25][4]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[4] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB14_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[25]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB4_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[25][4] ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_152  (.A(VCC), 
        .B(VCC), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/MGPIO3A_F2H_GPIN_net ), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/SPI0_SDO_F2H_SCP_net ), .IPC());
    CFG4 #( .INIT(16'hAC0F) )  
        \CoreGPIO_0/CONFIG_reg_o_2_31_am_RNO[4]  (.A(
        \CoreGPIO_0/CONFIG_reg[10][4] ), .B(
        \CoreGPIO_0/CONFIG_reg[26][4] ), .C(
        \CoreGPIO_0/CONFIG_reg_o_2_10_1_1[4] ), .D(
        \CoreAPB3_0_APBmslave3_PADDR[5] ), .Y(
        \CoreGPIO_0/CONFIG_reg_o_2_31_am_RNO[4]_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_4_[1]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[1] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB12_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_4__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_162_i ), .ADn(VCC), .SLn(
        VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_4_rs[1] ));
    CFG2 #( .INIT(4'h8) )  
        \reg_apb_wrp_0/reg16x8_0/mem_14__1_sqmuxa_0_a3  (.A(
        \reg_apb_wrp_0/reg16x8_0/N_503 ), .B(
        \reg_apb_wrp_0/wr_enable_net_1 ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_14__1_sqmuxa ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[3].REG_GEN.CONFIG_reg[3][5]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[5] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB9_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[3]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_YR ), .ADn(VCC), .SLn(
        VCC), .SD(GND), .LAT(GND), .Q(\CoreGPIO_0/CONFIG_reg[3][5] ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_132_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_85_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_132_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_132_rs_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_10_[3]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[3] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB1_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_10__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_197_i ), .ADn(VCC), .SLn(
        VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_10_rs[3] ));
    CFG3 #( .INIT(8'h20) )  
        \CoreGPIO_0/xhdl1.GEN_BITS[29].APB_32.edge_both_RNO[29]  (.A(
        \CoreGPIO_0/CONFIG_reg[29][3] ), .B(
        \CoreAPB3_0_APBmslave3_PWDATA[29] ), .C(
        \CoreGPIO_0/edge_pos[29] ), .Y(\CoreGPIO_0/edge_neg_415[29] ));
    CFG2 #( .INIT(4'h1) )  \reg_apb_wrp_0/rd_enable_RNO  (.A(
        CoreAPB3_0_APBmslave3_PWRITE), .B(\reg_apb_wrp_0/fsm[0]_net_1 )
        , .Y(\reg_apb_wrp_0/N_76 ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_109  (.A(VCC), 
        .B(VCC), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/FAB_XDATAIN_net[1] ), .IPB(), .IPC());
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_105  (.A(VCC), 
        .B(VCC), .C(VCC), .IPA(\FIC_MSS_0/MSS_ADLIB_INST/RCGF_net[5] ), 
        .IPB(\FIC_MSS_0/MSS_ADLIB_INST/FAB_LINESTATE_net[1] ), .IPC());
    CFG3 #( .INIT(8'hF2) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_147  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_2_[3]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_501 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_147_i ));
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_100  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_10_[7]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_491 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_100_net_1 ));
    sdf_IOPAD_TRI \GPIO_OUT_obuf[4]/U0/U_IOPAD  (.PAD(GPIO_OUT[4]), .D(
        \GPIO_OUT_obuf[4]/U0/DOUT ), .E(\GPIO_OUT_obuf[4]/U0/EOUT ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[24].REG_GEN.CONFIG_reg[24][0]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[0] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB16_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[24]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB6_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[24][0] ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[15].REG_GEN.CONFIG_reg[15][1]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[1] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB11_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[15]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB1_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[15][1] ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_120  (.A(VCC), 
        .B(VCC), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/FAB_VBUSVALID_net ), .IPB(), .IPC());
    CFG3 #( .INIT(8'hF2) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_245  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_14_[5]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_503 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_245_i ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_226  (.A(VCC), 
        .B(VCC), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[10] ), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[22] ), .IPC());
    CFG4 #( .INIT(16'hBBFB) )  \CoreGPIO_0/edge_neg_2_sqmuxa_11_i_0  (
        .A(\CoreGPIO_0/N_399 ), .B(\CoreGPIO_0/CONFIG_reg[1][3] ), .C(
        \CoreGPIO_0/INTR_reg21 ), .D(\CoreGPIO_0.N_247 ), .Y(
        \CoreGPIO_0/N_54 ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[15].APB_32.edge_pos[15]  (.D(
        \CoreGPIO_0/edge_pos_219[15] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB10_rgbr_net_1 ), .EN(
        \CoreGPIO_0/edge_pos_2_sqmuxa_7_i_1 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB0_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/edge_neg[15] ));
    CFG4 #( .INIT(16'h8F88) )  \FIC_MSS_0/MSS_ADLIB_INST_RNO_11  (.A(
        \CoreAPB3_0_APBmslave3_PRDATA[5] ), .B(
        CoreAPB3_0_APBmslave3_PSELx), .C(\CoreGPIO_0.N_247 ), .D(
        \FIC_MSS_0/CoreAPB3_0_APBmslave5_PRDATA_m_c_c_0[5] ), .Y(
        \FIC_MSS_0/CoreAPB3_0_APBmslave5_PRDATA_m_0_0[5] ));
    INV_BA AFLSDF_INV_51 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_51_net_1 ), .Y(
        AFLSDF_INV_51_net_1));
    CFG3 #( .INIT(8'hF2) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_251  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_15_[3]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_497 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_251_i ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[23].REG_GEN.CONFIG_reg[23][5]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[5] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB10_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[23]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB0_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[23][5] ));
    INV_BA AFLSDF_INV_90 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_114_net_1 ), .Y(
        AFLSDF_INV_90_net_1));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[8].REG_GEN.CONFIG_reg[8][0]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[0] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB11_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[8]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB1_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[8][0] ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[13].REG_GEN.CONFIG_reg[13][0]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[0] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB14_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[13]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB4_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[13][0] ));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/mem_2__RNIQB2N[6]  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_38_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_150_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_2_rs[6] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_2_[6]_net_1 ));
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_76  (
        .A(\reg_apb_wrp_0/reg16x8_0/mem_9_[4]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_492 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_76_net_1 ));
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_105  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_13_[1]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_500 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_105_net_1 ));
    CFG2 #( .INIT(4'h4) )  \CoreGPIO_0/edge_neg_2_sqmuxa_10_i_a2  (.A(
        \CoreGPIO_0/gpin2[2] ), .B(
        \CoreGPIO_0.xhdl1.GEN_BITS[2].gpin3[2] ), .Y(
        \CoreGPIO_0/N_395 ));
    CFG4 #( .INIT(16'h8000) )  
        \CoreGPIO_0/xhdl1.GEN_BITS[3].REG_GEN.CONFIG_reg[3]2_0_a4_0_a2  
        (.A(\CoreAPB3_0_APBmslave3_PADDR[3] ), .B(
        \CoreAPB3_0_APBmslave3_PADDR[2] ), .C(\CoreGPIO_0/N_604 ), .D(
        \CoreGPIO_0/N_606 ), .Y(\CoreGPIO_0/CONFIG_reg[3]2 ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[12].REG_GEN.CONFIG_reg[12][2]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[2] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB14_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[12]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB4_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[12][2] ));
    CFG3 #( .INIT(8'hFE) )  
        \CoreGPIO_0/xhdl1.GEN_BITS[0].REG_GEN.CONFIG_reg[0]2_0_a4_0_o2  
        (.A(\CoreAPB3_0_APBmslave3_PADDR[2] ), .B(
        \CoreAPB3_0_APBmslave3_PADDR[3] ), .C(
        \CoreAPB3_0_APBmslave3_PADDR[6] ), .Y(\CoreGPIO_0/N_243 ));
    CFG4 #( .INIT(16'h0F35) )  
        \CoreGPIO_0/CONFIG_reg_o_2_31_bm_RNO_1[2]  (.A(
        \CoreGPIO_0/CONFIG_reg[3][2] ), .B(
        \CoreGPIO_0/CONFIG_reg[19][2] ), .C(
        \CoreAPB3_0_APBmslave3_PADDR[6] ), .D(
        \CoreAPB3_0_APBmslave3_PADDR[5] ), .Y(
        \CoreGPIO_0/CONFIG_reg_o_2_25_1_1[2] ));
    CFG3 #( .INIT(8'hF2) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_164  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_4_[3]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_504 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_164_i ));
    IOTRI_OB_EB \GPIO_OUT_obuf[1]/U0/U_IOTRI  (.D(\GPIO_OUT_net_2[1] ), 
        .E(VCC), .DOUT(\GPIO_OUT_obuf[1]/U0/DOUT1 ), .EOUT(
        \GPIO_OUT_obuf[1]/U0/EOUT1 ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[9].REG_GEN.CONFIG_reg[9][1]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[1] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB16_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[9]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB6_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[9][1] ));
    CFG2 #( .INIT(4'h4) )  \CoreGPIO_0/PRDATA_0_iv_0_a2_0[12]  (.A(
        \CoreGPIO_0.N_247 ), .B(\CoreGPIO_0/INTR_reg[12] ), .Y(
        \CoreGPIO_0.N_562 ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_121_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB14_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_6__1_sqmuxa ), .ALn(
        AFLSDF_INV_1_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(GND), 
        .Q(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_121_set_net_1 ));
    CFG4 #( .INIT(16'hECA0) )  \FIC_MSS_0/MSS_ADLIB_INST_RNO_7  (.A(
        \CoreAPB3_0_APBmslave3_PRDATA[0] ), .B(
        CoreAPB3_0_APBmslave5_PSELx), .C(CoreAPB3_0_APBmslave3_PSELx), 
        .D(\CoreGPIO_0.PRDATA_iv_0_0_1[0] ), .Y(
        \FIC_MSS_0/CoreAPB3_0_APBmslave5_PRDATA_m_0_0[0] ));
    CFG4 #( .INIT(16'hEAFA) )  \FIC_MSS_0/MSS_ADLIB_INST_RNO  (.A(
        \FIC_MSS_0/CoreAPB3_0_APBmslave5_PRDATA_m_0_0[0] ), .B(
        \CoreGPIO_0.PRDATA_iv_0_0_0_0[0] ), .C(
        CoreAPB3_0_APBmslave5_PSELx), .D(
        \FIC_MSS_0/CoreAPB3_0_APBmslave5_PRDATA_m_0_1[0] ), .Y(
        \FIC_MSS_0/FIC_MSS_0_FIC_0_APB_MASTER_PRDATA[0] ));
    CFG2 #( .INIT(4'h8) )  \CoreAPB3_0/iPSELS[3]  (.A(
        \CoreAPB3_0.iPSELS_raw23 ), .B(
        FIC_MSS_0_FIC_0_APB_MASTER_PSELx), .Y(
        CoreAPB3_0_APBmslave3_PSELx));
    CFG4 #( .INIT(16'h4657) )  
        \CoreGPIO_0/CONFIG_reg_o_2_31_am_1_1[3]  (.A(
        \CoreAPB3_0_APBmslave3_PADDR[4] ), .B(
        \CoreAPB3_0_APBmslave3_PADDR[3] ), .C(
        \CoreGPIO_0/CONFIG_reg_o_2_31_am_1_1_RNO[3]_net_1 ), .D(
        \CoreGPIO_0/CONFIG_reg_o_2_31_am_1_RNO_0[3]_net_1 ), .Y(
        \CoreGPIO_0/CONFIG_reg_o_2_31_am_1[3] ));
    CFG4 #( .INIT(16'hDC00) )  \FIC_MSS_0/MSS_ADLIB_INST_RNO_21  (.A(
        \CoreGPIO_0.N_247 ), .B(\CoreGPIO_0.N_496 ), .C(
        \CoreGPIO_0.xhdl1.GEN_BITS[3].APB_32.INTR_reg[3] ), .D(
        CoreAPB3_0_APBmslave5_PSELx), .Y(
        \FIC_MSS_0/CoreAPB3_0_APBmslave5_PRDATA_m_d[3] ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[23].APB_32.edge_both[23]  (.D(
        \CoreGPIO_0/N_96_i_0 ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB10_rgbr_net_1 ), .EN(
        \CoreGPIO_0/edge_pos_2_sqmuxa_26_i_1 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB0_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/edge_neg[23] ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_87  (.A(VCC), 
        .B(VCC), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[28] ), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/RXDF_net[3] ), .IPC());
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_268  (.A(VCC), 
        .B(\FCCC_0/GL1_INST/U0_RGB1_YR ), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[28] ), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/CLK_BASE_net ), .IPC());
    IOINFF_BYPASS \FIC_MSS_0/MDDR_DQS_1_PAD/U_IOINFF  (.A(
        \FIC_MSS_0/MDDR_DQS_1_PAD_Y ), .Y(
        \FIC_MSS_0/MDDR_DQS_1_PAD/YIN ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_10  (.A(VCC), 
        .B(\FIC_MSS_0_FIC_0_APB_MASTER_PRDATA[15] ), .C(VCC), .IPA(), 
        .IPB(\FIC_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[15] ), .IPC());
    CFG4 #( .INIT(16'h330A) )  
        \CoreGPIO_0/xhdl1.GEN_BITS[9].APB_32.INTR_reg_126_0[9]  (.A(
        \CoreGPIO_0/INTR_reg[9] ), .B(
        \CoreGPIO_0/INTR_reg_126_0_o2_1[9] ), .C(
        \CoreAPB3_0_APBmslave3_PWDATA[9] ), .D(\CoreGPIO_0/N_248 ), .Y(
        \CoreGPIO_0/INTR_reg_126[9] ));
    CFG4 #( .INIT(16'h7350) )  
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_5[4]  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_14_[4]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/mem_6_[4]_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/N_503 ), .D(
        \reg_apb_wrp_0/reg16x8_0/N_493 ), .Y(
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_5[4]_net_1 ));
    CFG4 #( .INIT(16'h7530) )  
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_1[4]  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_15_[4]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/mem_7_[4]_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/N_498 ), .D(
        \reg_apb_wrp_0/reg16x8_0/N_497 ), .Y(
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_1[4]_net_1 ));
    CFG3 #( .INIT(8'hF2) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_246  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_14_[6]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_503 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_246_i ));
    CFG4 #( .INIT(16'hEFEE) )  
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_8[0]  (.A(
        \reg_apb_wrp_0/reg16x8_0/N_358 ), .B(
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_1[0]_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_5_[0]_net_1 ), .D(
        \reg_apb_wrp_0/reg16x8_0/N_490 ), .Y(
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_8[0]_net_1 ));
    CFG3 #( .INIT(8'hF2) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_238  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_13_[6]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_500 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_238_i ));
    RGB \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1  (.An(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_YNn_GSouth ), .ENn(GND), .YL()
        , .YR(\MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_YR ));
    CFG4 #( .INIT(16'hEFEE) )  
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_9[2]  (.A(
        \reg_apb_wrp_0/reg16x8_0/N_398 ), .B(
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_3[2]_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_1_[2]_net_1 ), .D(
        \reg_apb_wrp_0/reg16x8_0/N_502 ), .Y(
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_9[2]_net_1 ));
    CFG4 #( .INIT(16'h2000) )  
        \reg_apb_wrp_0/reg16x8_0/WRITE_GEN.mem_11__2_i_a2[6]  (.A(
        \CoreAPB3_0_APBmslave3_PADDR[3] ), .B(
        \CoreAPB3_0_APBmslave3_PADDR[2] ), .C(
        \CoreAPB3_0_APBmslave3_PADDR[0] ), .D(
        \CoreAPB3_0_APBmslave3_PADDR[1] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/N_505 ));
    INV_BA AFLSDF_INV_121 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_5_net_1 ), .Y(
        AFLSDF_INV_121_net_1));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_34_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB12_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_2__1_sqmuxa ), .ALn(
        AFLSDF_INV_2_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(GND), 
        .Q(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_34_set_net_1 ));
    CFG4 #( .INIT(16'hEC00) )  \CoreAPB3_0/u_mux_p_to_b3/PRDATA[15]  (
        .A(\CoreGPIO_0.xhdl1.GEN_BITS[0].APB_32.GPOUT_reg9 ), .B(
        \CoreGPIO_0.N_556 ), .C(
        \CoreGPIO_0.xhdl1.GEN_BITS[15].APB_32.GPOUT_reg[15] ), .D(
        CoreAPB3_0_APBmslave5_PSELx), .Y(
        \FIC_MSS_0_FIC_0_APB_MASTER_PRDATA[15] ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_191_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_97_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_191_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_191_rs_net_1 ));
    CFG4 #( .INIT(16'hAA08) )  
        \CoreGPIO_0/xhdl1.GEN_BITS[3].APB_32.edge_neg_51_iv_i_0[3]  (
        .A(\CoreGPIO_0/CONFIG_reg[3][3] ), .B(\CoreGPIO_0/edge_neg[3] )
        , .C(\CoreAPB3_0_APBmslave3_PWDATA[3] ), .D(\CoreGPIO_0/N_686 )
        , .Y(\CoreGPIO_0/edge_neg_51_iv_i_1[3] ));
    IOINFF_BYPASS \GPIO_IN_ibuf[1]/U0/U_IOINFF  (.A(
        \GPIO_IN_ibuf[1]/U0/YIN1 ), .Y(\GPIO_IN_ibuf[1]/U0/YIN ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_219_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_7_net_1 ), .EN(VCC), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_219_i ), .ADn(VCC), .SLn(
        VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_219_rs_net_1 ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[14].REG_GEN.CONFIG_reg[14][3]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[3] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB13_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[14]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB3_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[14][3] ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[27].APB_32.GPOUT_reg[27]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[27] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB10_rgbr_net_1 ), .EN(
        \CoreGPIO_0/GPOUT_reg_0_sqmuxa ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB0_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0.xhdl1.GEN_BITS[27].APB_32.GPOUT_reg[27] ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[12].REG_GEN.CONFIG_reg[12][6]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[6] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB12_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[12]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB2_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[12][6] ));
    INV_BA AFLSDF_INV_62 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_88_net_1 ), .Y(
        AFLSDF_INV_62_net_1));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_16_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB1_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_12__1_sqmuxa ), .ALn(
        AFLSDF_INV_3_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(GND), 
        .Q(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_16_set_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_192_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_33_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_192_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_192_rs_net_1 ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_99  (.A(VCC), 
        .B(VCC), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/GTX_CLKPF_net ), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/RCGF_net[6] ), .IPC());
    CFG4 #( .INIT(16'hA9FF) )  
        \CoreGPIO_0/xhdl1.GEN_BITS[29].APB_32.INTR_reg_386_0_o2_0_0[29]  
        (.A(\CoreGPIO_0/CONFIG_reg[29][7] ), .B(
        \CoreGPIO_0/CONFIG_reg[29][6] ), .C(
        \CoreGPIO_0/CONFIG_reg[29][5] ), .D(
        \CoreGPIO_0/CONFIG_reg[29][3] ), .Y(
        \CoreGPIO_0/INTR_reg_386_0_o2_0[29] ));
    CFG3 #( .INIT(8'hF2) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_214  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_11_[4]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_505 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_214_i ));
    IOIN_IB \GPIO_IN_ibuf[6]/U0/U_IOIN  (.YIN(\GPIO_IN_ibuf[6]/U0/YIN )
        , .E(GND), .Y(\GPIO_IN_c[6] ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_89_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB17_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_11__1_sqmuxa ), .ALn(
        AFLSDF_INV_4_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(GND), 
        .Q(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_89_set_net_1 ));
    CFG4 #( .INIT(16'hA9FF) )  
        \CoreGPIO_0/xhdl1.GEN_BITS[20].APB_32.INTR_reg_269_0_o2_0_0[20]  
        (.A(\CoreGPIO_0/CONFIG_reg[20][7] ), .B(
        \CoreGPIO_0/CONFIG_reg[20][6] ), .C(
        \CoreGPIO_0/CONFIG_reg[20][5] ), .D(
        \CoreGPIO_0/CONFIG_reg[20][3] ), .Y(
        \CoreGPIO_0/INTR_reg_269_0_o2_0[20] ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[13].APB_32.edge_both[13]  (.D(
        \CoreGPIO_0/edge_neg_191[13] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB11_rgbr_net_1 ), .EN(
        \CoreGPIO_0/edge_pos_2_sqmuxa_9_i_1 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB1_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/edge_neg[13] ));
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_71  (
        .A(\reg_apb_wrp_0/reg16x8_0/mem_8_[7]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_499 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_71_net_1 ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[1].APB_32.edge_neg[1]  (.D(
        \CoreGPIO_0/N_121 ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB16_rgbr_net_1 ), .EN(
        \CoreGPIO_0/N_54 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB6_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/edge_neg[1] ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[19].REG_GEN.CONFIG_reg[19][5]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[5] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB9_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[19]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_YR ), .ADn(VCC), .SLn(
        VCC), .SD(GND), .LAT(GND), .Q(\CoreGPIO_0/CONFIG_reg[19][5] ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_75_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB15_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_9__1_sqmuxa ), .ALn(
        AFLSDF_INV_5_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(GND), 
        .Q(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_75_set_net_1 ));
    CFG4 #( .INIT(16'h0008) )  
        \reg_apb_wrp_0/reg16x8_0/WRITE_GEN.mem_12__2_i_a2[6]  (.A(
        \CoreAPB3_0_APBmslave3_PADDR[3] ), .B(
        \CoreAPB3_0_APBmslave3_PADDR[2] ), .C(
        \CoreAPB3_0_APBmslave3_PADDR[0] ), .D(
        \CoreAPB3_0_APBmslave3_PADDR[1] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/N_495 ));
    IOINFF_BYPASS \FIC_MSS_0/MDDR_DM_RDQS_0_PAD/U_IOINFF  (.A(
        \FIC_MSS_0/MDDR_DM_RDQS_0_PAD_Y ), .Y(
        \FIC_MSS_0/MDDR_DM_RDQS_0_PAD/YIN ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[6].REG_GEN.CONFIG_reg[6][3]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[3] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB12_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[6]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB2_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[6][3] ));
    CFG4 #( .INIT(16'h7530) )  
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_0_7[5]  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_10_[5]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/mem_2_[5]_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/N_501 ), .D(
        \reg_apb_wrp_0/reg16x8_0/N_491 ), .Y(
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_0_7[5]_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_119_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB8_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_14__1_sqmuxa ), .ALn(
        AFLSDF_INV_6_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(GND), 
        .Q(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_119_set_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_10_[5]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[5] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB11_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_10__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_201_i ), .ADn(VCC), .SLn(
        VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_10_rs[5] ));
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_114  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_14_[2]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_503 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_114_net_1 ));
    CFG4 #( .INIT(16'h2000) )  
        \CoreGPIO_0/xhdl1.GEN_BITS[2].REG_GEN.CONFIG_reg[2]2_0_a4_0_a2  
        (.A(\CoreAPB3_0_APBmslave3_PADDR[3] ), .B(
        \CoreAPB3_0_APBmslave3_PADDR[2] ), .C(\CoreGPIO_0/N_604 ), .D(
        \CoreGPIO_0/N_606 ), .Y(\CoreGPIO_0/CONFIG_reg[2]2 ));
    CFG3 #( .INIT(8'hDF) )  \CoreGPIO_0/edge_both_2_sqmuxa_22_i_0_0  (
        .A(\CoreGPIO_0/CONFIG_reg[6][3] ), .B(\CoreGPIO_0/N_252_i ), 
        .C(\CoreGPIO_0/N_248 ), .Y(\CoreGPIO_0/N_78 ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[8].APB_32.edge_both[8]  (.D(
        \CoreGPIO_0/edge_neg_121[8] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB9_rgbr_net_1 ), .EN(
        \CoreGPIO_0/edge_neg_2_sqmuxa_4_i_1 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_YR ), .ADn(VCC), .SLn(
        VCC), .SD(GND), .LAT(GND), .Q(\CoreGPIO_0/edge_pos[8] ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[17].APB_32.edge_both[17]  (.D(
        \CoreGPIO_0/edge_neg_247[17] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB14_rgbr_net_1 ), .EN(
        \CoreGPIO_0/edge_pos_2_sqmuxa_30_i_1 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB4_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/edge_neg[17] ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[21].REG_GEN.CONFIG_reg[21][7]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[7] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB13_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[21]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB3_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[21][7] ));
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_127  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_7_[1]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_498 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_127_net_1 ));
    CFG3 #( .INIT(8'hF2) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_225  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_8_[3]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_499 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_225_i ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_26  (.A(GND), 
        .B(VCC), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[2] ), .IPB(), .IPC());
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_224  (.A(VCC), 
        .B(VCC), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[8] ), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[20] ), .IPC());
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[1].REG_GEN.CONFIG_reg[1][0]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[0] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB16_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[1]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB6_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[1][0] ));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_2_[2]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[2] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB12_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_2__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_146_i ), .ADn(VCC), .SLn(
        VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_2_rs[2] ));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_10_[4]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[4] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB9_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_10__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_199_i ), .ADn(VCC), .SLn(
        VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_10_rs[4] ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[5].REG_GEN.CONFIG_reg[5][3]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[3] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB13_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[5]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB3_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[5][3] ));
    GB \FCCC_0/GL1_INST  (.An(AFLSDF_INV_7_net_1), .ENn(GND), .YNn(
        \FCCC_0/GL1_INST/U0_YNn ), .YSn(
        \FCCC_0/GL1_INST/U0_YNn_GSouth ));
    CFG4 #( .INIT(16'h2000) )  \CoreAPB3_0/iPSELS[5]  (.A(
        FIC_MSS_0_FIC_0_APB_MASTER_PSELx), .B(
        \FIC_MSS_0_FIC_0_APB_MASTER_PADDR[31] ), .C(
        \FIC_MSS_0_FIC_0_APB_MASTER_PADDR[28] ), .D(
        \CoreAPB3_0/iPSELS_1[5] ), .Y(CoreAPB3_0_APBmslave5_PSELx));
    INV_BA AFLSDF_INV_9 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_28_net_1 ), .Y(
        AFLSDF_INV_9_net_1));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_45_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB16_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_1__1_sqmuxa ), .ALn(
        AFLSDF_INV_8_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(GND), 
        .Q(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_45_set_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_1_[0]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[0] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB14_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_1__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_136_i ), .ADn(VCC), .SLn(
        VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_1_rs[0] ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_262  (.A(VCC), 
        .B(VCC), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[10] ), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[22] ), .IPC());
    SLE \reg_apb_wrp_0/reg16x8_0/mem_9_[6]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[6] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB16_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_9__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_187_i ), .ADn(VCC), .SLn(
        VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_9_rs[6] ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_64  (.A(GND), 
        .B(VCC), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[25] ), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PREADY_net ), .IPC());
    CFG4 #( .INIT(16'h0040) )  
        \reg_apb_wrp_0/reg16x8_0/WRITE_GEN.mem_5__2_i_0_0_a2[5]  (.A(
        \CoreAPB3_0_APBmslave3_PADDR[3] ), .B(
        \CoreAPB3_0_APBmslave3_PADDR[2] ), .C(
        \CoreAPB3_0_APBmslave3_PADDR[0] ), .D(
        \CoreAPB3_0_APBmslave3_PADDR[1] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/N_490 ));
    CFG4 #( .INIT(16'h7530) )  
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_0_4[5]  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_12_[5]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/mem_4_[5]_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/N_504 ), .D(
        \reg_apb_wrp_0/reg16x8_0/N_495 ), .Y(
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_0_4[5]_net_1 ));
    CFG2 #( .INIT(4'h8) )  
        \reg_apb_wrp_0/reg16x8_0/mem_12__1_sqmuxa_0_a3  (.A(
        \reg_apb_wrp_0/reg16x8_0/N_495 ), .B(
        \reg_apb_wrp_0/wr_enable_net_1 ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_12__1_sqmuxa ));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/mem_3__RNISIGN[7]  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_55_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_160_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_3_rs[7] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_3_[7]_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_3_[3]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[3] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB17_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_3__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_155_i ), .ADn(VCC), .SLn(
        VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_3_rs[3] ));
    CFG3 #( .INIT(8'hF2) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_226  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_12_[2]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_495 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_226_i ));
    CFG3 #( .INIT(8'hB8) )  
        \CoreGPIO_0/xhdl1.GEN_BITS[3].REG_INT.un34_intr_1  (.A(
        \CoreGPIO_0/edge_neg[3] ), .B(\CoreGPIO_0/CONFIG_reg[3][5] ), 
        .C(\CoreGPIO_0/edge_pos[3] ), .Y(\CoreGPIO_0/N_4549 ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[13].REG_GEN.CONFIG_reg[13][3]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[3] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB13_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[13]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB3_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[13][3] ));
    CFG4 #( .INIT(16'h0F35) )  
        \CoreGPIO_0/CONFIG_reg_o_2_31_bm_1_RNO_2[1]  (.A(
        \CoreGPIO_0.xhdl1.GEN_BITS[1].REG_GEN.CONFIG_reg[1][1] ), .B(
        \CoreGPIO_0/CONFIG_reg[17][1] ), .C(
        \CoreAPB3_0_APBmslave3_PADDR[6] ), .D(
        \CoreAPB3_0_APBmslave3_PADDR[5] ), .Y(
        \CoreGPIO_0/CONFIG_reg_o_2_18_1[1] ));
    CFG4 #( .INIT(16'h7350) )  
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_5[3]  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_14_[3]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/mem_6_[3]_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/N_503 ), .D(
        \reg_apb_wrp_0/reg16x8_0/N_493 ), .Y(
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_5[3]_net_1 ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_167  (.A(VCC), 
        .B(VCC), .C(VCC), .IPA(), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/MMUART1_RTS_F2H_SCP_net ), .IPC());
    CFG2 #( .INIT(4'h4) )  \CoreGPIO_0/PRDATA_0_iv_0_a2_0[9]  (.A(
        \CoreGPIO_0.N_247 ), .B(\CoreGPIO_0/INTR_reg[9] ), .Y(
        \CoreGPIO_0.N_568 ));
    CFG2 #( .INIT(4'h7) )  \CoreGPIO_0/edge_both_2_sqmuxa_21_i  (.A(
        \CoreGPIO_0/N_248 ), .B(\CoreGPIO_0/CONFIG_reg[7][3] ), .Y(
        \CoreGPIO_0/edge_pos_2_sqmuxa_1_i_1 ));
    CFG4 #( .INIT(16'hF2F3) )  
        \CoreGPIO_0/xhdl1.GEN_BITS[25].APB_32.INTR_reg_334_0_o2_1_0[25]  
        (.A(\CoreGPIO_0/CONFIG_reg[25][6] ), .B(
        \CoreGPIO_0/edge_neg[25] ), .C(
        \CoreGPIO_0/INTR_reg_334_0_o2_0[25] ), .D(
        \CoreGPIO_0/CONFIG_reg[25][5] ), .Y(
        \CoreGPIO_0/INTR_reg_334_0_o2_1[25] ));
    CFG4 #( .INIT(16'h8000) )  
        \CoreGPIO_0/xhdl1.GEN_BITS[31].REG_GEN.CONFIG_reg[31]2_0_a4_0_a2  
        (.A(\CoreAPB3_0_APBmslave3_PADDR[3] ), .B(
        \CoreAPB3_0_APBmslave3_PADDR[2] ), .C(\CoreGPIO_0/N_598 ), .D(
        \CoreGPIO_0/N_605 ), .Y(\CoreGPIO_0/CONFIG_reg[31]2 ));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_40_set_RNIQICR  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_40_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_176_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_5_rs[2] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_5_[2]_net_1 ));
    CFG2 #( .INIT(4'h8) )  
        \reg_apb_wrp_0/reg16x8_0/mem_4__1_sqmuxa_0_a3  (.A(
        \reg_apb_wrp_0/reg16x8_0/N_504 ), .B(
        \reg_apb_wrp_0/wr_enable_net_1 ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_4__1_sqmuxa ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[15].REG_GEN.CONFIG_reg[15][6]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[6] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB10_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[15]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB0_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[15][6] ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[11].REG_GEN.CONFIG_reg[11][5]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[5] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB9_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[11]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_YR ), .ADn(VCC), .SLn(
        VCC), .SD(GND), .LAT(GND), .Q(\CoreGPIO_0/CONFIG_reg[11][5] ));
    IOENFF_BYPASS \GPIO_OUT_obuf[5]/U0/U_IOENFF  (.A(
        \GPIO_OUT_obuf[5]/U0/EOUT1 ), .Y(\GPIO_OUT_obuf[5]/U0/EOUT ));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_47_set_RNIO6TL  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_47_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_141_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_1_rs[5] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_1_[5]_net_1 ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_61  (.A(GND), 
        .B(VCC), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[22] ), .IPB(), .IPC()
        );
    SLE \reg_apb_wrp_0/reg16x8_0/mem_0_[1]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[1] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB2_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_0__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_128_i ), .ADn(VCC), .SLn(
        VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_0_rs[1] ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_160_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_55_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_160_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_160_rs_net_1 ));
    CFG4 #( .INIT(16'hEFEE) )  
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_8[6]  (.A(
        \reg_apb_wrp_0/reg16x8_0/N_450 ), .B(
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_1[6]_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_5_[6]_net_1 ), .D(
        \reg_apb_wrp_0/reg16x8_0/N_490 ), .Y(
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_8[6]_net_1 ));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_4_set_RNI519S  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_4_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_163_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_4_rs[2] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_4_[2]_net_1 ));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/mem_2__RNIJLTN[2]  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_30_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_146_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_2_rs[2] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_2_[2]_net_1 ));
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_66  (
        .A(\reg_apb_wrp_0/reg16x8_0/mem_8_[3]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_499 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_66_net_1 ));
    IOBI_IB_OB_EB \FIC_MSS_0/MDDR_DQ_3_PAD/U_IOBI  (.D(VCC), .E(VCC), 
        .YIN(\FIC_MSS_0/MDDR_DQ_3_PAD/YIN ), .DOUT(), .EOUT(), .Y());
    CFG4 #( .INIT(16'h330A) )  
        \CoreGPIO_0/xhdl1.GEN_BITS[29].APB_32.INTR_reg_386_0[29]  (.A(
        \CoreGPIO_0/INTR_reg[29] ), .B(
        \CoreGPIO_0/INTR_reg_386_0_o2_1[29] ), .C(
        \CoreAPB3_0_APBmslave3_PWDATA[29] ), .D(\CoreGPIO_0/N_248 ), 
        .Y(\CoreGPIO_0/INTR_reg_386[29] ));
    CFG4 #( .INIT(16'hB383) )  \CoreGPIO_0/CONFIG_reg_o_2_31_am[3]  (
        .A(\CoreGPIO_0/CONFIG_reg_o_2_31_am_RNO[3]_net_1 ), .B(
        \CoreGPIO_0/CONFIG_reg_o_2_31_am_1[3] ), .C(
        \CoreAPB3_0_APBmslave3_PADDR[3] ), .D(
        \CoreGPIO_0/CONFIG_reg_o_2_31_am_RNO_0[3]_net_1 ), .Y(
        \CONFIG_reg_o_2_31_am[3] ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_136  (.A(VCC), 
        .B(VCC), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/SMBSUS_NI0_net ), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/F_DMAREADY_net[0] ), .IPC());
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_88  (.A(VCC), 
        .B(VCC), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[29] ), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/RXDF_net[4] ), .IPC());
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_79  (
        .A(\reg_apb_wrp_0/reg16x8_0/mem_9_[7]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_492 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_79_net_1 ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[7].APB_32.edge_both[7]  (.D(
        \CoreGPIO_0/N_83_i_0 ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB10_rgbr_net_1 ), .EN(
        \CoreGPIO_0/edge_pos_2_sqmuxa_1_i_1 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB0_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/edge_pos[7] ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[13].APB_32.INTR_reg[13]  (.D(
        \CoreGPIO_0/INTR_reg_178[13] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB11_rgbr_net_1 ), .EN(VCC), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB1_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/INTR_reg[13] ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[31].REG_GEN.CONFIG_reg[31][5]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[5] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB10_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[31]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB0_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[31][5] ));
    CFG4 #( .INIT(16'h4657) )  
        \CoreGPIO_0/CONFIG_reg_o_2_31_bm_1_1[3]  (.A(
        \CoreAPB3_0_APBmslave3_PADDR[4] ), .B(
        \CoreAPB3_0_APBmslave3_PADDR[3] ), .C(
        \CoreGPIO_0/CONFIG_reg_o_2_31_bm_1_1_RNO[3]_net_1 ), .D(
        \CoreGPIO_0/CONFIG_reg_o_2_31_bm_1_RNO_0[3]_net_1 ), .Y(
        \CoreGPIO_0/CONFIG_reg_o_2_31_bm_1[3] ));
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_26  (
        .A(\reg_apb_wrp_0/reg16x8_0/mem_2_[0]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_501 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_26_net_1 ));
    CFG3 #( .INIT(8'h20) )  
        \CoreGPIO_0/xhdl1.GEN_BITS[27].APB_32.edge_both_RNO[27]  (.A(
        \CoreGPIO_0/CONFIG_reg[27][3] ), .B(
        \CoreAPB3_0_APBmslave3_PWDATA[27] ), .C(
        \CoreGPIO_0/edge_neg[27] ), .Y(\CoreGPIO_0/N_5912_i_0 ));
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_84  (
        .A(\reg_apb_wrp_0/reg16x8_0/mem_0_[3]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_496 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_84_net_1 ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[20].APB_32.GPOUT_reg[20]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[20] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB13_rgbr_net_1 ), .EN(
        \CoreGPIO_0/GPOUT_reg_0_sqmuxa ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB3_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0.xhdl1.GEN_BITS[20].APB_32.GPOUT_reg[20] ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_73  (.A(VCC), 
        .B(VCC), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[7] ), .IPB(), 
        .IPC());
    CFG3 #( .INIT(8'hF2) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_194  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_6_[3]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_493 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_194_i ));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_211_rs_RNI25BI  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_90_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_211_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_11_rs[2] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_11_[2]_net_1 ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[8].APB_32.GPOUT_reg[8]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[8] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB9_rgbr_net_1 ), .EN(
        \CoreGPIO_0/GPOUT_reg_0_sqmuxa ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_YR ), .ADn(VCC), .SLn(
        VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0.xhdl1.GEN_BITS[8].APB_32.GPOUT_reg[8] ));
    CFG4 #( .INIT(16'hAC0F) )  
        \CoreGPIO_0/CONFIG_reg_o_2_31_bm_RNO[4]  (.A(
        \CoreGPIO_0/CONFIG_reg[11][4] ), .B(
        \CoreGPIO_0/CONFIG_reg[27][4] ), .C(
        \CoreGPIO_0/CONFIG_reg_o_2_25_1_1[4] ), .D(
        \CoreAPB3_0_APBmslave3_PADDR[5] ), .Y(
        \CoreGPIO_0/CONFIG_reg_o_2_31_bm_RNO[4]_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_159_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_83_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_159_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_159_rs_net_1 ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[6].REG_GEN.CONFIG_reg[6][6]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[6] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB12_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[6]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB2_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[6][6] ));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_15_[1]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[1] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB5_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_15__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_249_i ), .ADn(VCC), .SLn(
        VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_15_rs[1] ));
    IOINFF_BYPASS \FIC_MSS_0/MDDR_DQ_11_PAD/U_IOINFF  (.A(
        \FIC_MSS_0/MDDR_DQ_11_PAD_Y ), .Y(
        \FIC_MSS_0/MDDR_DQ_11_PAD/YIN ));
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_94  (
        .A(\reg_apb_wrp_0/reg16x8_0/mem_11_[6]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_505 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_94_net_1 ));
    CFG4 #( .INIT(16'hEFEE) )  
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_9[7]  (.A(
        \reg_apb_wrp_0/reg16x8_0/N_478 ), .B(
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_3[7]_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_1_[7]_net_1 ), .D(
        \reg_apb_wrp_0/reg16x8_0/N_502 ), .Y(
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_9[7]_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/data_out[7]  (.D(
        \reg_apb_wrp_0/reg16x8_0/temp_data[7]_net_1 ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB12_rgbr_net_1 ), .EN(VCC), .ALn(
        VCC), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreAPB3_0_APBmslave3_PRDATA[7] ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_37  (.A(GND), 
        .B(VCC), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[20] ), .IPB(), .IPC());
    CFG2 #( .INIT(4'h2) )  \CoreGPIO_0/edge_pos_2_sqmuxa_i_a2  (.A(
        \CoreGPIO_0/gpin2[0] ), .B(
        \CoreGPIO_0.xhdl1.GEN_BITS[0].gpin3[0] ), .Y(
        \CoreGPIO_0/N_402 ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[19].REG_GEN.CONFIG_reg[19][4]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[4] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB10_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[19]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB0_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[19][4] ));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_15_[7]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[7] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB3_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_15__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_252_i ), .ADn(VCC), .SLn(
        VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_15_rs[7] ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[15].APB_32.INTR_reg[15]  (.D(
        \CoreGPIO_0/INTR_reg_204[15] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB9_rgbr_net_1 ), .EN(VCC), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_YR ), .ADn(VCC), .SLn(
        VCC), .SD(GND), .LAT(GND), .Q(\CoreGPIO_0/INTR_reg[15] ));
    sdf_IOPAD_TRI \GPIO_OUT_obuf[1]/U0/U_IOPAD  (.PAD(GPIO_OUT[1]), .D(
        \GPIO_OUT_obuf[1]/U0/DOUT ), .E(\GPIO_OUT_obuf[1]/U0/EOUT ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_231  (.A(VCC), 
        .B(VCC), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[29] ), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[41] ), .IPC());
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[5].REG_GEN.CONFIG_reg[5][6]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[6] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB13_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[5]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB3_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[5][6] ));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_236_rs_RNITBIQ  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_108_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_236_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_13_rs[4] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_13_[4]_net_1 ));
    CFG2 #( .INIT(4'h4) )  \CoreGPIO_0/PRDATA_0_iv_0_a2_0[30]  (.A(
        \CoreGPIO_0.N_247 ), .B(\CoreGPIO_0/INTR_reg[30] ), .Y(
        \CoreGPIO_0.N_526 ));
    CFG2 #( .INIT(4'h4) )  \CoreGPIO_0/PRDATA_0_iv_0_a2_0[15]  (.A(
        \CoreGPIO_0.N_247 ), .B(\CoreGPIO_0/INTR_reg[15] ), .Y(
        \CoreGPIO_0.N_556 ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_133  (.A(GND), 
        .B(VCC), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[15] ), .IPB(), 
        .IPC());
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[6].APB_32.edge_both[6]  (.D(
        \CoreGPIO_0/N_22_i_0 ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB12_rgbr_net_1 ), .EN(
        \CoreGPIO_0/N_78 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB2_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/edge_both[6] ));
    INV_BA AFLSDF_INV_13 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_108_net_1 ), .Y(
        AFLSDF_INV_13_net_1));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[28].REG_GEN.CONFIG_reg[28][7]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[7] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB12_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[28]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB2_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[28][7] ));
    CFG2 #( .INIT(4'h2) )  
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_a3_3[3]  (.A(
        \reg_apb_wrp_0/reg16x8_0/N_500 ), .B(
        \reg_apb_wrp_0/reg16x8_0/mem_13_[3]_net_1 ), .Y(
        \reg_apb_wrp_0/reg16x8_0/N_406 ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[13].REG_GEN.CONFIG_reg[13][4]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[4] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB14_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[13]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB4_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[13][4] ));
    CFG4 #( .INIT(16'hAC0F) )  
        \CoreGPIO_0/CONFIG_reg_o_2_31_bm_1_1_RNO[3]  (.A(
        \CoreGPIO_0/CONFIG_reg[13][3] ), .B(
        \CoreGPIO_0/CONFIG_reg[29][3] ), .C(
        \CoreGPIO_0/CONFIG_reg_o_2_21_1[3] ), .D(
        \CoreAPB3_0_APBmslave3_PADDR[5] ), .Y(
        \CoreGPIO_0/CONFIG_reg_o_2_31_bm_1_1_RNO[3]_net_1 ));
    CFG4 #( .INIT(16'hAC0F) )  
        \CoreGPIO_0/CONFIG_reg_o_2_31_am_1_1_RNO[0]  (.A(
        \CoreGPIO_0/CONFIG_reg[12][0] ), .B(
        \CoreGPIO_0/CONFIG_reg[28][0] ), .C(
        \CoreGPIO_0/CONFIG_reg_o_2_6_1[0] ), .D(
        \CoreAPB3_0_APBmslave3_PADDR[5] ), .Y(
        \CoreGPIO_0/CONFIG_reg_o_2_31_am_1_1_RNO[0]_net_1 ));
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_50  (
        .A(\reg_apb_wrp_0/reg16x8_0/mem_3_[4]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_494 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_50_net_1 ));
    sdf_IOPAD_BI \FIC_MSS_0/MDDR_DQ_4_PAD/U_IOPAD  (.PAD(MDDR_DQ[4]), 
        .D(\FIC_MSS_0/DRAM_DQ_OUT_net_0[4] ), .E(
        \FIC_MSS_0/DRAM_DQ_OE_net_0[4] ), .Y(
        \FIC_MSS_0/MDDR_DQ_4_PAD_Y ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_192  (.A(GND), 
        .B(VCC), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/F_AWID_HSEL0_net[0] ), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[8] ), .IPC(
        \FIC_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[20] ));
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_61  (
        .A(\reg_apb_wrp_0/reg16x8_0/mem_15_[3]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_497 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_61_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_173_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_71_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_173_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_173_rs_net_1 ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[18].REG_GEN.CONFIG_reg[18][2]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[2] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB16_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[18]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB6_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[18][2] ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[23].REG_GEN.CONFIG_reg[23][7]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[7] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB10_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[23]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB0_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[23][7] ));
    CFG3 #( .INIT(8'h01) )  \reg_apb_wrp_0/reg16x8_0/temp_data_RNO[7]  
        (.A(\reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_8[7]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_13[7]_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_9[7]_net_1 ), .Y(
        \reg_apb_wrp_0/reg16x8_0/N_86_i_0 ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[3].REG_GEN.CONFIG_reg[3][0]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[0] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB9_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[3]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_YR ), .ADn(VCC), .SLn(
        VCC), .SD(GND), .LAT(GND), .Q(\CoreGPIO_0/CONFIG_reg[3][0] ));
    CFG4 #( .INIT(16'h330A) )  
        \CoreGPIO_0/xhdl1.GEN_BITS[30].APB_32.INTR_reg_399_0[30]  (.A(
        \CoreGPIO_0/INTR_reg[30] ), .B(
        \CoreGPIO_0/INTR_reg_399_0_o2_1[30] ), .C(
        \CoreAPB3_0_APBmslave3_PWDATA[30] ), .D(\CoreGPIO_0/N_248 ), 
        .Y(\CoreGPIO_0/INTR_reg_399[30] ));
    CFG4 #( .INIT(16'hAC0F) )  
        \CoreGPIO_0/CONFIG_reg_o_2_31_am_RNO_0[7]  (.A(
        \CoreGPIO_0/CONFIG_reg[14][7] ), .B(
        \CoreGPIO_0/CONFIG_reg[30][7] ), .C(
        \CoreGPIO_0/CONFIG_reg_o_2_13_1_1[7] ), .D(
        \CoreAPB3_0_APBmslave3_PADDR[5] ), .Y(
        \CoreGPIO_0/CONFIG_reg_o_2_31_am_RNO_0[7]_net_1 ));
    CFG4 #( .INIT(16'h0F35) )  
        \CoreGPIO_0/CONFIG_reg_o_2_31_bm_RNO_1[0]  (.A(
        \CoreGPIO_0/CONFIG_reg[3][0] ), .B(
        \CoreGPIO_0/CONFIG_reg[19][0] ), .C(
        \CoreAPB3_0_APBmslave3_PADDR[6] ), .D(
        \CoreAPB3_0_APBmslave3_PADDR[5] ), .Y(
        \CoreGPIO_0/CONFIG_reg_o_2_25_1_1[0] ));
    CFG3 #( .INIT(8'hF2) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_254  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_15_[5]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_497 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_254_i ));
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_21  (
        .A(\reg_apb_wrp_0/reg16x8_0/mem_12_[5]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_495 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_21_net_1 ));
    CFG4 #( .INIT(16'hAC0F) )  
        \CoreGPIO_0/CONFIG_reg_o_2_31_bm_RNO_0[4]  (.A(
        \CoreGPIO_0/CONFIG_reg[15][4] ), .B(
        \CoreGPIO_0/CONFIG_reg[31][4] ), .C(
        \CoreGPIO_0/CONFIG_reg_o_2_28_1_1[4] ), .D(
        \CoreAPB3_0_APBmslave3_PADDR[5] ), .Y(
        \CoreGPIO_0/CONFIG_reg_o_2_31_bm_RNO_0[4]_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_5_[0]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[0] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB12_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_5__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_172_i ), .ADn(VCC), .SLn(
        VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_5_rs[0] ));
    CFG4 #( .INIT(16'h330A) )  
        \CoreGPIO_0/xhdl1.GEN_BITS[27].APB_32.INTR_reg_360_0[27]  (.A(
        \CoreGPIO_0/INTR_reg[27] ), .B(
        \CoreGPIO_0/INTR_reg_360_0_o2_1[27] ), .C(
        \CoreAPB3_0_APBmslave3_PWDATA[27] ), .D(\CoreGPIO_0/N_248 ), 
        .Y(\CoreGPIO_0/INTR_reg_360[27] ));
    INV_BA AFLSDF_INV_16 (.A(\MSS_RESET_N_F2M_ibuf/U0/YIN1 ), .Y(
        AFLSDF_INV_16_net_1));
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_75  (
        .A(\reg_apb_wrp_0/reg16x8_0/mem_9_[3]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_492 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_75_net_1 ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_54  (.A(GND), 
        .B(GND), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[8] ), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[15] ), .IPC());
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[21].APB_32.INTR_reg[21]  (.D(
        \CoreGPIO_0/INTR_reg_282[21] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB13_rgbr_net_1 ), .EN(VCC), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB3_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/INTR_reg[21] ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[13].REG_GEN.CONFIG_reg[13][6]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[6] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB13_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[13]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB3_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[13][6] ));
    IOINFF_BYPASS \FIC_MSS_0/MDDR_DQS_0_PAD/U_IOINFF  (.A(
        \FIC_MSS_0/MDDR_DQS_0_PAD_Y ), .Y(
        \FIC_MSS_0/MDDR_DQS_0_PAD/YIN ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[8].REG_GEN.CONFIG_reg[8][3]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[3] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB9_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[8]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_YR ), .ADn(VCC), .SLn(
        VCC), .SD(GND), .LAT(GND), .Q(\CoreGPIO_0/CONFIG_reg[8][3] ));
    INV_BA AFLSDF_INV_25 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_109_net_1 ), .Y(
        AFLSDF_INV_25_net_1));
    CFG3 #( .INIT(8'hF2) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_154  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_3_[2]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_494 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_154_i ));
    CFG4 #( .INIT(16'hEFEE) )  
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_10[0]  (.A(
        \reg_apb_wrp_0/reg16x8_0/N_360 ), .B(
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_5[0]_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_4_[0]_net_1 ), .D(
        \reg_apb_wrp_0/reg16x8_0/N_504 ), .Y(
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_10[0]_net_1 ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[5].APB_32.INTR_reg[5]  (.D(
        \CoreGPIO_0/INTR_reg_74[5] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB10_rgbr_net_1 ), .EN(VCC), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB0_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0.xhdl1.GEN_BITS[5].APB_32.INTR_reg[5] ));
    INV_BA AFLSDF_INV_85 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_105_net_1 ), .Y(
        AFLSDF_INV_85_net_1));
    CFG4 #( .INIT(16'hAA08) )  
        \CoreGPIO_0/xhdl1.GEN_BITS[2].APB_32.edge_both_37_iv_i_0[2]  (
        .A(\CoreGPIO_0/CONFIG_reg[2][3] ), .B(
        \CoreGPIO_0/edge_both[2] ), .C(
        \CoreAPB3_0_APBmslave3_PWDATA[2] ), .D(\CoreGPIO_0/N_144_i ), 
        .Y(\CoreGPIO_0/N_93 ));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_14_[0]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[0] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB6_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_14__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_240_i ), .ADn(VCC), .SLn(
        VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_14_rs[0] ));
    IOTRI_OB_EB \FIC_MSS_0/MDDR_ADDR_4_PAD/U_IOOUT  (.D(VCC), .E(VCC), 
        .DOUT(), .EOUT(\FIC_MSS_0/MDDR_ADDR_4_PAD/EOUT ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_171  (.A(VCC), 
        .B(VCC), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/MMUART1_DCD_F2H_SCP_net ), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/MGPIO17B_F2H_GPIN_net ), .IPC());
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_28_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB1_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_2__1_sqmuxa ), .ALn(
        AFLSDF_INV_9_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(GND), 
        .Q(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_28_set_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_12_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB14_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_1__1_sqmuxa ), .ALn(
        AFLSDF_INV_10_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(GND)
        , .Q(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_12_set_net_1 ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[26].REG_GEN.CONFIG_reg[26][5]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[5] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB17_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[26]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB7_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[26][5] ));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_129_rs_RNIPFDM  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_82_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_129_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_0_rs[2] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_0_[2]_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_9_[3]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[3] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB15_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_9__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_181_i ), .ADn(VCC), .SLn(
        VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_9_rs[3] ));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/mem_10__RNIDMMI[0]  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_97_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_191_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_10_rs[0] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_10_[0]_net_1 ));
    CFG4 #( .INIT(16'hAA08) )  
        \CoreGPIO_0/xhdl1.GEN_BITS[6].APB_32.edge_neg_93_iv_i_0_0[6]  
        (.A(\CoreGPIO_0/CONFIG_reg[6][3] ), .B(
        \CoreGPIO_0/edge_neg[6] ), .C(
        \CoreAPB3_0_APBmslave3_PWDATA[6] ), .D(\CoreGPIO_0/N_688 ), .Y(
        \CoreGPIO_0/N_113 ));
    sdf_IOPADP_TRI \FIC_MSS_0/MDDR_CLK_PAD/U_IOPADP  (.PAD_P(MDDR_CLK), 
        .OIN_P(\FIC_MSS_0/MSS_ADLIB_INST_DRAM_CLK ), .EIN_P(VCC));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_200_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_121_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_200_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_200_rs_net_1 ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_44  (.A(GND), 
        .B(VCC), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[27] ), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_READY_net ), .IPC());
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_82  (
        .A(\reg_apb_wrp_0/reg16x8_0/mem_0_[2]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_496 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_82_net_1 ));
    CFG4 #( .INIT(16'h5D55) )  
        \CoreAPB3_0/u_mux_p_to_b3/PRDATA_0_iv[7]  (.A(
        \CoreAPB3_0/u_mux_p_to_b3/PRDATA_0_iv_1[7]_net_1 ), .B(
        \CoreGPIO_0.CONFIG_reg_o_2[7] ), .C(
        \CoreAPB3_0_APBmslave3_PADDR[7] ), .D(
        CoreAPB3_0_APBmslave5_PSELx), .Y(
        \FIC_MSS_0_FIC_0_APB_MASTER_PRDATA[7] ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[6].gpin1[6]  (.D(\GPIO_IN_c[6] ), 
        .CLK(\FCCC_0/GL1_INST/U0_RGB1_RGB12_rgbr_net_1 ), .EN(VCC), 
        .ALn(\MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB2_rgbr_net_1 ), 
        .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/gpin1[6] ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_4_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB11_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_4__1_sqmuxa ), .ALn(
        AFLSDF_INV_11_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(GND)
        , .Q(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_4_set_net_1 ));
    CFG4 #( .INIT(16'hB383) )  \CoreGPIO_0/CONFIG_reg_o_2_31_bm[0]  (
        .A(\CoreGPIO_0/CONFIG_reg_o_2_31_bm_RNO[0]_net_1 ), .B(
        \CoreGPIO_0/CONFIG_reg_o_2_31_bm_1[0] ), .C(
        \CoreAPB3_0_APBmslave3_PADDR[3] ), .D(
        \CoreGPIO_0/CONFIG_reg_o_2_31_bm_RNO_0[0]_net_1 ), .Y(
        \CoreGPIO_0/CONFIG_reg_o_2_31_bm[0]_net_1 ));
    CFG4 #( .INIT(16'hF2F3) )  
        \CoreGPIO_0/xhdl1.GEN_BITS[23].APB_32.INTR_reg_308_0_o2_1_0[23]  
        (.A(\CoreGPIO_0/CONFIG_reg[23][6] ), .B(
        \CoreGPIO_0/edge_neg[23] ), .C(
        \CoreGPIO_0/INTR_reg_308_0_o2_0[23] ), .D(
        \CoreGPIO_0/CONFIG_reg[23][5] ), .Y(
        \CoreGPIO_0/INTR_reg_308_0_o2_1[23] ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[23].REG_GEN.CONFIG_reg[23][2]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[2] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB11_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[23]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB1_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[23][2] ));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_15_[6]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[6] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB7_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_15__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_255_i ), .ADn(VCC), .SLn(
        VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_15_rs[6] ));
    CFG4 #( .INIT(16'hC480) )  
        \CoreGPIO_0/xhdl1.GEN_BITS[6].APB_32.INTR_reg_87_0_0_RNO[6]  (
        .A(\CoreGPIO_0/CONFIG_reg[6][7] ), .B(
        \CoreGPIO_0/CONFIG_reg[6][3] ), .C(
        \CoreGPIO_0/INTR_reg_87_0_0_55_tz_1 ), .D(
        \CoreGPIO_0/INTR_reg_87_0_0_m2[6] ), .Y(\CoreGPIO_0/N_1580_tz )
        );
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[12].REG_GEN.CONFIG_reg[12][3]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[3] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB12_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[12]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB2_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[12][3] ));
    CFG4 #( .INIT(16'h0F35) )  
        \CoreGPIO_0/CONFIG_reg_o_2_31_am_RNO_2[0]  (.A(
        \CoreGPIO_0/CONFIG_reg[6][0] ), .B(
        \CoreGPIO_0/CONFIG_reg[22][0] ), .C(
        \CoreAPB3_0_APBmslave3_PADDR[6] ), .D(
        \CoreAPB3_0_APBmslave3_PADDR[5] ), .Y(
        \CoreGPIO_0/CONFIG_reg_o_2_13_1_1[0] ));
    CFG4 #( .INIT(16'h0F35) )  
        \CoreGPIO_0/CONFIG_reg_o_2_31_am_RNO_1[4]  (.A(
        \CoreGPIO_0/CONFIG_reg[2][4] ), .B(
        \CoreGPIO_0/CONFIG_reg[18][4] ), .C(
        \CoreAPB3_0_APBmslave3_PADDR[6] ), .D(
        \CoreAPB3_0_APBmslave3_PADDR[5] ), .Y(
        \CoreGPIO_0/CONFIG_reg_o_2_10_1_1[4] ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_51  (.A(GND), 
        .B(GND), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[5] ), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[12] ), .IPC());
    CFG4 #( .INIT(16'h7350) )  
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_3[1]  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_11_[1]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/mem_3_[1]_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/N_505 ), .D(
        \reg_apb_wrp_0/reg16x8_0/N_494 ), .Y(
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_3[1]_net_1 ));
    IOBI_IB_OB_EB \FIC_MSS_0/MDDR_DQ_14_PAD/U_IOBI  (.D(VCC), .E(VCC), 
        .YIN(\FIC_MSS_0/MDDR_DQ_14_PAD/YIN ), .DOUT(), .EOUT(), .Y());
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_92  (
        .A(\reg_apb_wrp_0/reg16x8_0/mem_11_[4]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_505 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_92_net_1 ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[0].REG_GEN.CONFIG_reg[0][2]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[2] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB15_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[0]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB5_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[0][2] ));
    CFG4 #( .INIT(16'h0200) )  
        \reg_apb_wrp_0/reg16x8_0/WRITE_GEN.mem_10__2_i_a2[7]  (.A(
        \CoreAPB3_0_APBmslave3_PADDR[3] ), .B(
        \CoreAPB3_0_APBmslave3_PADDR[2] ), .C(
        \CoreAPB3_0_APBmslave3_PADDR[0] ), .D(
        \CoreAPB3_0_APBmslave3_PADDR[1] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/N_491 ));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_84_set_RNIK14P  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_84_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_130_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_0_rs[3] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_0_[3]_net_1 ));
    CFG3 #( .INIT(8'h4C) )  \FIC_MSS_0/MSS_ADLIB_INST_RNO_16  (.A(
        \CoreGPIO_0.xhdl1.GEN_BITS[0].APB_32.GPOUT_reg9 ), .B(
        \FIC_MSS_0/CoreAPB3_0_APBmslave5_PRDATA_m_0_1_0[1] ), .C(
        \CoreGPIO_0.xhdl1.GEN_BITS[1].APB_32.GPOUT_reg[1] ), .Y(
        \FIC_MSS_0/CoreAPB3_0_APBmslave5_PRDATA_m_0_1_1[1] ));
    sdf_IOPADN_BI \FIC_MSS_0/MDDR_DQS_0_PAD/U_IOPADN  (.PAD_P(
        MDDR_DQS_N[0]), .OIN_P(\FIC_MSS_0/DRAM_DQS_OUT_net_0[0] ), 
        .EIN_P(\FIC_MSS_0/DRAM_DQS_OE_net_0[0] ), .N2POUT_P(
        \FIC_MSS_0/MDDR_DQS_0_PAD/U2_N2P ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_238  (.A(VCC), 
        .B(VCC), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[36] ), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[48] ), .IPC());
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_77  (
        .A(\reg_apb_wrp_0/reg16x8_0/mem_9_[5]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_492 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_77_net_1 ));
    CFG4 #( .INIT(16'h4657) )  
        \CoreGPIO_0/CONFIG_reg_o_2_31_am_1_1[6]  (.A(
        \CoreAPB3_0_APBmslave3_PADDR[4] ), .B(
        \CoreAPB3_0_APBmslave3_PADDR[3] ), .C(
        \CoreGPIO_0/CONFIG_reg_o_2_31_am_1_1_RNO[6]_net_1 ), .D(
        \CoreGPIO_0/CONFIG_reg_o_2_31_am_1_RNO_0[6]_net_1 ), .Y(
        \CoreGPIO_0/CONFIG_reg_o_2_31_am_1[6] ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[29].APB_32.edge_both[29]  (.D(
        \CoreGPIO_0/edge_neg_415[29] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB13_rgbr_net_1 ), .EN(
        \CoreGPIO_0/N_190 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB3_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/edge_pos[29] ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[8].APB_32.INTR_reg[8]  (.D(
        \CoreGPIO_0/INTR_reg_113[8] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB9_rgbr_net_1 ), .EN(VCC), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_YR ), .ADn(VCC), .SLn(
        VCC), .SD(GND), .LAT(GND), .Q(\CoreGPIO_0/INTR_reg[8] ));
    CFG4 #( .INIT(16'h0F35) )  
        \CoreGPIO_0/CONFIG_reg_o_2_31_bm_RNO_1[1]  (.A(
        \CoreGPIO_0.xhdl1.GEN_BITS[3].REG_GEN.CONFIG_reg[3][1] ), .B(
        \CoreGPIO_0/CONFIG_reg[19][1] ), .C(
        \CoreAPB3_0_APBmslave3_PADDR[6] ), .D(
        \CoreAPB3_0_APBmslave3_PADDR[5] ), .Y(
        \CoreGPIO_0/CONFIG_reg_o_2_25_1_1[1] ));
    CFG3 #( .INIT(8'hF2) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_174  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_5_[1]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_490 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_174_i ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[14].APB_32.edge_both[14]  (.D(
        \CoreGPIO_0/edge_neg_205[14] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB13_rgbr_net_1 ), .EN(
        \CoreGPIO_0/edge_pos_2_sqmuxa_8_i_1 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB3_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/edge_neg[14] ));
    CFG3 #( .INIT(8'hF2) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_203  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_10_[6]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_491 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_203_i ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_41  (.A(GND), 
        .B(GND), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[24] ), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[31] ), .IPC());
    CFG4 #( .INIT(16'hA9FF) )  
        \CoreGPIO_0/xhdl1.GEN_BITS[8].APB_32.INTR_reg_113_0_o2_0_0[8]  
        (.A(\CoreGPIO_0/CONFIG_reg[8][7] ), .B(
        \CoreGPIO_0/CONFIG_reg[8][6] ), .C(
        \CoreGPIO_0/CONFIG_reg[8][5] ), .D(
        \CoreGPIO_0/CONFIG_reg[8][3] ), .Y(
        \CoreGPIO_0/INTR_reg_113_0_o2_0[8] ));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/mem_15__RNIL8TK[1]  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_59_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_249_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_15_rs[1] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_15_[1]_net_1 ));
    CFG4 #( .INIT(16'hEAFA) )  \FIC_MSS_0/MSS_ADLIB_INST_RNO_0  (.A(
        \FIC_MSS_0/CoreAPB3_0_APBmslave5_PRDATA_m_0_0[1] ), .B(
        \CoreGPIO_0.PRDATA_iv_0_0_0_0[1] ), .C(
        CoreAPB3_0_APBmslave5_PSELx), .D(
        \FIC_MSS_0/CoreAPB3_0_APBmslave5_PRDATA_m_0_1_1[1] ), .Y(
        \FIC_MSS_0/FIC_MSS_0_FIC_0_APB_MASTER_PRDATA[1] ));
    CFG2 #( .INIT(4'h8) )  \FIC_MSS_0/MSS_ADLIB_INST_RNO_26  (.A(
        CoreAPB3_0_APBmslave5_PSELx), .B(
        \CoreGPIO_0.xhdl1.GEN_BITS[6].APB_32.INTR_reg[6] ), .Y(
        \FIC_MSS_0/CoreAPB3_0_APBmslave5_PRDATA_m_c_c_0[6] ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_87_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB16_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_0__1_sqmuxa ), .ALn(
        AFLSDF_INV_12_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(GND)
        , .Q(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_87_set_net_1 ));
    CFG4 #( .INIT(16'hCC0A) )  
        \CoreGPIO_0/xhdl1.GEN_BITS[4].APB_32.INTR_reg_61_0_0[4]  (.A(
        \CoreGPIO_0.xhdl1.GEN_BITS[4].APB_32.INTR_reg[4] ), .B(
        \CoreGPIO_0/N_1578_tz ), .C(\CoreAPB3_0_APBmslave3_PWDATA[4] ), 
        .D(\CoreGPIO_0/N_248 ), .Y(\CoreGPIO_0/INTR_reg_61[4] ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_230_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_22_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_230_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_230_rs_net_1 ));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/mem_3__RNITLDU[5]  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_52_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_157_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_3_rs[5] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_3_[5]_net_1 ));
    sdf_IOPAD_BI \FIC_MSS_0/MDDR_DQ_2_PAD/U_IOPAD  (.PAD(MDDR_DQ[2]), 
        .D(\FIC_MSS_0/DRAM_DQ_OUT_net_0[2] ), .E(
        \FIC_MSS_0/DRAM_DQ_OE_net_0[2] ), .Y(
        \FIC_MSS_0/MDDR_DQ_2_PAD_Y ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_108_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB5_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_13__1_sqmuxa ), .ALn(
        AFLSDF_INV_13_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(GND)
        , .Q(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_108_set_net_1 ));
    CFG4 #( .INIT(16'hC480) )  
        \CoreGPIO_0/xhdl1.GEN_BITS[2].APB_32.INTR_reg_35_0_0_RNO[2]  (
        .A(\CoreGPIO_0/CONFIG_reg[2][7] ), .B(
        \CoreGPIO_0/CONFIG_reg[2][3] ), .C(
        \CoreGPIO_0/INTR_reg_35_0_0_52_tz_1 ), .D(\CoreGPIO_0/N_178 ), 
        .Y(\CoreGPIO_0/N_1577_tz ));
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_69  (
        .A(\reg_apb_wrp_0/reg16x8_0/mem_8_[5]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_499 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_69_net_1 ));
    CFG4 #( .INIT(16'hF2F3) )  
        \CoreGPIO_0/xhdl1.GEN_BITS[29].APB_32.INTR_reg_386_0_o2_1_0[29]  
        (.A(\CoreGPIO_0/CONFIG_reg[29][6] ), .B(
        \CoreGPIO_0/edge_pos[29] ), .C(
        \CoreGPIO_0/INTR_reg_386_0_o2_0[29] ), .D(
        \CoreGPIO_0/CONFIG_reg[29][5] ), .Y(
        \CoreGPIO_0/INTR_reg_386_0_o2_1[29] ));
    IOIN_IB \GPIO_IN_ibuf[0]/U0/U_IOIN  (.YIN(\GPIO_IN_ibuf[0]/U0/YIN )
        , .E(GND), .Y(\GPIO_IN_c[0] ));
    CFG4 #( .INIT(16'h8000) )  
        \reg_apb_wrp_0/reg16x8_0/WRITE_GEN.mem_15__2_i_a2[7]  (.A(
        \CoreAPB3_0_APBmslave3_PADDR[3] ), .B(
        \CoreAPB3_0_APBmslave3_PADDR[2] ), .C(
        \CoreAPB3_0_APBmslave3_PADDR[0] ), .D(
        \CoreAPB3_0_APBmslave3_PADDR[1] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/N_497 ));
    IOINFF_BYPASS \GPIO_IN_ibuf[5]/U0/U_IOINFF  (.A(
        \GPIO_IN_ibuf[5]/U0/YIN1 ), .Y(\GPIO_IN_ibuf[5]/U0/YIN ));
    CFG3 #( .INIT(8'hF2) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_168  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_4_[6]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_504 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_168_i ));
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_29  (
        .A(\reg_apb_wrp_0/reg16x8_0/mem_6_[0]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_493 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_29_net_1 ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[27].REG_GEN.CONFIG_reg[27][7]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[7] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB9_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[27]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_YR ), .ADn(VCC), .SLn(
        VCC), .SD(GND), .LAT(GND), .Q(\CoreGPIO_0/CONFIG_reg[27][7] ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[1].REG_GEN.CONFIG_reg[1][3]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[3] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB15_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[1]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB5_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[1][3] ));
    CFG4 #( .INIT(16'hEC00) )  \CoreAPB3_0/u_mux_p_to_b3/PRDATA[31]  (
        .A(\CoreGPIO_0.xhdl1.GEN_BITS[0].APB_32.GPOUT_reg9 ), .B(
        \CoreGPIO_0.N_524 ), .C(
        \CoreGPIO_0.xhdl1.GEN_BITS[31].APB_32.GPOUT_reg[31] ), .D(
        CoreAPB3_0_APBmslave5_PSELx), .Y(
        \FIC_MSS_0_FIC_0_APB_MASTER_PRDATA[31] ));
    CFG4 #( .INIT(16'h0F35) )  
        \CoreGPIO_0/CONFIG_reg_o_2_31_bm_RNO_1[6]  (.A(
        \CoreGPIO_0/CONFIG_reg[3][6] ), .B(
        \CoreGPIO_0/CONFIG_reg[19][6] ), .C(
        \CoreAPB3_0_APBmslave3_PADDR[6] ), .D(
        \CoreAPB3_0_APBmslave3_PADDR[5] ), .Y(
        \CoreGPIO_0/CONFIG_reg_o_2_25_1_1[6] ));
    IOINFF_BYPASS \FIC_MSS_0/MDDR_DQ_10_PAD/U_IOINFF  (.A(
        \FIC_MSS_0/MDDR_DQ_10_PAD_Y ), .Y(
        \FIC_MSS_0/MDDR_DQ_10_PAD/YIN ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[26].REG_GEN.CONFIG_reg[26][0]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[0] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB16_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[26]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB6_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[26][0] ));
    CFG4 #( .INIT(16'h7350) )  
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_0[4]  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_13_[4]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/mem_5_[4]_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/N_500 ), .D(
        \reg_apb_wrp_0/reg16x8_0/N_490 ), .Y(
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_0[4]_net_1 ));
    IOENFF_BYPASS \GPIO_OUT_obuf[2]/U0/U_IOENFF  (.A(
        \GPIO_OUT_obuf[2]/U0/EOUT1 ), .Y(\GPIO_OUT_obuf[2]/U0/EOUT ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_38  (.A(GND), 
        .B(VCC), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[21] ), .IPB(), .IPC());
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_149  (.A(VCC), 
        .B(VCC), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/I2C1_SCL_F2H_SCP_net ), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/MGPIO5A_F2H_GPIN_net ), .IPC());
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_145  (.A(GND), 
        .B(VCC), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/SLEEPHOLDREQ_net ), .IPB(), .IPC());
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[7].REG_GEN.CONFIG_reg[7][1]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[1] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB11_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[7]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB1_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[7][1] ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_106  (.A(VCC), 
        .B(VCC), .C(VCC), .IPA(), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/FAB_TXREADY_net ), .IPC());
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_65  (.A(GND), 
        .B(VCC), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[26] ), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PSLVERR_net ), .IPC());
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[23].REG_GEN.CONFIG_reg[23][6]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[6] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB10_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[23]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB0_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[23][6] ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_183_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_76_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_183_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_183_rs_net_1 ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[22].APB_32.INTR_reg[22]  (.D(
        \CoreGPIO_0/INTR_reg_295[22] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB13_rgbr_net_1 ), .EN(VCC), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB3_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/INTR_reg[22] ));
    CFG4 #( .INIT(16'hA9FF) )  
        \CoreGPIO_0/xhdl1.GEN_BITS[13].APB_32.INTR_reg_178_0_o2_0_0[13]  
        (.A(\CoreGPIO_0/CONFIG_reg[13][7] ), .B(
        \CoreGPIO_0/CONFIG_reg[13][6] ), .C(
        \CoreGPIO_0/CONFIG_reg[13][5] ), .D(
        \CoreGPIO_0/CONFIG_reg[13][3] ), .Y(
        \CoreGPIO_0/INTR_reg_178_0_o2_0[13] ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_70  (.A(VCC), 
        .B(VCC), .C(VCC), .IPA(), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[4] ), .IPC());
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_160  (.A(VCC), 
        .B(VCC), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/MGPIO11A_F2H_GPIN_net ), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/MGPIO14A_F2H_GPIN_net ), .IPC());
    IOTRI_OB_EB \GPIO_OUT_obuf[5]/U0/U_IOTRI  (.D(\GPIO_OUT_net_2[5] ), 
        .E(VCC), .DOUT(\GPIO_OUT_obuf[5]/U0/DOUT1 ), .EOUT(
        \GPIO_OUT_obuf[5]/U0/EOUT1 ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_266  (.A(VCC), 
        .B(GND), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[26] ), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/F_ARLOCK_HMASTLOCK1_net[0] ), .IPC());
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/mem_2__RNIRDSQ[4]  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_34_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_148_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_2_rs[4] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_2_[4]_net_1 ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_23  (.A(VCC), 
        .B(GND), .C(VCC), .IPA(), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_TRANS1_net ), .IPC());
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_14_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB15_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_1__1_sqmuxa ), .ALn(
        AFLSDF_INV_14_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(GND)
        , .Q(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_14_set_net_1 ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[7].APB_32.GPOUT_reg[7]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[7] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB11_rgbr_net_1 ), .EN(
        \CoreGPIO_0/GPOUT_reg_0_sqmuxa ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB1_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/GPOUT_reg[7] ));
    IOTRI_OB_EB \FIC_MSS_0/MDDR_ADDR_5_PAD/U_IOOUT  (.D(VCC), .E(VCC), 
        .DOUT(), .EOUT(\FIC_MSS_0/MDDR_ADDR_5_PAD/EOUT ));
    INV_BA AFLSDF_INV_107 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_30_net_1 ), .Y(
        AFLSDF_INV_107_net_1));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[8].REG_GEN.CONFIG_reg[8][6]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[6] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB9_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[8]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_YR ), .ADn(VCC), .SLn(
        VCC), .SD(GND), .LAT(GND), .Q(\CoreGPIO_0/CONFIG_reg[8][6] ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[25].REG_GEN.CONFIG_reg[25][5]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[5] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB15_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[25]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB5_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[25][5] ));
    CFG4 #( .INIT(16'hA9FF) )  
        \CoreGPIO_0/xhdl1.GEN_BITS[22].APB_32.INTR_reg_295_0_o2_0_0[22]  
        (.A(\CoreGPIO_0/CONFIG_reg[22][7] ), .B(
        \CoreGPIO_0/CONFIG_reg[22][6] ), .C(
        \CoreGPIO_0/CONFIG_reg[22][5] ), .D(
        \CoreGPIO_0/CONFIG_reg[22][3] ), .Y(
        \CoreGPIO_0/INTR_reg_295_0_o2_0[22] ));
    CFG4 #( .INIT(16'hF2F3) )  
        \CoreGPIO_0/xhdl1.GEN_BITS[18].APB_32.INTR_reg_243_0_o2_1_0[18]  
        (.A(\CoreGPIO_0/CONFIG_reg[18][6] ), .B(
        \CoreGPIO_0/edge_neg[18] ), .C(
        \CoreGPIO_0/INTR_reg_243_0_o2_0[18] ), .D(
        \CoreGPIO_0/CONFIG_reg[18][5] ), .Y(
        \CoreGPIO_0/INTR_reg_243_0_o2_1[18] ));
    INV_BA AFLSDF_INV_65 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_116_net_1 ), .Y(
        AFLSDF_INV_65_net_1));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_38_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB13_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_2__1_sqmuxa ), .ALn(
        AFLSDF_INV_15_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(GND)
        , .Q(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_38_set_net_1 ));
    INV_BA AFLSDF_INV_43 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_126_net_1 ), .Y(
        AFLSDF_INV_43_net_1));
    CFG4 #( .INIT(16'h0F35) )  
        \CoreGPIO_0/CONFIG_reg_o_2_31_bm_1_RNO_2[7]  (.A(
        \CoreGPIO_0/CONFIG_reg[1][7] ), .B(
        \CoreGPIO_0/CONFIG_reg[17][7] ), .C(
        \CoreAPB3_0_APBmslave3_PADDR[6] ), .D(
        \CoreAPB3_0_APBmslave3_PADDR[5] ), .Y(
        \CoreGPIO_0/CONFIG_reg_o_2_18_1[7] ));
    CFG4 #( .INIT(16'h4657) )  
        \CoreGPIO_0/CONFIG_reg_o_2_31_am_1_1[4]  (.A(
        \CoreAPB3_0_APBmslave3_PADDR[4] ), .B(
        \CoreAPB3_0_APBmslave3_PADDR[3] ), .C(
        \CoreGPIO_0/CONFIG_reg_o_2_31_am_1_1_RNO[4]_net_1 ), .D(
        \CoreGPIO_0/CONFIG_reg_o_2_31_am_1_RNO_0[4]_net_1 ), .Y(
        \CoreGPIO_0/CONFIG_reg_o_2_31_am_1[4] ));
    IOTRI_OB_EB \FIC_MSS_0/MDDR_ADDR_0_PAD/U_IOOUT  (.D(VCC), .E(VCC), 
        .DOUT(), .EOUT(\FIC_MSS_0/MDDR_ADDR_0_PAD/EOUT ));
    INV_BA AFLSDF_INV_21 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_122_net_1 ), .Y(
        AFLSDF_INV_21_net_1));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_155_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_48_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_155_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_155_rs_net_1 ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_232  (.A(VCC), 
        .B(VCC), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[30] ), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[42] ), .IPC());
    INV_BA AFLSDF_INV_81 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_50_net_1 ), .Y(
        AFLSDF_INV_81_net_1));
    CFG4 #( .INIT(16'hAC0F) )  
        \CoreGPIO_0/CONFIG_reg_o_2_31_am_1_1_RNO[4]  (.A(
        \CoreGPIO_0/CONFIG_reg[12][4] ), .B(
        \CoreGPIO_0/CONFIG_reg[28][4] ), .C(
        \CoreGPIO_0/CONFIG_reg_o_2_6_1[4] ), .D(
        \CoreAPB3_0_APBmslave3_PADDR[5] ), .Y(
        \CoreGPIO_0/CONFIG_reg_o_2_31_am_1_1_RNO[4]_net_1 ));
    CFG4 #( .INIT(16'hB383) )  \CoreGPIO_0/CONFIG_reg_o_2_31_am[1]  (
        .A(\CoreGPIO_0/CONFIG_reg_o_2_31_am_RNO[1]_net_1 ), .B(
        \CoreGPIO_0/CONFIG_reg_o_2_31_am_1[1] ), .C(
        \CoreAPB3_0_APBmslave3_PADDR[3] ), .D(
        \CoreGPIO_0/CONFIG_reg_o_2_31_am_RNO_0[1]_net_1 ), .Y(
        \CoreGPIO_0/CONFIG_reg_o_2_31_am[1]_net_1 ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_14  (.A(
        \FIC_MSS_0_FIC_0_APB_MASTER_PRDATA[19] ), .B(VCC), .C(VCC), 
        .IPA(\FIC_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[19] ), .IPB(), 
        .IPC());
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_201  (.A(VCC), 
        .B(VCC), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[5] ), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[17] ), .IPC());
    CFG4 #( .INIT(16'hEFEE) )  
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_11[2]  (.A(
        \reg_apb_wrp_0/reg16x8_0/N_400 ), .B(
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_7[2]_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_0_[2]_net_1 ), .D(
        \reg_apb_wrp_0/reg16x8_0/N_496 ), .Y(
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_11[2]_net_1 ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_97  (.A(VCC), 
        .B(VCC), .C(VCC), .IPA(\FIC_MSS_0/MSS_ADLIB_INST/COLF_net ), 
        .IPB(), .IPC());
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_119  (.A(VCC), 
        .B(VCC), .C(VCC), .IPA(), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/FAB_RXERROR_net ), .IPC());
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_115  (.A(VCC), 
        .B(VCC), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/FAB_XDATAIN_net[7] ), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/FAB_VSTATUS_net[4] ), .IPC());
    CFG4 #( .INIT(16'h0F35) )  
        \CoreGPIO_0/CONFIG_reg_o_2_31_bm_RNO_2[4]  (.A(
        \CoreGPIO_0/CONFIG_reg[7][4] ), .B(
        \CoreGPIO_0/CONFIG_reg[23][4] ), .C(
        \CoreAPB3_0_APBmslave3_PADDR[6] ), .D(
        \CoreAPB3_0_APBmslave3_PADDR[5] ), .Y(
        \CoreGPIO_0/CONFIG_reg_o_2_28_1_1[4] ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[24].REG_GEN.CONFIG_reg[24][6]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[6] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB11_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[24]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB1_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[24][6] ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_103  (.A(VCC), 
        .B(VCC), .C(VCC), .IPA(\FIC_MSS_0/MSS_ADLIB_INST/RCGF_net[3] ), 
        .IPB(\FIC_MSS_0/MSS_ADLIB_INST/XCLK_FAB_net ), .IPC());
    INV_BA AFLSDF_INV_46 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_101_net_1 ), .Y(
        AFLSDF_INV_46_net_1));
    CFG3 #( .INIT(8'h32) )  \reg_apb_wrp_0/fsm_ns_1_0_.m2  (.A(
        \reg_apb_wrp_0/fsm[1]_net_1 ), .B(\reg_apb_wrp_0/fsm[0]_net_1 )
        , .C(CoreAPB3_0_APBmslave3_PSELx), .Y(
        \reg_apb_wrp_0/fsm_ns[0] ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_247_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_119_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_247_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_247_rs_net_1 ));
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_118  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_14_[6]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_503 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_118_net_1 ));
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_65  (
        .A(\reg_apb_wrp_0/reg16x8_0/mem_4_[4]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_504 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_65_net_1 ));
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_4_[0]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_504 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_net_1 ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_137  (.A(VCC), 
        .B(VCC), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/I2C1_BCLK_net ), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/F_DMAREADY_net[1] ), .IPC());
    CFG4 #( .INIT(16'hAA08) )  
        \CoreGPIO_0/xhdl1.GEN_BITS[1].APB_32.edge_neg_23_iv_i_0[1]  (
        .A(\CoreGPIO_0/CONFIG_reg[1][3] ), .B(\CoreGPIO_0/edge_neg[1] )
        , .C(\CoreAPB3_0_APBmslave3_PWDATA[1] ), .D(\CoreGPIO_0/N_399 )
        , .Y(\CoreGPIO_0/N_121 ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_181  (.A(VCC), 
        .B(VCC), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/MMUART0_DCD_F2H_SCP_net ), .IPB(), 
        .IPC());
    CFG3 #( .INIT(8'h20) )  
        \CoreGPIO_0/xhdl1.GEN_BITS[22].APB_32.edge_both_RNO[22]  (.A(
        \CoreGPIO_0/CONFIG_reg[22][3] ), .B(
        \CoreAPB3_0_APBmslave3_PWDATA[22] ), .C(
        \CoreGPIO_0/edge_neg[22] ), .Y(\CoreGPIO_0/edge_neg_317[22] ));
    CFG4 #( .INIT(16'h7350) )  
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_3[3]  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_11_[3]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/mem_3_[3]_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/N_505 ), .D(
        \reg_apb_wrp_0/reg16x8_0/N_494 ), .Y(
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_3[3]_net_1 ));
    IOINFF_BYPASS \FIC_MSS_0/MDDR_DQ_7_PAD/U_IOINFF  (.A(
        \FIC_MSS_0/MDDR_DQ_7_PAD_Y ), .Y(\FIC_MSS_0/MDDR_DQ_7_PAD/YIN )
        );
    CFG3 #( .INIT(8'hF2) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_163  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_4_[2]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_504 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_163_i ));
    GB MSS_RESET_N_F2M_ibuf_RNIBBDD (.An(AFLSDF_INV_16_net_1), .ENn(
        GND), .YNn(), .YSn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_YNn_GSouth ));
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_25  (
        .A(\reg_apb_wrp_0/reg16x8_0/mem_5_[6]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_490 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_25_net_1 ));
    CFG2 #( .INIT(4'h8) )  
        \CoreGPIO_0/xhdl1.GEN_BITS[5].REG_GPOUT.un54_GPIO_OUT_i  (.A(
        \CoreGPIO_0.xhdl1.GEN_BITS[5].APB_32.GPOUT_reg[5] ), .B(
        \CoreGPIO_0/CONFIG_reg[5][0] ), .Y(\GPIO_OUT_net_2[5] ));
    CFG4 #( .INIT(16'h7530) )  
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_1[3]  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_15_[3]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/mem_7_[3]_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/N_498 ), .D(
        \reg_apb_wrp_0/reg16x8_0/N_497 ), .Y(
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_1[3]_net_1 ));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/mem_3__RNI5HO01[1]  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_124_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_153_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_3_rs[1] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_3_[1]_net_1 ));
    sdf_IOPAD_IN \GPIO_IN_ibuf[2]/U0/U_IOPAD  (.PAD(GPIO_IN[2]), .Y(
        \GPIO_IN_ibuf[2]/U0/YIN1 ));
    CFG4 #( .INIT(16'h5410) )  \CoreGPIO_0/PRDATA_iv_0_0_1[4]  (.A(
        \CoreAPB3_0_APBmslave3_PADDR[7] ), .B(
        \CoreAPB3_0_APBmslave3_PADDR[2] ), .C(
        \CoreGPIO_0/CONFIG_reg_o_2_31_am[4]_net_1 ), .D(
        \CoreGPIO_0/CONFIG_reg_o_2_31_bm[4]_net_1 ), .Y(
        \CoreGPIO_0.PRDATA_iv_0_0_1[4] ));
    CFG2 #( .INIT(4'h4) )  \CoreGPIO_0/PRDATA_0_iv_0_a2_0[23]  (.A(
        \CoreGPIO_0.N_247 ), .B(\CoreGPIO_0/INTR_reg[23] ), .Y(
        \CoreGPIO_0.N_540 ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[21].REG_GEN.CONFIG_reg[21][4]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[4] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB14_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[21]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB4_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[21][4] ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_11  (.A(VCC), 
        .B(\FIC_MSS_0_FIC_0_APB_MASTER_PRDATA[16] ), .C(VCC), .IPA(), 
        .IPB(\FIC_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[16] ), .IPC());
    SLE \reg_apb_wrp_0/fsm[0]  (.D(\reg_apb_wrp_0/fsm_ns[0] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB12_rgbr_net_1 ), .EN(VCC), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB2_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/fsm[0]_net_1 ));
    CFG4 #( .INIT(16'hB383) )  \CoreGPIO_0/CONFIG_reg_o_2_31_bm[4]  (
        .A(\CoreGPIO_0/CONFIG_reg_o_2_31_bm_RNO[4]_net_1 ), .B(
        \CoreGPIO_0/CONFIG_reg_o_2_31_bm_1[4] ), .C(
        \CoreAPB3_0_APBmslave3_PADDR[3] ), .D(
        \CoreGPIO_0/CONFIG_reg_o_2_31_bm_RNO_0[4]_net_1 ), .Y(
        \CoreGPIO_0/CONFIG_reg_o_2_31_bm[4]_net_1 ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[0].gpin2[0]  (.D(
        \CoreGPIO_0/gpin1[0] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB9_rgbr_net_1 ), .EN(VCC), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_YR ), .ADn(VCC), .SLn(
        VCC), .SD(GND), .LAT(GND), .Q(\CoreGPIO_0/gpin2[0] ));
    CFG4 #( .INIT(16'hAA08) )  
        \CoreGPIO_0/xhdl1.GEN_BITS[0].APB_32.edge_both_9_iv_i_0[0]  (
        .A(\CoreGPIO_0/CONFIG_reg[0][3] ), .B(
        \CoreGPIO_0/edge_both[0] ), .C(
        \CoreAPB3_0_APBmslave3_PWDATA[0] ), .D(\CoreGPIO_0/N_141_i ), 
        .Y(\CoreGPIO_0/N_97 ));
    CFG4 #( .INIT(16'hAC0F) )  
        \CoreGPIO_0/CONFIG_reg_o_2_31_am_RNO_0[3]  (.A(
        \CoreGPIO_0/CONFIG_reg[14][3] ), .B(
        \CoreGPIO_0/CONFIG_reg[30][3] ), .C(
        \CoreGPIO_0/CONFIG_reg_o_2_13_1_1[3] ), .D(
        \CoreAPB3_0_APBmslave3_PADDR[5] ), .Y(
        \CoreGPIO_0/CONFIG_reg_o_2_31_am_RNO_0[3]_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_227_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_19_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_227_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_227_rs_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_11_[2]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[2] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB17_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_11__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_211_i ), .ADn(VCC), .SLn(
        VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_11_rs[2] ));
    INV_BA AFLSDF_INV_39 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_73_net_1 ), .Y(
        AFLSDF_INV_39_net_1));
    CFG3 #( .INIT(8'hF2) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_161  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_4_[0]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_504 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_161_i ));
    IOBI_IB_OB_EB \FIC_MSS_0/MDDR_DQ_4_PAD/U_IOBI  (.D(VCC), .E(VCC), 
        .YIN(\FIC_MSS_0/MDDR_DQ_4_PAD/YIN ), .DOUT(), .EOUT(), .Y());
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_71_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB10_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_8__1_sqmuxa ), .ALn(
        AFLSDF_INV_17_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(GND)
        , .Q(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_71_set_net_1 ));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_134_rs_RNIUS2Q  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_87_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_134_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_0_rs[6] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_0_[6]_net_1 ));
    INV_BA AFLSDF_INV_37 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_1_net_1 ), .Y(
        AFLSDF_INV_37_net_1));
    CFG2 #( .INIT(4'h8) )  
        \reg_apb_wrp_0/reg16x8_0/mem_5__1_sqmuxa_0_a2_0_a3  (.A(
        \reg_apb_wrp_0/reg16x8_0/N_490 ), .B(
        \reg_apb_wrp_0/wr_enable_net_1 ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_5__1_sqmuxa ));
    CFG3 #( .INIT(8'hF2) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_210  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_7_[3]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_498 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_210_i ));
    CFG4 #( .INIT(16'h4657) )  
        \CoreGPIO_0/CONFIG_reg_o_2_31_bm_1_1[6]  (.A(
        \CoreAPB3_0_APBmslave3_PADDR[4] ), .B(
        \CoreAPB3_0_APBmslave3_PADDR[3] ), .C(
        \CoreGPIO_0/CONFIG_reg_o_2_31_bm_1_1_RNO[6]_net_1 ), .D(
        \CoreGPIO_0/CONFIG_reg_o_2_31_bm_1_RNO_0[6]_net_1 ), .Y(
        \CoreGPIO_0/CONFIG_reg_o_2_31_bm_1[6] ));
    IOTRI_OB_EB \GPIO_OUT_obuf[6]/U0/U_IOTRI  (.D(\GPIO_OUT_net_2[6] ), 
        .E(VCC), .DOUT(\GPIO_OUT_obuf[6]/U0/DOUT1 ), .EOUT(
        \GPIO_OUT_obuf[6]/U0/EOUT1 ));
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_67  (
        .A(\reg_apb_wrp_0/reg16x8_0/mem_4_[5]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_504 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_67_net_1 ));
    CFG3 #( .INIT(8'h40) )  \CoreGPIO_0/PRDATA_0_iv_0_a2[26]  (.A(
        \CoreGPIO_0.N_246 ), .B(\CoreGPIO_0/GPOUT_reg[26] ), .C(
        \CoreAPB3_0_APBmslave3_PADDR[5] ), .Y(\CoreGPIO_0.N_533 ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_264  (.A(VCC), 
        .B(GND), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[24] ), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/F_ARBURST_HTRANS1_net[0] ), .IPC(
        \FIC_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PENABLE_net ));
    sdf_IOPAD_TRI \FIC_MSS_0/MDDR_ADDR_2_PAD/U_IOPAD  (.PAD(
        MDDR_ADDR[2]), .D(\FIC_MSS_0/DRAM_ADDR_net_0[2] ), .E(
        \FIC_MSS_0/MDDR_ADDR_2_PAD/EOUT ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[1].REG_GEN.CONFIG_reg[1][6]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[6] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB15_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[1]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB5_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[1][6] ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[23].REG_GEN.CONFIG_reg[23][1]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[1] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB11_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[23]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB1_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[23][1] ));
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_36  (
        .A(\reg_apb_wrp_0/reg16x8_0/mem_2_[5]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_501 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_36_net_1 ));
    CFG3 #( .INIT(8'hF2) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_212  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_11_[3]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_505 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_212_i ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[13].APB_32.GPOUT_reg[13]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[13] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB11_rgbr_net_1 ), .EN(
        \CoreGPIO_0/GPOUT_reg_0_sqmuxa ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB1_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0.xhdl1.GEN_BITS[13].APB_32.GPOUT_reg[13] ));
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_27  (
        .A(\reg_apb_wrp_0/reg16x8_0/mem_5_[7]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_490 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_27_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_8_[4]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[4] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB18_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_8__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_167_i ), .ADn(VCC), .SLn(
        VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_8_rs[4] ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_80_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB2_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_0__1_sqmuxa ), .ALn(
        AFLSDF_INV_18_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(GND)
        , .Q(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_80_set_net_1 ));
    CFG2 #( .INIT(4'hE) )  
        \CoreGPIO_0/xhdl1.GEN_BITS[0].APB_32.un5_PRDATA_o_0_a2_0_o2_x  
        (.A(\CoreGPIO_0/un5_PRDATA_o_0_a2_0_o2_sx ), .B(
        \CoreAPB3_0_APBmslave3_PADDR[6] ), .Y(
        \xhdl1.GEN_BITS[0].APB_32.un5_PRDATA_o_0_a2_0_o2_x ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[20].REG_GEN.CONFIG_reg[20][1]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[1] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB12_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[20]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB2_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[20][1] ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[31].APB_32.INTR_reg[31]  (.D(
        \CoreGPIO_0/INTR_reg_412[31] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB9_rgbr_net_1 ), .EN(VCC), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_YR ), .ADn(VCC), .SLn(
        VCC), .SD(GND), .LAT(GND), .Q(\CoreGPIO_0/INTR_reg[31] ));
    CFG4 #( .INIT(16'hEC00) )  \CoreAPB3_0/u_mux_p_to_b3/PRDATA[30]  (
        .A(\CoreGPIO_0.xhdl1.GEN_BITS[0].APB_32.GPOUT_reg9 ), .B(
        \CoreGPIO_0.N_526 ), .C(
        \CoreGPIO_0.xhdl1.GEN_BITS[30].APB_32.GPOUT_reg[30] ), .D(
        CoreAPB3_0_APBmslave5_PSELx), .Y(
        \FIC_MSS_0_FIC_0_APB_MASTER_PRDATA[30] ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_143_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_24_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_143_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_143_rs_net_1 ));
    CFG3 #( .INIT(8'h20) )  
        \CoreGPIO_0/xhdl1.GEN_BITS[8].APB_32.edge_both_RNO[8]  (.A(
        \CoreGPIO_0/CONFIG_reg[8][3] ), .B(
        \CoreAPB3_0_APBmslave3_PWDATA[8] ), .C(
        \CoreGPIO_0/edge_pos[8] ), .Y(\CoreGPIO_0/edge_neg_121[8] ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_41_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB15_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_1__1_sqmuxa ), .ALn(
        AFLSDF_INV_19_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(GND)
        , .Q(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_41_set_net_1 ));
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_113  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_14_[1]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_503 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_113_net_1 ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_208  (.A(VCC), 
        .B(GND), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[26] ), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/F_AWBURST_HTRANS0_net[0] ), .IPC());
    RGB \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB1  (.An(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_YNn_GSouth ), .ENn(GND), .YL(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB1_rgbl_net_1 ), .YR(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB1_rgbr_net_1 ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[12].APB_32.GPOUT_reg[12]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[12] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB13_rgbr_net_1 ), .EN(
        \CoreGPIO_0/GPOUT_reg_0_sqmuxa ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB3_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0.xhdl1.GEN_BITS[12].APB_32.GPOUT_reg[12] ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_229  (.A(VCC), 
        .B(VCC), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[27] ), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[39] ), .IPC(
        \FIC_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[51] ));
    INV_BA AFLSDF_INV_111 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_62_net_1 ), .Y(
        AFLSDF_INV_111_net_1));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[3].REG_GEN.CONFIG_reg[3][3]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[3] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB9_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[3]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_YR ), .ADn(VCC), .SLn(
        VCC), .SD(GND), .LAT(GND), .Q(\CoreGPIO_0/CONFIG_reg[3][3] ));
    CFG3 #( .INIT(8'h20) )  
        \CoreGPIO_0/xhdl1.GEN_BITS[13].APB_32.edge_both_RNO[13]  (.A(
        \CoreGPIO_0/CONFIG_reg[13][3] ), .B(
        \CoreAPB3_0_APBmslave3_PWDATA[13] ), .C(
        \CoreGPIO_0/edge_neg[13] ), .Y(\CoreGPIO_0/edge_neg_191[13] ));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/mem_2__RNIVPBK[5]  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_36_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_149_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_2_rs[5] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_2_[5]_net_1 ));
    CFG4 #( .INIT(16'hEAFA) )  \FIC_MSS_0/MSS_ADLIB_INST_RNO_1  (.A(
        \FIC_MSS_0/CoreAPB3_0_APBmslave5_PRDATA_m_0_0[2] ), .B(
        \CoreGPIO_0.PRDATA_iv_0_0_0_0[2] ), .C(
        CoreAPB3_0_APBmslave5_PSELx), .D(
        \FIC_MSS_0/CoreAPB3_0_APBmslave5_PRDATA_m_0_1[2] ), .Y(
        \FIC_MSS_0/FIC_MSS_0_FIC_0_APB_MASTER_PRDATA[2] ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_55  (.A(GND), 
        .B(GND), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[9] ), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[16] ), .IPC());
    SLE \reg_apb_wrp_0/reg16x8_0/mem_3_[1]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[1] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB15_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_3__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_153_i ), .ADn(VCC), .SLn(
        VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_3_rs[1] ));
    sdf_IOPAD_BI \FIC_MSS_0/MDDR_DQ_14_PAD/U_IOPAD  (.PAD(MDDR_DQ[14]), 
        .D(\FIC_MSS_0/DRAM_DQ_OUT_net_0[14] ), .E(
        \FIC_MSS_0/DRAM_DQ_OE_net_0[14] ), .Y(
        \FIC_MSS_0/MDDR_DQ_14_PAD_Y ));
    CFG4 #( .INIT(16'h8000) )  
        \CoreGPIO_0/xhdl1.GEN_BITS[15].REG_GEN.CONFIG_reg[15]2_0_a4_0_a2  
        (.A(\CoreAPB3_0_APBmslave3_PADDR[3] ), .B(
        \CoreAPB3_0_APBmslave3_PADDR[2] ), .C(\CoreGPIO_0/N_604 ), .D(
        \CoreGPIO_0/N_605 ), .Y(\CoreGPIO_0/CONFIG_reg[15]2 ));
    CFG3 #( .INIT(8'hF2) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_208  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_7_[2]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_498 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_208_i ));
    IP_INTERFACE ip_interface_inst (.A(VCC), .B(ff_to_start_net), .C(
        VCC), .IPA(), .IPB(), .IPC());
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_203_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_103_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_203_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_203_rs_net_1 ));
    CFG4 #( .INIT(16'hB383) )  \CoreGPIO_0/CONFIG_reg_o_2_31_am[6]  (
        .A(\CoreGPIO_0/CONFIG_reg_o_2_31_am_RNO[6]_net_1 ), .B(
        \CoreGPIO_0/CONFIG_reg_o_2_31_am_1[6] ), .C(
        \CoreAPB3_0_APBmslave3_PADDR[3] ), .D(
        \CoreGPIO_0/CONFIG_reg_o_2_31_am_RNO_0[6]_net_1 ), .Y(
        \CoreGPIO_0/CONFIG_reg_o_2_31_am[6]_net_1 ));
    CFG4 #( .INIT(16'h0020) )  
        \reg_apb_wrp_0/reg16x8_0/WRITE_GEN.mem_9__2_i_a2[7]  (.A(
        \CoreAPB3_0_APBmslave3_PADDR[3] ), .B(
        \CoreAPB3_0_APBmslave3_PADDR[2] ), .C(
        \CoreAPB3_0_APBmslave3_PADDR[0] ), .D(
        \CoreAPB3_0_APBmslave3_PADDR[1] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/N_492 ));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_4_[5]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[5] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB16_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_4__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_166_i ), .ADn(VCC), .SLn(
        VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_4_rs[5] ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[15].REG_GEN.CONFIG_reg[15][2]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[2] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB11_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[15]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB1_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[15][2] ));
    CFG4 #( .INIT(16'h0001) )  
        \reg_apb_wrp_0/reg16x8_0/temp_data_RNO[5]  (.A(
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_0_0[5]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_0_1[5]_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_0_13[5]_net_1 ), .D(
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_0_9[5]_net_1 ), .Y(
        \reg_apb_wrp_0/reg16x8_0/N_25_i_0 ));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_164_rs_RNI9DOL  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_6_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_164_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_4_rs[3] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_4_[3]_net_1 ));
    INV_BA AFLSDF_INV_61 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_97_net_1 ), .Y(
        AFLSDF_INV_61_net_1));
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_111  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_13_[7]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_500 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_111_net_1 ));
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_78  (
        .A(\reg_apb_wrp_0/reg16x8_0/mem_9_[6]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_492 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_78_net_1 ));
    CFG3 #( .INIT(8'hF2) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_198  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_6_[5]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_493 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_198_i ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_83_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB17_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_3__1_sqmuxa ), .ALn(
        AFLSDF_INV_20_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(GND)
        , .Q(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_83_set_net_1 ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_45  (.A(GND), 
        .B(GND), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[28] ), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_ENABLE_net ), .IPC());
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_177_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_73_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_177_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_177_rs_net_1 ));
    CFG4 #( .INIT(16'hFFEA) )  \FIC_MSS_0/MSS_ADLIB_INST_RNO_2  (.A(
        \FIC_MSS_0/CoreAPB3_0_APBmslave5_PRDATA_m_0_0[3] ), .B(
        \FIC_MSS_0/CoreAPB3_0_APBmslave5_PRDATA_m_0_1[3] ), .C(
        CoreAPB3_0_APBmslave5_PSELx), .D(
        \FIC_MSS_0/CoreAPB3_0_APBmslave5_PRDATA_m_d[3] ), .Y(
        \FIC_MSS_0/FIC_MSS_0_FIC_0_APB_MASTER_PRDATA[3] ));
    CFG3 #( .INIT(8'hF2) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_184  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_5_[6]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_490 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_184_i ));
    MSS_010_IP #( .INIT(1438'h00000000003612000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000F00000000F000000000000000000000000000000007FFFFFFFB000001007C33C00020200609280104003FFFFE400000000000050000000000001C0000007EDFDC010842108421000001FE34001FF8000000400000000020091007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF)
        , .ACT_UBITS(56'hFFFFFFFFFFFFFF), .MEMORYFILE("ENVM_init.mem")
        , .RTC_MAIN_XTL_FREQ(0.0), .RTC_MAIN_XTL_MODE("") )  
        \FIC_MSS_0/MSS_ADLIB_INST/INST_MSS_010_IP  (
        .CAN_RXBUS_MGPIO3A_H2F_A(), .CAN_RXBUS_MGPIO3A_H2F_B(), 
        .CAN_TX_EBL_MGPIO4A_H2F_A(), .CAN_TX_EBL_MGPIO4A_H2F_B(), 
        .CAN_TXBUS_MGPIO2A_H2F_A(), .CAN_TXBUS_MGPIO2A_H2F_B(), 
        .CLK_CONFIG_APB(), .COMMS_INT(), .CONFIG_PRESET_N(), 
        .EDAC_ERROR({nc0, nc1, nc2, nc3, nc4, nc5, nc6, nc7}), 
        .F_FM0_RDATA({nc8, nc9, nc10, nc11, nc12, nc13, nc14, nc15, 
        nc16, nc17, nc18, nc19, nc20, nc21, nc22, nc23, nc24, nc25, 
        nc26, nc27, nc28, nc29, nc30, nc31, nc32, nc33, nc34, nc35, 
        nc36, nc37, nc38, nc39}), .F_FM0_READYOUT(), .F_FM0_RESP(), 
        .F_HM0_ADDR({\FIC_MSS_0_FIC_0_APB_MASTER_PADDR[31] , 
        \FIC_MSS_0_FIC_0_APB_MASTER_PADDR[30] , 
        \FIC_MSS_0_FIC_0_APB_MASTER_PADDR[29] , 
        \FIC_MSS_0_FIC_0_APB_MASTER_PADDR[28] , nc40, nc41, nc42, nc43, 
        nc44, nc45, nc46, nc47, nc48, nc49, nc50, nc51, nc52, nc53, 
        nc54, nc55, nc56, nc57, nc58, nc59, 
        \CoreAPB3_0_APBmslave3_PADDR[7] , 
        \CoreAPB3_0_APBmslave3_PADDR[6] , 
        \CoreAPB3_0_APBmslave3_PADDR[5] , 
        \CoreAPB3_0_APBmslave3_PADDR[4] , 
        \CoreAPB3_0_APBmslave3_PADDR[3] , 
        \CoreAPB3_0_APBmslave3_PADDR[2] , 
        \CoreAPB3_0_APBmslave3_PADDR[1] , 
        \CoreAPB3_0_APBmslave3_PADDR[0] }), .F_HM0_ENABLE(
        CoreAPB3_0_APBmslave3_PENABLE), .F_HM0_SEL(
        FIC_MSS_0_FIC_0_APB_MASTER_PSELx), .F_HM0_SIZE({nc60, nc61}), 
        .F_HM0_TRANS1(), .F_HM0_WDATA({
        \CoreAPB3_0_APBmslave3_PWDATA[31] , 
        \CoreAPB3_0_APBmslave3_PWDATA[30] , 
        \CoreAPB3_0_APBmslave3_PWDATA[29] , 
        \CoreAPB3_0_APBmslave3_PWDATA[28] , 
        \CoreAPB3_0_APBmslave3_PWDATA[27] , 
        \CoreAPB3_0_APBmslave3_PWDATA[26] , 
        \CoreAPB3_0_APBmslave3_PWDATA[25] , 
        \CoreAPB3_0_APBmslave3_PWDATA[24] , 
        \CoreAPB3_0_APBmslave3_PWDATA[23] , 
        \CoreAPB3_0_APBmslave3_PWDATA[22] , 
        \CoreAPB3_0_APBmslave3_PWDATA[21] , 
        \CoreAPB3_0_APBmslave3_PWDATA[20] , 
        \CoreAPB3_0_APBmslave3_PWDATA[19] , 
        \CoreAPB3_0_APBmslave3_PWDATA[18] , 
        \CoreAPB3_0_APBmslave3_PWDATA[17] , 
        \CoreAPB3_0_APBmslave3_PWDATA[16] , 
        \CoreAPB3_0_APBmslave3_PWDATA[15] , 
        \CoreAPB3_0_APBmslave3_PWDATA[14] , 
        \CoreAPB3_0_APBmslave3_PWDATA[13] , 
        \CoreAPB3_0_APBmslave3_PWDATA[12] , 
        \CoreAPB3_0_APBmslave3_PWDATA[11] , 
        \CoreAPB3_0_APBmslave3_PWDATA[10] , 
        \CoreAPB3_0_APBmslave3_PWDATA[9] , 
        \CoreAPB3_0_APBmslave3_PWDATA[8] , 
        \CoreAPB3_0_APBmslave3_PWDATA[7] , 
        \CoreAPB3_0_APBmslave3_PWDATA[6] , 
        \CoreAPB3_0_APBmslave3_PWDATA[5] , 
        \CoreAPB3_0_APBmslave3_PWDATA[4] , 
        \CoreAPB3_0_APBmslave3_PWDATA[3] , 
        \CoreAPB3_0_APBmslave3_PWDATA[2] , 
        \CoreAPB3_0_APBmslave3_PWDATA[1] , 
        \CoreAPB3_0_APBmslave3_PWDATA[0] }), .F_HM0_WRITE(
        CoreAPB3_0_APBmslave3_PWRITE), .FAB_CHRGVBUS(), 
        .FAB_DISCHRGVBUS(), .FAB_DMPULLDOWN(), .FAB_DPPULLDOWN(), 
        .FAB_DRVVBUS(), .FAB_IDPULLUP(), .FAB_OPMODE({nc62, nc63}), 
        .FAB_SUSPENDM(), .FAB_TERMSEL(), .FAB_TXVALID(), .FAB_VCONTROL({
        nc64, nc65, nc66, nc67}), .FAB_VCONTROLLOADM(), .FAB_XCVRSEL({
        nc68, nc69}), .FAB_XDATAOUT({nc70, nc71, nc72, nc73, nc74, 
        nc75, nc76, nc77}), .FACC_GLMUX_SEL(), .FIC32_0_MASTER({nc78, 
        nc79}), .FIC32_1_MASTER({nc80, nc81}), .FPGA_RESET_N(), 
        .GTX_CLK(), .H2F_INTERRUPT({nc82, nc83, nc84, nc85, nc86, nc87, 
        nc88, nc89, nc90, nc91, nc92, nc93, nc94, nc95, nc96, nc97}), 
        .H2F_NMI(), .H2FCALIB(), .I2C0_SCL_MGPIO31B_H2F_A(), 
        .I2C0_SCL_MGPIO31B_H2F_B(), .I2C0_SDA_MGPIO30B_H2F_A(), 
        .I2C0_SDA_MGPIO30B_H2F_B(), .I2C1_SCL_MGPIO1A_H2F_A(), 
        .I2C1_SCL_MGPIO1A_H2F_B(), .I2C1_SDA_MGPIO0A_H2F_A(), 
        .I2C1_SDA_MGPIO0A_H2F_B(), .MDCF(), .MDOENF(), .MDOF(), 
        .MMUART0_CTS_MGPIO19B_H2F_A(), .MMUART0_CTS_MGPIO19B_H2F_B(), 
        .MMUART0_DCD_MGPIO22B_H2F_A(), .MMUART0_DCD_MGPIO22B_H2F_B(), 
        .MMUART0_DSR_MGPIO20B_H2F_A(), .MMUART0_DSR_MGPIO20B_H2F_B(), 
        .MMUART0_DTR_MGPIO18B_H2F_A(), .MMUART0_DTR_MGPIO18B_H2F_B(), 
        .MMUART0_RI_MGPIO21B_H2F_A(), .MMUART0_RI_MGPIO21B_H2F_B(), 
        .MMUART0_RTS_MGPIO17B_H2F_A(), .MMUART0_RTS_MGPIO17B_H2F_B(), 
        .MMUART0_RXD_MGPIO28B_H2F_A(), .MMUART0_RXD_MGPIO28B_H2F_B(), 
        .MMUART0_SCK_MGPIO29B_H2F_A(), .MMUART0_SCK_MGPIO29B_H2F_B(), 
        .MMUART0_TXD_MGPIO27B_H2F_A(), .MMUART0_TXD_MGPIO27B_H2F_B(), 
        .MMUART1_DTR_MGPIO12B_H2F_A(), .MMUART1_RTS_MGPIO11B_H2F_A(), 
        .MMUART1_RTS_MGPIO11B_H2F_B(), .MMUART1_RXD_MGPIO26B_H2F_A(), 
        .MMUART1_RXD_MGPIO26B_H2F_B(), .MMUART1_SCK_MGPIO25B_H2F_A(), 
        .MMUART1_SCK_MGPIO25B_H2F_B(), .MMUART1_TXD_MGPIO24B_H2F_A(), 
        .MMUART1_TXD_MGPIO24B_H2F_B(), .MPLL_LOCK(), 
        .PER2_FABRIC_PADDR({nc98, nc99, nc100, nc101, nc102, nc103, 
        nc104, nc105, nc106, nc107, nc108, nc109, nc110, nc111}), 
        .PER2_FABRIC_PENABLE(), .PER2_FABRIC_PSEL(), 
        .PER2_FABRIC_PWDATA({nc112, nc113, nc114, nc115, nc116, nc117, 
        nc118, nc119, nc120, nc121, nc122, nc123, nc124, nc125, nc126, 
        nc127, nc128, nc129, nc130, nc131, nc132, nc133, nc134, nc135, 
        nc136, nc137, nc138, nc139, nc140, nc141, nc142, nc143}), 
        .PER2_FABRIC_PWRITE(), .RTC_MATCH(), .SLEEPDEEP(), 
        .SLEEPHOLDACK(), .SLEEPING(), .SMBALERT_NO0(), .SMBALERT_NO1(), 
        .SMBSUS_NO0(), .SMBSUS_NO1(), .SPI0_CLK_OUT(), 
        .SPI0_SDI_MGPIO5A_H2F_A(), .SPI0_SDI_MGPIO5A_H2F_B(), 
        .SPI0_SDO_MGPIO6A_H2F_A(), .SPI0_SDO_MGPIO6A_H2F_B(), 
        .SPI0_SS0_MGPIO7A_H2F_A(), .SPI0_SS0_MGPIO7A_H2F_B(), 
        .SPI0_SS1_MGPIO8A_H2F_A(), .SPI0_SS1_MGPIO8A_H2F_B(), 
        .SPI0_SS2_MGPIO9A_H2F_A(), .SPI0_SS2_MGPIO9A_H2F_B(), 
        .SPI0_SS3_MGPIO10A_H2F_A(), .SPI0_SS3_MGPIO10A_H2F_B(), 
        .SPI0_SS4_MGPIO19A_H2F_A(), .SPI0_SS5_MGPIO20A_H2F_A(), 
        .SPI0_SS6_MGPIO21A_H2F_A(), .SPI0_SS7_MGPIO22A_H2F_A(), 
        .SPI1_CLK_OUT(), .SPI1_SDI_MGPIO11A_H2F_A(), 
        .SPI1_SDI_MGPIO11A_H2F_B(), .SPI1_SDO_MGPIO12A_H2F_A(), 
        .SPI1_SDO_MGPIO12A_H2F_B(), .SPI1_SS0_MGPIO13A_H2F_A(), 
        .SPI1_SS0_MGPIO13A_H2F_B(), .SPI1_SS1_MGPIO14A_H2F_A(), 
        .SPI1_SS1_MGPIO14A_H2F_B(), .SPI1_SS2_MGPIO15A_H2F_A(), 
        .SPI1_SS2_MGPIO15A_H2F_B(), .SPI1_SS3_MGPIO16A_H2F_A(), 
        .SPI1_SS3_MGPIO16A_H2F_B(), .SPI1_SS4_MGPIO17A_H2F_A(), 
        .SPI1_SS5_MGPIO18A_H2F_A(), .SPI1_SS6_MGPIO23A_H2F_A(), 
        .SPI1_SS7_MGPIO24A_H2F_A(), .TCGF({nc144, nc145, nc146, nc147, 
        nc148, nc149, nc150, nc151, nc152, nc153}), .TRACECLK(), 
        .TRACEDATA({nc154, nc155, nc156, nc157}), .TX_CLK(), .TX_ENF(), 
        .TX_ERRF(), .TXCTL_EN_RIF(), .TXD_RIF({nc158, nc159, nc160, 
        nc161}), .TXDF({nc162, nc163, nc164, nc165, nc166, nc167, 
        nc168, nc169}), .TXEV(), .WDOGTIMEOUT(), .F_ARREADY_HREADYOUT1(
        ), .F_AWREADY_HREADYOUT0(), .F_BID({nc170, nc171, nc172, nc173})
        , .F_BRESP_HRESP0({nc174, nc175}), .F_BVALID(), 
        .F_RDATA_HRDATA01({nc176, nc177, nc178, nc179, nc180, nc181, 
        nc182, nc183, nc184, nc185, nc186, nc187, nc188, nc189, nc190, 
        nc191, nc192, nc193, nc194, nc195, nc196, nc197, nc198, nc199, 
        nc200, nc201, nc202, nc203, nc204, nc205, nc206, nc207, nc208, 
        nc209, nc210, nc211, nc212, nc213, nc214, nc215, nc216, nc217, 
        nc218, nc219, nc220, nc221, nc222, nc223, nc224, nc225, nc226, 
        nc227, nc228, nc229, nc230, nc231, nc232, nc233, nc234, nc235, 
        nc236, nc237, nc238, nc239}), .F_RID({nc240, nc241, nc242, 
        nc243}), .F_RLAST(), .F_RRESP_HRESP1({nc244, nc245}), 
        .F_RVALID(), .F_WREADY(), .MDDR_FABRIC_PRDATA({nc246, nc247, 
        nc248, nc249, nc250, nc251, nc252, nc253, nc254, nc255, nc256, 
        nc257, nc258, nc259, nc260, nc261}), .MDDR_FABRIC_PREADY(), 
        .MDDR_FABRIC_PSLVERR(), .CAN_RXBUS_F2H_SCP(
        \FIC_MSS_0/MSS_ADLIB_INST/CAN_RXBUS_F2H_SCP_net ), 
        .CAN_TX_EBL_F2H_SCP(
        \FIC_MSS_0/MSS_ADLIB_INST/CAN_TX_EBL_F2H_SCP_net ), 
        .CAN_TXBUS_F2H_SCP(
        \FIC_MSS_0/MSS_ADLIB_INST/CAN_TXBUS_F2H_SCP_net ), .COLF(
        \FIC_MSS_0/MSS_ADLIB_INST/COLF_net ), .CRSF(
        \FIC_MSS_0/MSS_ADLIB_INST/CRSF_net ), .F2_DMAREADY({
        \FIC_MSS_0/MSS_ADLIB_INST/F2_DMAREADY_net[1] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F2_DMAREADY_net[0] }), 
        .F2H_INTERRUPT({
        \FIC_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[15] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[14] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[13] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[12] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[11] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[10] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[9] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[8] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[7] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[6] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[5] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[4] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[3] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[2] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[1] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[0] }), .F2HCALIB(
        \FIC_MSS_0/MSS_ADLIB_INST/F2HCALIB_net ), .F_DMAREADY({
        \FIC_MSS_0/MSS_ADLIB_INST/F_DMAREADY_net[1] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_DMAREADY_net[0] }), .F_FM0_ADDR({
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[31] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[30] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[29] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[28] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[27] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[26] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[25] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[24] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[23] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[22] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[21] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[20] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[19] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[18] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[17] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[16] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[15] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[14] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[13] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[12] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[11] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[10] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[9] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[8] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[7] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[6] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[5] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[4] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[3] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[2] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[1] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[0] }), .F_FM0_ENABLE(
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_ENABLE_net ), .F_FM0_MASTLOCK(
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_MASTLOCK_net ), .F_FM0_READY(
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_READY_net ), .F_FM0_SEL(
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_SEL_net ), .F_FM0_SIZE({
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_SIZE_net[1] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_SIZE_net[0] }), .F_FM0_TRANS1(
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_TRANS1_net ), .F_FM0_WDATA({
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[31] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[30] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[29] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[28] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[27] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[26] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[25] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[24] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[23] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[22] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[21] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[20] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[19] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[18] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[17] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[16] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[15] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[14] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[13] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[12] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[11] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[10] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[9] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[8] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[7] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[6] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[5] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[4] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[3] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[2] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[1] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[0] }), .F_FM0_WRITE(
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_WRITE_net ), .F_HM0_RDATA({
        \FIC_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[31] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[30] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[29] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[28] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[27] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[26] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[25] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[24] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[23] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[22] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[21] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[20] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[19] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[18] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[17] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[16] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[15] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[14] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[13] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[12] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[11] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[10] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[9] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[8] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[7] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[6] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[5] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[4] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[3] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[2] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[1] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[0] }), .F_HM0_READY(
        \FIC_MSS_0/MSS_ADLIB_INST/F_HM0_READY_net ), .F_HM0_RESP(
        \FIC_MSS_0/MSS_ADLIB_INST/F_HM0_RESP_net ), .FAB_AVALID(
        \FIC_MSS_0/MSS_ADLIB_INST/FAB_AVALID_net ), .FAB_HOSTDISCON(
        \FIC_MSS_0/MSS_ADLIB_INST/FAB_HOSTDISCON_net ), .FAB_IDDIG(
        \FIC_MSS_0/MSS_ADLIB_INST/FAB_IDDIG_net ), .FAB_LINESTATE({
        \FIC_MSS_0/MSS_ADLIB_INST/FAB_LINESTATE_net[1] , 
        \FIC_MSS_0/MSS_ADLIB_INST/FAB_LINESTATE_net[0] }), 
        .FAB_M3_RESET_N(\FIC_MSS_0/MSS_ADLIB_INST/FAB_M3_RESET_N_net ), 
        .FAB_PLL_LOCK(\FIC_MSS_0/MSS_ADLIB_INST/FAB_PLL_LOCK_net ), 
        .FAB_RXACTIVE(\FIC_MSS_0/MSS_ADLIB_INST/FAB_RXACTIVE_net ), 
        .FAB_RXERROR(\FIC_MSS_0/MSS_ADLIB_INST/FAB_RXERROR_net ), 
        .FAB_RXVALID(\FIC_MSS_0/MSS_ADLIB_INST/FAB_RXVALID_net ), 
        .FAB_RXVALIDH(\FIC_MSS_0/MSS_ADLIB_INST/FAB_RXVALIDH_net ), 
        .FAB_SESSEND(\FIC_MSS_0/MSS_ADLIB_INST/FAB_SESSEND_net ), 
        .FAB_TXREADY(\FIC_MSS_0/MSS_ADLIB_INST/FAB_TXREADY_net ), 
        .FAB_VBUSVALID(\FIC_MSS_0/MSS_ADLIB_INST/FAB_VBUSVALID_net ), 
        .FAB_VSTATUS({\FIC_MSS_0/MSS_ADLIB_INST/FAB_VSTATUS_net[7] , 
        \FIC_MSS_0/MSS_ADLIB_INST/FAB_VSTATUS_net[6] , 
        \FIC_MSS_0/MSS_ADLIB_INST/FAB_VSTATUS_net[5] , 
        \FIC_MSS_0/MSS_ADLIB_INST/FAB_VSTATUS_net[4] , 
        \FIC_MSS_0/MSS_ADLIB_INST/FAB_VSTATUS_net[3] , 
        \FIC_MSS_0/MSS_ADLIB_INST/FAB_VSTATUS_net[2] , 
        \FIC_MSS_0/MSS_ADLIB_INST/FAB_VSTATUS_net[1] , 
        \FIC_MSS_0/MSS_ADLIB_INST/FAB_VSTATUS_net[0] }), .FAB_XDATAIN({
        \FIC_MSS_0/MSS_ADLIB_INST/FAB_XDATAIN_net[7] , 
        \FIC_MSS_0/MSS_ADLIB_INST/FAB_XDATAIN_net[6] , 
        \FIC_MSS_0/MSS_ADLIB_INST/FAB_XDATAIN_net[5] , 
        \FIC_MSS_0/MSS_ADLIB_INST/FAB_XDATAIN_net[4] , 
        \FIC_MSS_0/MSS_ADLIB_INST/FAB_XDATAIN_net[3] , 
        \FIC_MSS_0/MSS_ADLIB_INST/FAB_XDATAIN_net[2] , 
        \FIC_MSS_0/MSS_ADLIB_INST/FAB_XDATAIN_net[1] , 
        \FIC_MSS_0/MSS_ADLIB_INST/FAB_XDATAIN_net[0] }), .GTX_CLKPF(
        \FIC_MSS_0/MSS_ADLIB_INST/GTX_CLKPF_net ), .I2C0_BCLK(
        \FIC_MSS_0/MSS_ADLIB_INST/I2C0_BCLK_net ), .I2C0_SCL_F2H_SCP(
        \FIC_MSS_0/MSS_ADLIB_INST/I2C0_SCL_F2H_SCP_net ), 
        .I2C0_SDA_F2H_SCP(
        \FIC_MSS_0/MSS_ADLIB_INST/I2C0_SDA_F2H_SCP_net ), .I2C1_BCLK(
        \FIC_MSS_0/MSS_ADLIB_INST/I2C1_BCLK_net ), .I2C1_SCL_F2H_SCP(
        \FIC_MSS_0/MSS_ADLIB_INST/I2C1_SCL_F2H_SCP_net ), 
        .I2C1_SDA_F2H_SCP(
        \FIC_MSS_0/MSS_ADLIB_INST/I2C1_SDA_F2H_SCP_net ), .MDIF(
        \FIC_MSS_0/MSS_ADLIB_INST/MDIF_net ), .MGPIO0A_F2H_GPIN(
        \FIC_MSS_0/MSS_ADLIB_INST/MGPIO0A_F2H_GPIN_net ), 
        .MGPIO10A_F2H_GPIN(
        \FIC_MSS_0/MSS_ADLIB_INST/MGPIO10A_F2H_GPIN_net ), 
        .MGPIO11A_F2H_GPIN(
        \FIC_MSS_0/MSS_ADLIB_INST/MGPIO11A_F2H_GPIN_net ), 
        .MGPIO11B_F2H_GPIN(
        \FIC_MSS_0/MSS_ADLIB_INST/MGPIO11B_F2H_GPIN_net ), 
        .MGPIO12A_F2H_GPIN(
        \FIC_MSS_0/MSS_ADLIB_INST/MGPIO12A_F2H_GPIN_net ), 
        .MGPIO13A_F2H_GPIN(
        \FIC_MSS_0/MSS_ADLIB_INST/MGPIO13A_F2H_GPIN_net ), 
        .MGPIO14A_F2H_GPIN(
        \FIC_MSS_0/MSS_ADLIB_INST/MGPIO14A_F2H_GPIN_net ), 
        .MGPIO15A_F2H_GPIN(
        \FIC_MSS_0/MSS_ADLIB_INST/MGPIO15A_F2H_GPIN_net ), 
        .MGPIO16A_F2H_GPIN(
        \FIC_MSS_0/MSS_ADLIB_INST/MGPIO16A_F2H_GPIN_net ), 
        .MGPIO17B_F2H_GPIN(
        \FIC_MSS_0/MSS_ADLIB_INST/MGPIO17B_F2H_GPIN_net ), 
        .MGPIO18B_F2H_GPIN(
        \FIC_MSS_0/MSS_ADLIB_INST/MGPIO18B_F2H_GPIN_net ), 
        .MGPIO19B_F2H_GPIN(
        \FIC_MSS_0/MSS_ADLIB_INST/MGPIO19B_F2H_GPIN_net ), 
        .MGPIO1A_F2H_GPIN(
        \FIC_MSS_0/MSS_ADLIB_INST/MGPIO1A_F2H_GPIN_net ), 
        .MGPIO20B_F2H_GPIN(
        \FIC_MSS_0/MSS_ADLIB_INST/MGPIO20B_F2H_GPIN_net ), 
        .MGPIO21B_F2H_GPIN(
        \FIC_MSS_0/MSS_ADLIB_INST/MGPIO21B_F2H_GPIN_net ), 
        .MGPIO22B_F2H_GPIN(
        \FIC_MSS_0/MSS_ADLIB_INST/MGPIO22B_F2H_GPIN_net ), 
        .MGPIO24B_F2H_GPIN(
        \FIC_MSS_0/MSS_ADLIB_INST/MGPIO24B_F2H_GPIN_net ), 
        .MGPIO25B_F2H_GPIN(
        \FIC_MSS_0/MSS_ADLIB_INST/MGPIO25B_F2H_GPIN_net ), 
        .MGPIO26B_F2H_GPIN(
        \FIC_MSS_0/MSS_ADLIB_INST/MGPIO26B_F2H_GPIN_net ), 
        .MGPIO27B_F2H_GPIN(
        \FIC_MSS_0/MSS_ADLIB_INST/MGPIO27B_F2H_GPIN_net ), 
        .MGPIO28B_F2H_GPIN(
        \FIC_MSS_0/MSS_ADLIB_INST/MGPIO28B_F2H_GPIN_net ), 
        .MGPIO29B_F2H_GPIN(
        \FIC_MSS_0/MSS_ADLIB_INST/MGPIO29B_F2H_GPIN_net ), 
        .MGPIO2A_F2H_GPIN(
        \FIC_MSS_0/MSS_ADLIB_INST/MGPIO2A_F2H_GPIN_net ), 
        .MGPIO30B_F2H_GPIN(
        \FIC_MSS_0/MSS_ADLIB_INST/MGPIO30B_F2H_GPIN_net ), 
        .MGPIO31B_F2H_GPIN(
        \FIC_MSS_0/MSS_ADLIB_INST/MGPIO31B_F2H_GPIN_net ), 
        .MGPIO3A_F2H_GPIN(
        \FIC_MSS_0/MSS_ADLIB_INST/MGPIO3A_F2H_GPIN_net ), 
        .MGPIO4A_F2H_GPIN(
        \FIC_MSS_0/MSS_ADLIB_INST/MGPIO4A_F2H_GPIN_net ), 
        .MGPIO5A_F2H_GPIN(
        \FIC_MSS_0/MSS_ADLIB_INST/MGPIO5A_F2H_GPIN_net ), 
        .MGPIO6A_F2H_GPIN(
        \FIC_MSS_0/MSS_ADLIB_INST/MGPIO6A_F2H_GPIN_net ), 
        .MGPIO7A_F2H_GPIN(
        \FIC_MSS_0/MSS_ADLIB_INST/MGPIO7A_F2H_GPIN_net ), 
        .MGPIO8A_F2H_GPIN(
        \FIC_MSS_0/MSS_ADLIB_INST/MGPIO8A_F2H_GPIN_net ), 
        .MGPIO9A_F2H_GPIN(
        \FIC_MSS_0/MSS_ADLIB_INST/MGPIO9A_F2H_GPIN_net ), 
        .MMUART0_CTS_F2H_SCP(
        \FIC_MSS_0/MSS_ADLIB_INST/MMUART0_CTS_F2H_SCP_net ), 
        .MMUART0_DCD_F2H_SCP(
        \FIC_MSS_0/MSS_ADLIB_INST/MMUART0_DCD_F2H_SCP_net ), 
        .MMUART0_DSR_F2H_SCP(
        \FIC_MSS_0/MSS_ADLIB_INST/MMUART0_DSR_F2H_SCP_net ), 
        .MMUART0_DTR_F2H_SCP(
        \FIC_MSS_0/MSS_ADLIB_INST/MMUART0_DTR_F2H_SCP_net ), 
        .MMUART0_RI_F2H_SCP(
        \FIC_MSS_0/MSS_ADLIB_INST/MMUART0_RI_F2H_SCP_net ), 
        .MMUART0_RTS_F2H_SCP(
        \FIC_MSS_0/MSS_ADLIB_INST/MMUART0_RTS_F2H_SCP_net ), 
        .MMUART0_RXD_F2H_SCP(
        \FIC_MSS_0/MSS_ADLIB_INST/MMUART0_RXD_F2H_SCP_net ), 
        .MMUART0_SCK_F2H_SCP(
        \FIC_MSS_0/MSS_ADLIB_INST/MMUART0_SCK_F2H_SCP_net ), 
        .MMUART0_TXD_F2H_SCP(
        \FIC_MSS_0/MSS_ADLIB_INST/MMUART0_TXD_F2H_SCP_net ), 
        .MMUART1_CTS_F2H_SCP(
        \FIC_MSS_0/MSS_ADLIB_INST/MMUART1_CTS_F2H_SCP_net ), 
        .MMUART1_DCD_F2H_SCP(
        \FIC_MSS_0/MSS_ADLIB_INST/MMUART1_DCD_F2H_SCP_net ), 
        .MMUART1_DSR_F2H_SCP(
        \FIC_MSS_0/MSS_ADLIB_INST/MMUART1_DSR_F2H_SCP_net ), 
        .MMUART1_RI_F2H_SCP(
        \FIC_MSS_0/MSS_ADLIB_INST/MMUART1_RI_F2H_SCP_net ), 
        .MMUART1_RTS_F2H_SCP(
        \FIC_MSS_0/MSS_ADLIB_INST/MMUART1_RTS_F2H_SCP_net ), 
        .MMUART1_RXD_F2H_SCP(
        \FIC_MSS_0/MSS_ADLIB_INST/MMUART1_RXD_F2H_SCP_net ), 
        .MMUART1_SCK_F2H_SCP(
        \FIC_MSS_0/MSS_ADLIB_INST/MMUART1_SCK_F2H_SCP_net ), 
        .MMUART1_TXD_F2H_SCP(
        \FIC_MSS_0/MSS_ADLIB_INST/MMUART1_TXD_F2H_SCP_net ), 
        .PER2_FABRIC_PRDATA({
        \FIC_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[31] , 
        \FIC_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[30] , 
        \FIC_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[29] , 
        \FIC_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[28] , 
        \FIC_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[27] , 
        \FIC_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[26] , 
        \FIC_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[25] , 
        \FIC_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[24] , 
        \FIC_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[23] , 
        \FIC_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[22] , 
        \FIC_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[21] , 
        \FIC_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[20] , 
        \FIC_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[19] , 
        \FIC_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[18] , 
        \FIC_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[17] , 
        \FIC_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[16] , 
        \FIC_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[15] , 
        \FIC_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[14] , 
        \FIC_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[13] , 
        \FIC_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[12] , 
        \FIC_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[11] , 
        \FIC_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[10] , 
        \FIC_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[9] , 
        \FIC_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[8] , 
        \FIC_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[7] , 
        \FIC_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[6] , 
        \FIC_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[5] , 
        \FIC_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[4] , 
        \FIC_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[3] , 
        \FIC_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[2] , 
        \FIC_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[1] , 
        \FIC_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[0] }), 
        .PER2_FABRIC_PREADY(
        \FIC_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PREADY_net ), 
        .PER2_FABRIC_PSLVERR(
        \FIC_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PSLVERR_net ), .RCGF({
        \FIC_MSS_0/MSS_ADLIB_INST/RCGF_net[9] , 
        \FIC_MSS_0/MSS_ADLIB_INST/RCGF_net[8] , 
        \FIC_MSS_0/MSS_ADLIB_INST/RCGF_net[7] , 
        \FIC_MSS_0/MSS_ADLIB_INST/RCGF_net[6] , 
        \FIC_MSS_0/MSS_ADLIB_INST/RCGF_net[5] , 
        \FIC_MSS_0/MSS_ADLIB_INST/RCGF_net[4] , 
        \FIC_MSS_0/MSS_ADLIB_INST/RCGF_net[3] , 
        \FIC_MSS_0/MSS_ADLIB_INST/RCGF_net[2] , 
        \FIC_MSS_0/MSS_ADLIB_INST/RCGF_net[1] , 
        \FIC_MSS_0/MSS_ADLIB_INST/RCGF_net[0] }), .RX_CLKPF(
        \FIC_MSS_0/MSS_ADLIB_INST/RX_CLKPF_net ), .RX_DVF(
        \FIC_MSS_0/MSS_ADLIB_INST/RX_DVF_net ), .RX_ERRF(
        \FIC_MSS_0/MSS_ADLIB_INST/RX_ERRF_net ), .RX_EV(
        \FIC_MSS_0/MSS_ADLIB_INST/RX_EV_net ), .RXDF({
        \FIC_MSS_0/MSS_ADLIB_INST/RXDF_net[7] , 
        \FIC_MSS_0/MSS_ADLIB_INST/RXDF_net[6] , 
        \FIC_MSS_0/MSS_ADLIB_INST/RXDF_net[5] , 
        \FIC_MSS_0/MSS_ADLIB_INST/RXDF_net[4] , 
        \FIC_MSS_0/MSS_ADLIB_INST/RXDF_net[3] , 
        \FIC_MSS_0/MSS_ADLIB_INST/RXDF_net[2] , 
        \FIC_MSS_0/MSS_ADLIB_INST/RXDF_net[1] , 
        \FIC_MSS_0/MSS_ADLIB_INST/RXDF_net[0] }), .SLEEPHOLDREQ(
        \FIC_MSS_0/MSS_ADLIB_INST/SLEEPHOLDREQ_net ), .SMBALERT_NI0(
        \FIC_MSS_0/MSS_ADLIB_INST/SMBALERT_NI0_net ), .SMBALERT_NI1(
        \FIC_MSS_0/MSS_ADLIB_INST/SMBALERT_NI1_net ), .SMBSUS_NI0(
        \FIC_MSS_0/MSS_ADLIB_INST/SMBSUS_NI0_net ), .SMBSUS_NI1(
        \FIC_MSS_0/MSS_ADLIB_INST/SMBSUS_NI1_net ), .SPI0_CLK_IN(
        \FIC_MSS_0/MSS_ADLIB_INST/SPI0_CLK_IN_net ), .SPI0_SDI_F2H_SCP(
        \FIC_MSS_0/MSS_ADLIB_INST/SPI0_SDI_F2H_SCP_net ), 
        .SPI0_SDO_F2H_SCP(
        \FIC_MSS_0/MSS_ADLIB_INST/SPI0_SDO_F2H_SCP_net ), 
        .SPI0_SS0_F2H_SCP(
        \FIC_MSS_0/MSS_ADLIB_INST/SPI0_SS0_F2H_SCP_net ), 
        .SPI0_SS1_F2H_SCP(
        \FIC_MSS_0/MSS_ADLIB_INST/SPI0_SS1_F2H_SCP_net ), 
        .SPI0_SS2_F2H_SCP(
        \FIC_MSS_0/MSS_ADLIB_INST/SPI0_SS2_F2H_SCP_net ), 
        .SPI0_SS3_F2H_SCP(
        \FIC_MSS_0/MSS_ADLIB_INST/SPI0_SS3_F2H_SCP_net ), .SPI1_CLK_IN(
        \FIC_MSS_0/MSS_ADLIB_INST/SPI1_CLK_IN_net ), .SPI1_SDI_F2H_SCP(
        \FIC_MSS_0/MSS_ADLIB_INST/SPI1_SDI_F2H_SCP_net ), 
        .SPI1_SDO_F2H_SCP(
        \FIC_MSS_0/MSS_ADLIB_INST/SPI1_SDO_F2H_SCP_net ), 
        .SPI1_SS0_F2H_SCP(
        \FIC_MSS_0/MSS_ADLIB_INST/SPI1_SS0_F2H_SCP_net ), 
        .SPI1_SS1_F2H_SCP(
        \FIC_MSS_0/MSS_ADLIB_INST/SPI1_SS1_F2H_SCP_net ), 
        .SPI1_SS2_F2H_SCP(
        \FIC_MSS_0/MSS_ADLIB_INST/SPI1_SS2_F2H_SCP_net ), 
        .SPI1_SS3_F2H_SCP(
        \FIC_MSS_0/MSS_ADLIB_INST/SPI1_SS3_F2H_SCP_net ), .TX_CLKPF(
        \FIC_MSS_0/MSS_ADLIB_INST/TX_CLKPF_net ), 
        .USER_MSS_GPIO_RESET_N(
        \FIC_MSS_0/MSS_ADLIB_INST/USER_MSS_GPIO_RESET_N_net ), 
        .USER_MSS_RESET_N(
        \FIC_MSS_0/MSS_ADLIB_INST/USER_MSS_RESET_N_net ), .XCLK_FAB(
        \FIC_MSS_0/MSS_ADLIB_INST/XCLK_FAB_net ), .CLK_BASE(
        \FIC_MSS_0/MSS_ADLIB_INST/CLK_BASE_net ), .CLK_MDDR_APB(
        \FIC_MSS_0/MSS_ADLIB_INST/CLK_MDDR_APB_net ), .F_ARADDR_HADDR1({
        \FIC_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[31] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[30] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[29] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[28] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[27] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[26] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[25] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[24] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[23] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[22] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[21] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[20] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[19] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[18] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[17] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[16] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[15] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[14] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[13] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[12] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[11] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[10] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[9] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[8] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[7] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[6] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[5] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[4] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[3] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[2] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[1] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[0] }), 
        .F_ARBURST_HTRANS1({
        \FIC_MSS_0/MSS_ADLIB_INST/F_ARBURST_HTRANS1_net[1] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_ARBURST_HTRANS1_net[0] }), 
        .F_ARID_HSEL1({\FIC_MSS_0/MSS_ADLIB_INST/F_ARID_HSEL1_net[3] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_ARID_HSEL1_net[2] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_ARID_HSEL1_net[1] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_ARID_HSEL1_net[0] }), 
        .F_ARLEN_HBURST1({
        \FIC_MSS_0/MSS_ADLIB_INST/F_ARLEN_HBURST1_net[3] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_ARLEN_HBURST1_net[2] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_ARLEN_HBURST1_net[1] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_ARLEN_HBURST1_net[0] }), 
        .F_ARLOCK_HMASTLOCK1({
        \FIC_MSS_0/MSS_ADLIB_INST/F_ARLOCK_HMASTLOCK1_net[1] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_ARLOCK_HMASTLOCK1_net[0] }), 
        .F_ARSIZE_HSIZE1({
        \FIC_MSS_0/MSS_ADLIB_INST/F_ARSIZE_HSIZE1_net[1] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_ARSIZE_HSIZE1_net[0] }), 
        .F_ARVALID_HWRITE1(
        \FIC_MSS_0/MSS_ADLIB_INST/F_ARVALID_HWRITE1_net ), 
        .F_AWADDR_HADDR0({
        \FIC_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[31] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[30] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[29] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[28] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[27] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[26] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[25] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[24] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[23] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[22] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[21] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[20] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[19] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[18] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[17] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[16] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[15] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[14] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[13] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[12] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[11] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[10] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[9] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[8] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[7] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[6] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[5] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[4] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[3] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[2] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[1] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[0] }), 
        .F_AWBURST_HTRANS0({
        \FIC_MSS_0/MSS_ADLIB_INST/F_AWBURST_HTRANS0_net[1] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_AWBURST_HTRANS0_net[0] }), 
        .F_AWID_HSEL0({\FIC_MSS_0/MSS_ADLIB_INST/F_AWID_HSEL0_net[3] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_AWID_HSEL0_net[2] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_AWID_HSEL0_net[1] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_AWID_HSEL0_net[0] }), 
        .F_AWLEN_HBURST0({
        \FIC_MSS_0/MSS_ADLIB_INST/F_AWLEN_HBURST0_net[3] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_AWLEN_HBURST0_net[2] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_AWLEN_HBURST0_net[1] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_AWLEN_HBURST0_net[0] }), 
        .F_AWLOCK_HMASTLOCK0({
        \FIC_MSS_0/MSS_ADLIB_INST/F_AWLOCK_HMASTLOCK0_net[1] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_AWLOCK_HMASTLOCK0_net[0] }), 
        .F_AWSIZE_HSIZE0({
        \FIC_MSS_0/MSS_ADLIB_INST/F_AWSIZE_HSIZE0_net[1] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_AWSIZE_HSIZE0_net[0] }), 
        .F_AWVALID_HWRITE0(
        \FIC_MSS_0/MSS_ADLIB_INST/F_AWVALID_HWRITE0_net ), .F_BREADY(
        \FIC_MSS_0/MSS_ADLIB_INST/F_BREADY_net ), .F_RMW_AXI(
        \FIC_MSS_0/MSS_ADLIB_INST/F_RMW_AXI_net ), .F_RREADY(
        \FIC_MSS_0/MSS_ADLIB_INST/F_RREADY_net ), .F_WDATA_HWDATA01({
        \FIC_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[63] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[62] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[61] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[60] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[59] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[58] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[57] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[56] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[55] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[54] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[53] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[52] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[51] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[50] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[49] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[48] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[47] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[46] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[45] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[44] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[43] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[42] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[41] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[40] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[39] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[38] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[37] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[36] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[35] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[34] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[33] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[32] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[31] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[30] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[29] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[28] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[27] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[26] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[25] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[24] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[23] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[22] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[21] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[20] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[19] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[18] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[17] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[16] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[15] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[14] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[13] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[12] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[11] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[10] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[9] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[8] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[7] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[6] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[5] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[4] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[3] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[2] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[1] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[0] }), 
        .F_WID_HREADY01({
        \FIC_MSS_0/MSS_ADLIB_INST/F_WID_HREADY01_net[3] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_WID_HREADY01_net[2] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_WID_HREADY01_net[1] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_WID_HREADY01_net[0] }), .F_WLAST(
        \FIC_MSS_0/MSS_ADLIB_INST/F_WLAST_net ), .F_WSTRB({
        \FIC_MSS_0/MSS_ADLIB_INST/F_WSTRB_net[7] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_WSTRB_net[6] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_WSTRB_net[5] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_WSTRB_net[4] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_WSTRB_net[3] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_WSTRB_net[2] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_WSTRB_net[1] , 
        \FIC_MSS_0/MSS_ADLIB_INST/F_WSTRB_net[0] }), .F_WVALID(
        \FIC_MSS_0/MSS_ADLIB_INST/F_WVALID_net ), .FPGA_MDDR_ARESET_N(
        \FIC_MSS_0/MSS_ADLIB_INST/FPGA_MDDR_ARESET_N_net ), 
        .MDDR_FABRIC_PADDR({
        \FIC_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PADDR_net[10] , 
        \FIC_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PADDR_net[9] , 
        \FIC_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PADDR_net[8] , 
        \FIC_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PADDR_net[7] , 
        \FIC_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PADDR_net[6] , 
        \FIC_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PADDR_net[5] , 
        \FIC_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PADDR_net[4] , 
        \FIC_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PADDR_net[3] , 
        \FIC_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PADDR_net[2] }), 
        .MDDR_FABRIC_PENABLE(
        \FIC_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PENABLE_net ), 
        .MDDR_FABRIC_PSEL(
        \FIC_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PSEL_net ), 
        .MDDR_FABRIC_PWDATA({
        \FIC_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[15] , 
        \FIC_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[14] , 
        \FIC_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[13] , 
        \FIC_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[12] , 
        \FIC_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[11] , 
        \FIC_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[10] , 
        \FIC_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[9] , 
        \FIC_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[8] , 
        \FIC_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[7] , 
        \FIC_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[6] , 
        \FIC_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[5] , 
        \FIC_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[4] , 
        \FIC_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[3] , 
        \FIC_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[2] , 
        \FIC_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[1] , 
        \FIC_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[0] }), 
        .MDDR_FABRIC_PWRITE(
        \FIC_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWRITE_net ), .PRESET_N(
        \FIC_MSS_0/MSS_ADLIB_INST/PRESET_N_net ), 
        .CAN_RXBUS_USBA_DATA1_MGPIO3A_IN(GND), 
        .CAN_TX_EBL_USBA_DATA2_MGPIO4A_IN(GND), 
        .CAN_TXBUS_USBA_DATA0_MGPIO2A_IN(GND), .DM_IN({GND, 
        \FIC_MSS_0/MDDR_DM_RDQS_1_PAD_Y , 
        \FIC_MSS_0/MDDR_DM_RDQS_0_PAD_Y }), .DRAM_DQ_IN({GND, GND, 
        \FIC_MSS_0/MDDR_DQ_15_PAD_Y , \FIC_MSS_0/MDDR_DQ_14_PAD_Y , 
        \FIC_MSS_0/MDDR_DQ_13_PAD_Y , \FIC_MSS_0/MDDR_DQ_12_PAD_Y , 
        \FIC_MSS_0/MDDR_DQ_11_PAD_Y , \FIC_MSS_0/MDDR_DQ_10_PAD_Y , 
        \FIC_MSS_0/MDDR_DQ_9_PAD_Y , \FIC_MSS_0/MDDR_DQ_8_PAD_Y , 
        \FIC_MSS_0/MDDR_DQ_7_PAD_Y , \FIC_MSS_0/MDDR_DQ_6_PAD_Y , 
        \FIC_MSS_0/MDDR_DQ_5_PAD_Y , \FIC_MSS_0/MDDR_DQ_4_PAD_Y , 
        \FIC_MSS_0/MDDR_DQ_3_PAD_Y , \FIC_MSS_0/MDDR_DQ_2_PAD_Y , 
        \FIC_MSS_0/MDDR_DQ_1_PAD_Y , \FIC_MSS_0/MDDR_DQ_0_PAD_Y }), 
        .DRAM_DQS_IN({GND, \FIC_MSS_0/MDDR_DQS_1_PAD_Y , 
        \FIC_MSS_0/MDDR_DQS_0_PAD_Y }), .DRAM_FIFO_WE_IN({GND, 
        \FIC_MSS_0/MDDR_DQS_TMATCH_0_IN_PAD_Y }), 
        .I2C0_SCL_USBC_DATA1_MGPIO31B_IN(GND), 
        .I2C0_SDA_USBC_DATA0_MGPIO30B_IN(GND), 
        .I2C1_SCL_USBA_DATA4_MGPIO1A_IN(GND), 
        .I2C1_SDA_USBA_DATA3_MGPIO0A_IN(GND), 
        .MMUART0_CTS_USBC_DATA7_MGPIO19B_IN(GND), 
        .MMUART0_DCD_MGPIO22B_IN(GND), .MMUART0_DSR_MGPIO20B_IN(GND), 
        .MMUART0_DTR_USBC_DATA6_MGPIO18B_IN(GND), 
        .MMUART0_RI_MGPIO21B_IN(GND), 
        .MMUART0_RTS_USBC_DATA5_MGPIO17B_IN(GND), 
        .MMUART0_RXD_USBC_STP_MGPIO28B_IN(
        \FIC_MSS_0/MMUART_0_RXD_PAD_Y ), 
        .MMUART0_SCK_USBC_NXT_MGPIO29B_IN(GND), 
        .MMUART0_TXD_USBC_DIR_MGPIO27B_IN(GND), 
        .MMUART1_RXD_USBC_DATA3_MGPIO26B_IN(GND), 
        .MMUART1_SCK_USBC_DATA4_MGPIO25B_IN(GND), 
        .MMUART1_TXD_USBC_DATA2_MGPIO24B_IN(GND), 
        .RGMII_GTX_CLK_RMII_CLK_USBB_XCLK_IN(GND), 
        .RGMII_MDC_RMII_MDC_IN(GND), 
        .RGMII_MDIO_RMII_MDIO_USBB_DATA7_IN(GND), .RGMII_RX_CLK_IN(GND)
        , .RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_IN(GND), 
        .RGMII_RXD0_RMII_RXD0_USBB_DATA0_IN(GND), 
        .RGMII_RXD1_RMII_RXD1_USBB_DATA1_IN(GND), 
        .RGMII_RXD2_RMII_RX_ER_USBB_DATA3_IN(GND), 
        .RGMII_RXD3_USBB_DATA4_IN(GND), .RGMII_TX_CLK_IN(GND), 
        .RGMII_TX_CTL_RMII_TX_EN_USBB_NXT_IN(GND), 
        .RGMII_TXD0_RMII_TXD0_USBB_DIR_IN(GND), 
        .RGMII_TXD1_RMII_TXD1_USBB_STP_IN(GND), 
        .RGMII_TXD2_USBB_DATA5_IN(GND), .RGMII_TXD3_USBB_DATA6_IN(GND), 
        .SPI0_SCK_USBA_XCLK_IN(GND), .SPI0_SDI_USBA_DIR_MGPIO5A_IN(GND)
        , .SPI0_SDO_USBA_STP_MGPIO6A_IN(GND), 
        .SPI0_SS0_USBA_NXT_MGPIO7A_IN(GND), 
        .SPI0_SS1_USBA_DATA5_MGPIO8A_IN(GND), 
        .SPI0_SS2_USBA_DATA6_MGPIO9A_IN(GND), 
        .SPI0_SS3_USBA_DATA7_MGPIO10A_IN(GND), .SPI1_SCK_IN(GND), 
        .SPI1_SDI_MGPIO11A_IN(GND), .SPI1_SDO_MGPIO12A_IN(GND), 
        .SPI1_SS0_MGPIO13A_IN(GND), .SPI1_SS1_MGPIO14A_IN(GND), 
        .SPI1_SS2_MGPIO15A_IN(GND), .SPI1_SS3_MGPIO16A_IN(GND), 
        .SPI1_SS4_MGPIO17A_IN(GND), .SPI1_SS5_MGPIO18A_IN(GND), 
        .SPI1_SS6_MGPIO23A_IN(GND), .SPI1_SS7_MGPIO24A_IN(GND), 
        .USBC_XCLK_IN(GND), .CAN_RXBUS_USBA_DATA1_MGPIO3A_OUT(), 
        .CAN_TX_EBL_USBA_DATA2_MGPIO4A_OUT(), 
        .CAN_TXBUS_USBA_DATA0_MGPIO2A_OUT(), .DRAM_ADDR({
        \FIC_MSS_0/DRAM_ADDR_net_0[15] , 
        \FIC_MSS_0/DRAM_ADDR_net_0[14] , 
        \FIC_MSS_0/DRAM_ADDR_net_0[13] , 
        \FIC_MSS_0/DRAM_ADDR_net_0[12] , 
        \FIC_MSS_0/DRAM_ADDR_net_0[11] , 
        \FIC_MSS_0/DRAM_ADDR_net_0[10] , 
        \FIC_MSS_0/DRAM_ADDR_net_0[9] , \FIC_MSS_0/DRAM_ADDR_net_0[8] , 
        \FIC_MSS_0/DRAM_ADDR_net_0[7] , \FIC_MSS_0/DRAM_ADDR_net_0[6] , 
        \FIC_MSS_0/DRAM_ADDR_net_0[5] , \FIC_MSS_0/DRAM_ADDR_net_0[4] , 
        \FIC_MSS_0/DRAM_ADDR_net_0[3] , \FIC_MSS_0/DRAM_ADDR_net_0[2] , 
        \FIC_MSS_0/DRAM_ADDR_net_0[1] , \FIC_MSS_0/DRAM_ADDR_net_0[0] })
        , .DRAM_BA({\FIC_MSS_0/DRAM_BA_net_0[2] , 
        \FIC_MSS_0/DRAM_BA_net_0[1] , \FIC_MSS_0/DRAM_BA_net_0[0] }), 
        .DRAM_CASN(\FIC_MSS_0/MSS_ADLIB_INST_DRAM_CASN ), .DRAM_CKE(
        \FIC_MSS_0/MSS_ADLIB_INST_DRAM_CKE ), .DRAM_CLK(
        \FIC_MSS_0/MSS_ADLIB_INST_DRAM_CLK ), .DRAM_CSN(
        \FIC_MSS_0/MSS_ADLIB_INST_DRAM_CSN ), .DRAM_DM_RDQS_OUT({nc262, 
        \FIC_MSS_0/DRAM_DM_RDQS_OUT_net_0[1] , 
        \FIC_MSS_0/DRAM_DM_RDQS_OUT_net_0[0] }), .DRAM_DQ_OUT({nc263, 
        nc264, \FIC_MSS_0/DRAM_DQ_OUT_net_0[15] , 
        \FIC_MSS_0/DRAM_DQ_OUT_net_0[14] , 
        \FIC_MSS_0/DRAM_DQ_OUT_net_0[13] , 
        \FIC_MSS_0/DRAM_DQ_OUT_net_0[12] , 
        \FIC_MSS_0/DRAM_DQ_OUT_net_0[11] , 
        \FIC_MSS_0/DRAM_DQ_OUT_net_0[10] , 
        \FIC_MSS_0/DRAM_DQ_OUT_net_0[9] , 
        \FIC_MSS_0/DRAM_DQ_OUT_net_0[8] , 
        \FIC_MSS_0/DRAM_DQ_OUT_net_0[7] , 
        \FIC_MSS_0/DRAM_DQ_OUT_net_0[6] , 
        \FIC_MSS_0/DRAM_DQ_OUT_net_0[5] , 
        \FIC_MSS_0/DRAM_DQ_OUT_net_0[4] , 
        \FIC_MSS_0/DRAM_DQ_OUT_net_0[3] , 
        \FIC_MSS_0/DRAM_DQ_OUT_net_0[2] , 
        \FIC_MSS_0/DRAM_DQ_OUT_net_0[1] , 
        \FIC_MSS_0/DRAM_DQ_OUT_net_0[0] }), .DRAM_DQS_OUT({nc265, 
        \FIC_MSS_0/DRAM_DQS_OUT_net_0[1] , 
        \FIC_MSS_0/DRAM_DQS_OUT_net_0[0] }), .DRAM_FIFO_WE_OUT({nc266, 
        \FIC_MSS_0/DRAM_FIFO_WE_OUT_net_0[0] }), .DRAM_ODT(
        \FIC_MSS_0/MSS_ADLIB_INST_DRAM_ODT ), .DRAM_RASN(
        \FIC_MSS_0/MSS_ADLIB_INST_DRAM_RASN ), .DRAM_RSTN(
        \FIC_MSS_0/MSS_ADLIB_INST_DRAM_RSTN ), .DRAM_WEN(
        \FIC_MSS_0/MSS_ADLIB_INST_DRAM_WEN ), 
        .I2C0_SCL_USBC_DATA1_MGPIO31B_OUT(), 
        .I2C0_SDA_USBC_DATA0_MGPIO30B_OUT(), 
        .I2C1_SCL_USBA_DATA4_MGPIO1A_OUT(), 
        .I2C1_SDA_USBA_DATA3_MGPIO0A_OUT(), 
        .MMUART0_CTS_USBC_DATA7_MGPIO19B_OUT(), 
        .MMUART0_DCD_MGPIO22B_OUT(), .MMUART0_DSR_MGPIO20B_OUT(), 
        .MMUART0_DTR_USBC_DATA6_MGPIO18B_OUT(), 
        .MMUART0_RI_MGPIO21B_OUT(), 
        .MMUART0_RTS_USBC_DATA5_MGPIO17B_OUT(), 
        .MMUART0_RXD_USBC_STP_MGPIO28B_OUT(), 
        .MMUART0_SCK_USBC_NXT_MGPIO29B_OUT(), 
        .MMUART0_TXD_USBC_DIR_MGPIO27B_OUT(
        \FIC_MSS_0/MSS_ADLIB_INST_MMUART0_TXD_USBC_DIR_MGPIO27B_OUT ), 
        .MMUART1_RXD_USBC_DATA3_MGPIO26B_OUT(), 
        .MMUART1_SCK_USBC_DATA4_MGPIO25B_OUT(), 
        .MMUART1_TXD_USBC_DATA2_MGPIO24B_OUT(), 
        .RGMII_GTX_CLK_RMII_CLK_USBB_XCLK_OUT(), 
        .RGMII_MDC_RMII_MDC_OUT(), 
        .RGMII_MDIO_RMII_MDIO_USBB_DATA7_OUT(), .RGMII_RX_CLK_OUT(), 
        .RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_OUT(), 
        .RGMII_RXD0_RMII_RXD0_USBB_DATA0_OUT(), 
        .RGMII_RXD1_RMII_RXD1_USBB_DATA1_OUT(), 
        .RGMII_RXD2_RMII_RX_ER_USBB_DATA3_OUT(), 
        .RGMII_RXD3_USBB_DATA4_OUT(), .RGMII_TX_CLK_OUT(), 
        .RGMII_TX_CTL_RMII_TX_EN_USBB_NXT_OUT(), 
        .RGMII_TXD0_RMII_TXD0_USBB_DIR_OUT(), 
        .RGMII_TXD1_RMII_TXD1_USBB_STP_OUT(), 
        .RGMII_TXD2_USBB_DATA5_OUT(), .RGMII_TXD3_USBB_DATA6_OUT(), 
        .SPI0_SCK_USBA_XCLK_OUT(), .SPI0_SDI_USBA_DIR_MGPIO5A_OUT(), 
        .SPI0_SDO_USBA_STP_MGPIO6A_OUT(), 
        .SPI0_SS0_USBA_NXT_MGPIO7A_OUT(), 
        .SPI0_SS1_USBA_DATA5_MGPIO8A_OUT(), 
        .SPI0_SS2_USBA_DATA6_MGPIO9A_OUT(), 
        .SPI0_SS3_USBA_DATA7_MGPIO10A_OUT(), .SPI1_SCK_OUT(), 
        .SPI1_SDI_MGPIO11A_OUT(), .SPI1_SDO_MGPIO12A_OUT(), 
        .SPI1_SS0_MGPIO13A_OUT(), .SPI1_SS1_MGPIO14A_OUT(), 
        .SPI1_SS2_MGPIO15A_OUT(), .SPI1_SS3_MGPIO16A_OUT(), 
        .SPI1_SS4_MGPIO17A_OUT(), .SPI1_SS5_MGPIO18A_OUT(), 
        .SPI1_SS6_MGPIO23A_OUT(), .SPI1_SS7_MGPIO24A_OUT(), 
        .USBC_XCLK_OUT(), .CAN_RXBUS_USBA_DATA1_MGPIO3A_OE(), 
        .CAN_TX_EBL_USBA_DATA2_MGPIO4A_OE(), 
        .CAN_TXBUS_USBA_DATA0_MGPIO2A_OE(), .DM_OE({nc267, 
        \FIC_MSS_0/DM_OE_net_0[1] , \FIC_MSS_0/DM_OE_net_0[0] }), 
        .DRAM_DQ_OE({nc268, nc269, \FIC_MSS_0/DRAM_DQ_OE_net_0[15] , 
        \FIC_MSS_0/DRAM_DQ_OE_net_0[14] , 
        \FIC_MSS_0/DRAM_DQ_OE_net_0[13] , 
        \FIC_MSS_0/DRAM_DQ_OE_net_0[12] , 
        \FIC_MSS_0/DRAM_DQ_OE_net_0[11] , 
        \FIC_MSS_0/DRAM_DQ_OE_net_0[10] , 
        \FIC_MSS_0/DRAM_DQ_OE_net_0[9] , 
        \FIC_MSS_0/DRAM_DQ_OE_net_0[8] , 
        \FIC_MSS_0/DRAM_DQ_OE_net_0[7] , 
        \FIC_MSS_0/DRAM_DQ_OE_net_0[6] , 
        \FIC_MSS_0/DRAM_DQ_OE_net_0[5] , 
        \FIC_MSS_0/DRAM_DQ_OE_net_0[4] , 
        \FIC_MSS_0/DRAM_DQ_OE_net_0[3] , 
        \FIC_MSS_0/DRAM_DQ_OE_net_0[2] , 
        \FIC_MSS_0/DRAM_DQ_OE_net_0[1] , 
        \FIC_MSS_0/DRAM_DQ_OE_net_0[0] }), .DRAM_DQS_OE({nc270, 
        \FIC_MSS_0/DRAM_DQS_OE_net_0[1] , 
        \FIC_MSS_0/DRAM_DQS_OE_net_0[0] }), 
        .I2C0_SCL_USBC_DATA1_MGPIO31B_OE(), 
        .I2C0_SDA_USBC_DATA0_MGPIO30B_OE(), 
        .I2C1_SCL_USBA_DATA4_MGPIO1A_OE(), 
        .I2C1_SDA_USBA_DATA3_MGPIO0A_OE(), 
        .MMUART0_CTS_USBC_DATA7_MGPIO19B_OE(), 
        .MMUART0_DCD_MGPIO22B_OE(), .MMUART0_DSR_MGPIO20B_OE(), 
        .MMUART0_DTR_USBC_DATA6_MGPIO18B_OE(), .MMUART0_RI_MGPIO21B_OE(
        ), .MMUART0_RTS_USBC_DATA5_MGPIO17B_OE(), 
        .MMUART0_RXD_USBC_STP_MGPIO28B_OE(), 
        .MMUART0_SCK_USBC_NXT_MGPIO29B_OE(), 
        .MMUART0_TXD_USBC_DIR_MGPIO27B_OE(
        \FIC_MSS_0/MSS_ADLIB_INST_MMUART0_TXD_USBC_DIR_MGPIO27B_OE ), 
        .MMUART1_RXD_USBC_DATA3_MGPIO26B_OE(), 
        .MMUART1_SCK_USBC_DATA4_MGPIO25B_OE(), 
        .MMUART1_TXD_USBC_DATA2_MGPIO24B_OE(), 
        .RGMII_GTX_CLK_RMII_CLK_USBB_XCLK_OE(), .RGMII_MDC_RMII_MDC_OE(
        ), .RGMII_MDIO_RMII_MDIO_USBB_DATA7_OE(), .RGMII_RX_CLK_OE(), 
        .RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_OE(), 
        .RGMII_RXD0_RMII_RXD0_USBB_DATA0_OE(), 
        .RGMII_RXD1_RMII_RXD1_USBB_DATA1_OE(), 
        .RGMII_RXD2_RMII_RX_ER_USBB_DATA3_OE(), 
        .RGMII_RXD3_USBB_DATA4_OE(), .RGMII_TX_CLK_OE(), 
        .RGMII_TX_CTL_RMII_TX_EN_USBB_NXT_OE(), 
        .RGMII_TXD0_RMII_TXD0_USBB_DIR_OE(), 
        .RGMII_TXD1_RMII_TXD1_USBB_STP_OE(), .RGMII_TXD2_USBB_DATA5_OE(
        ), .RGMII_TXD3_USBB_DATA6_OE(), .SPI0_SCK_USBA_XCLK_OE(), 
        .SPI0_SDI_USBA_DIR_MGPIO5A_OE(), .SPI0_SDO_USBA_STP_MGPIO6A_OE(
        ), .SPI0_SS0_USBA_NXT_MGPIO7A_OE(), 
        .SPI0_SS1_USBA_DATA5_MGPIO8A_OE(), 
        .SPI0_SS2_USBA_DATA6_MGPIO9A_OE(), 
        .SPI0_SS3_USBA_DATA7_MGPIO10A_OE(), .SPI1_SCK_OE(), 
        .SPI1_SDI_MGPIO11A_OE(), .SPI1_SDO_MGPIO12A_OE(), 
        .SPI1_SS0_MGPIO13A_OE(), .SPI1_SS1_MGPIO14A_OE(), 
        .SPI1_SS2_MGPIO15A_OE(), .SPI1_SS3_MGPIO16A_OE(), 
        .SPI1_SS4_MGPIO17A_OE(), .SPI1_SS5_MGPIO18A_OE(), 
        .SPI1_SS6_MGPIO23A_OE(), .SPI1_SS7_MGPIO24A_OE(), 
        .USBC_XCLK_OE());
    CFG4 #( .INIT(16'hAA08) )  
        \CoreGPIO_0/xhdl1.GEN_BITS[4].APB_32.edge_both_65_iv_i_0[4]  (
        .A(\CoreGPIO_0/CONFIG_reg[4][3] ), .B(
        \CoreGPIO_0/edge_both[4] ), .C(
        \CoreAPB3_0_APBmslave3_PWDATA[4] ), .D(\CoreGPIO_0/N_143_i ), 
        .Y(\CoreGPIO_0/N_91 ));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_166_rs_RNI4KVK  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_67_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_166_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_4_rs[5] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_4_[5]_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_130_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_84_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_130_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_130_rs_net_1 ));
    CFG4 #( .INIT(16'hF2F3) )  
        \CoreGPIO_0/xhdl1.GEN_BITS[16].APB_32.INTR_reg_217_0_o2_1_0[16]  
        (.A(\CoreGPIO_0/CONFIG_reg[16][6] ), .B(
        \CoreGPIO_0/edge_neg[16] ), .C(
        \CoreGPIO_0/INTR_reg_217_0_o2_0[16] ), .D(
        \CoreGPIO_0/CONFIG_reg[16][5] ), .Y(
        \CoreGPIO_0/INTR_reg_217_0_o2_1[16] ));
    IOIN_IB \FIC_MSS_0/MMUART_0_RXD_PAD/U_IOIN  (.YIN(
        \FIC_MSS_0/MMUART_0_RXD_PAD/YIN ), .E(GND), .Y());
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_245_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_117_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_245_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_245_rs_net_1 ));
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_31  (
        .A(\reg_apb_wrp_0/reg16x8_0/mem_6_[1]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_493 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_31_net_1 ));
    CFG2 #( .INIT(4'h6) )  \CoreGPIO_0/edge_both_2_sqmuxa_15_i_x2  (.A(
        \CoreGPIO_0/gpin2[0] ), .B(
        \CoreGPIO_0.xhdl1.GEN_BITS[0].gpin3[0] ), .Y(
        \CoreGPIO_0/N_141_i ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_275  (.A(GND), 
        .B(GND), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/F_ARLEN_HBURST1_net[3] ), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/PRESET_N_net ), .IPC());
    sdf_IOPAD_TRI \FIC_MSS_0/MDDR_CAS_N_PAD/U_IOPAD  (.PAD(MDDR_CAS_N), 
        .D(\FIC_MSS_0/MSS_ADLIB_INST_DRAM_CASN ), .E(
        \FIC_MSS_0/MDDR_CAS_N_PAD/EOUT ));
    CFG4 #( .INIT(16'hEC00) )  \CoreAPB3_0/u_mux_p_to_b3/PRDATA[19]  (
        .A(\CoreGPIO_0.xhdl1.GEN_BITS[0].APB_32.GPOUT_reg9 ), .B(
        \CoreGPIO_0.N_548 ), .C(
        \CoreGPIO_0.xhdl1.GEN_BITS[19].APB_32.GPOUT_reg[19] ), .D(
        CoreAPB3_0_APBmslave5_PSELx), .Y(
        \FIC_MSS_0_FIC_0_APB_MASTER_PRDATA[19] ));
    CFG4 #( .INIT(16'h4657) )  
        \CoreGPIO_0/CONFIG_reg_o_2_31_bm_1_1[4]  (.A(
        \CoreAPB3_0_APBmslave3_PADDR[4] ), .B(
        \CoreAPB3_0_APBmslave3_PADDR[3] ), .C(
        \CoreGPIO_0/CONFIG_reg_o_2_31_bm_1_1_RNO[4]_net_1 ), .D(
        \CoreGPIO_0/CONFIG_reg_o_2_31_bm_1_RNO_0[4]_net_1 ), .Y(
        \CoreGPIO_0/CONFIG_reg_o_2_31_bm_1[4] ));
    CFG3 #( .INIT(8'hF2) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_237  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_13_[5]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_500 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_237_i ));
    INV_BA AFLSDF_INV_53 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_3_net_1 ), .Y(
        AFLSDF_INV_53_net_1));
    CFG4 #( .INIT(16'hAC0F) )  
        \CoreGPIO_0/CONFIG_reg_o_2_31_bm_RNO_0[5]  (.A(
        \CoreGPIO_0/CONFIG_reg[15][5] ), .B(
        \CoreGPIO_0/CONFIG_reg[31][5] ), .C(
        \CoreGPIO_0/CONFIG_reg_o_2_28_1_1[5] ), .D(
        \CoreAPB3_0_APBmslave3_PADDR[5] ), .Y(
        \CoreGPIO_0/CONFIG_reg_o_2_31_bm_RNO_0[5]_net_1 ));
    CFG3 #( .INIT(8'hF2) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_231  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_12_[7]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_495 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_231_i ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_98  (.A(VCC), 
        .B(VCC), .C(VCC), .IPA(\FIC_MSS_0/MSS_ADLIB_INST/MDIF_net ), 
        .IPB(), .IPC());
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_242_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_114_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_242_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_242_rs_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_122_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB15_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_3__1_sqmuxa ), .ALn(
        AFLSDF_INV_21_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(GND)
        , .Q(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_122_set_net_1 ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_20  (.A(
        \FIC_MSS_0_FIC_0_APB_MASTER_PRDATA[25] ), .B(GND), .C(VCC), 
        .IPA(\FIC_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[25] ), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_MASTLOCK_net ), .IPC());
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[24].REG_GEN.CONFIG_reg[24][3]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[3] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB11_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[24]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB1_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[24][3] ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_233_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_105_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_233_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_233_rs_net_1 ));
    CFG3 #( .INIT(8'hF2) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_146  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_2_[2]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_501 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_146_i ));
    CFG4 #( .INIT(16'h0F35) )  
        \CoreGPIO_0/CONFIG_reg_o_2_31_am_1_RNO_2[0]  (.A(
        \CoreGPIO_0/CONFIG_reg[0][0] ), .B(
        \CoreGPIO_0/CONFIG_reg[16][0] ), .C(
        \CoreAPB3_0_APBmslave3_PADDR[6] ), .D(
        \CoreAPB3_0_APBmslave3_PADDR[5] ), .Y(
        \CoreGPIO_0/CONFIG_reg_o_2_3_1[0] ));
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_7  (
        .A(\reg_apb_wrp_0/reg16x8_0/mem_8_[0]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_499 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_7_net_1 ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_128  (.A(GND), 
        .B(GND), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[3] ), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[10] ), .IPC());
    CFG4 #( .INIT(16'h8000) )  
        \CoreGPIO_0/xhdl1.GEN_BITS[11].REG_GEN.CONFIG_reg[11]2_0_a4_0_a2  
        (.A(\CoreAPB3_0_APBmslave3_PADDR[3] ), .B(
        \CoreAPB3_0_APBmslave3_PADDR[2] ), .C(\CoreGPIO_0/N_604 ), .D(
        \CoreGPIO_0/N_610 ), .Y(\CoreGPIO_0/CONFIG_reg[11]2 ));
    IP_INTERFACE \FCCC_0/CCC_INST/IP_INTERFACE_10  (.A(VCC), .B(VCC), 
        .C(VCC), .IPA(\FCCC_0/CCC_INST/PLL_ARST_N_net ), .IPB(
        \FCCC_0/CCC_INST/NGMUX2_HOLD_N_net ), .IPC());
    SLE \reg_apb_wrp_0/reg16x8_0/temp_data[0]  (.D(
        \reg_apb_wrp_0/reg16x8_0/N_5_i_0 ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB12_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/rd_enable_net_1 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB2_rgbl_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/temp_data[0]_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_225_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_66_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_225_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_225_rs_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_4_[7]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[7] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB13_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_4__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_170_i ), .ADn(VCC), .SLn(
        VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_4_rs[7] ));
    sdf_IOPAD_TRI \GPIO_OUT_obuf[6]/U0/U_IOPAD  (.PAD(GPIO_OUT[6]), .D(
        \GPIO_OUT_obuf[6]/U0/DOUT ), .E(\GPIO_OUT_obuf[6]/U0/EOUT ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_172  (.A(VCC), 
        .B(VCC), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/MGPIO24B_F2H_GPIN_net ), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/MMUART0_RTS_F2H_SCP_net ), .IPC());
    INV_BA AFLSDF_INV_56 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_61_net_1 ), .Y(
        AFLSDF_INV_56_net_1));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_120_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB11_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_2__1_sqmuxa ), .ALn(
        AFLSDF_INV_22_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(GND)
        , .Q(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_120_set_net_1 ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_202  (.A(VCC), 
        .B(VCC), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[6] ), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[18] ), .IPC());
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_111_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB4_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_13__1_sqmuxa ), .ALn(
        AFLSDF_INV_23_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(GND)
        , .Q(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_111_set_net_1 ));
    IOENFF_BYPASS \GPIO_OUT_obuf[0]/U0/U_IOENFF  (.A(
        \GPIO_OUT_obuf[0]/U0/EOUT1 ), .Y(\GPIO_OUT_obuf[0]/U0/EOUT ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[19].REG_GEN.CONFIG_reg[19][3]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[3] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB9_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[19]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_YR ), .ADn(VCC), .SLn(
        VCC), .SD(GND), .LAT(GND), .Q(\CoreGPIO_0/CONFIG_reg[19][3] ));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_168_rs_RNIJ8NM  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_9_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_168_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_4_rs[6] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_4_[6]_net_1 ));
    CFG4 #( .INIT(16'hAC0F) )  
        \CoreGPIO_0/CONFIG_reg_o_2_31_bm_1_RNO_0[2]  (.A(
        \CoreGPIO_0/CONFIG_reg[9][2] ), .B(
        \CoreGPIO_0/CONFIG_reg[25][2] ), .C(
        \CoreGPIO_0/CONFIG_reg_o_2_18_1[2] ), .D(
        \CoreAPB3_0_APBmslave3_PADDR[5] ), .Y(
        \CoreGPIO_0/CONFIG_reg_o_2_31_bm_1_RNO_0[2]_net_1 ));
    CFG4 #( .INIT(16'h0F35) )  
        \CoreGPIO_0/CONFIG_reg_o_2_31_bm_1_RNO_1[0]  (.A(
        \CoreGPIO_0/CONFIG_reg[5][0] ), .B(
        \CoreGPIO_0/CONFIG_reg[21][0] ), .C(
        \CoreAPB3_0_APBmslave3_PADDR[6] ), .D(
        \CoreAPB3_0_APBmslave3_PADDR[5] ), .Y(
        \CoreGPIO_0/CONFIG_reg_o_2_21_1[0] ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[14].REG_GEN.CONFIG_reg[14][2]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[2] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB14_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[14]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB4_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[14][2] ));
    IP_INTERFACE \FCCC_0/CCC_INST/IP_INTERFACE_0  (.A(VCC), .B(VCC), 
        .C(VCC), .IPA(\FCCC_0/CCC_INST/CLK0_net ), .IPB(
        \FCCC_0/CCC_INST/PSEL_net ), .IPC());
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_222_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_16_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_222_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_222_rs_net_1 ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[3].gpin2[3]  (.D(
        \CoreGPIO_0/gpin1[3] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB9_rgbr_net_1 ), .EN(VCC), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_YR ), .ADn(VCC), .SLn(
        VCC), .SD(GND), .LAT(GND), .Q(\CoreGPIO_0/gpin2[3] ));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_14_[1]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[1] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB6_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_14__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_241_i ), .ADn(VCC), .SLn(
        VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_14_rs[1] ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[4].REG_GEN.CONFIG_reg[4][1]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[1] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB12_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[4]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB2_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0.xhdl1.GEN_BITS[4].REG_GEN.CONFIG_reg[4][1] ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[29].REG_GEN.CONFIG_reg[29][5]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[5] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB13_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[29]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB3_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[29][5] ));
    CFG3 #( .INIT(8'hF2) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_158  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_7_[4]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_498 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_158_i ));
    CFG3 #( .INIT(8'hF2) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_193  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_10_[1]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_491 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_193_i ));
    CFG4 #( .INIT(16'h0001) )  
        \reg_apb_wrp_0/reg16x8_0/temp_data_RNO[2]  (.A(
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_11[2]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_10[2]_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_9[2]_net_1 ), .D(
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_8[2]_net_1 ), .Y(
        \reg_apb_wrp_0/reg16x8_0/N_9_i_0 ));
    sdf_IOPAD_TRI \GPIO_OUT_obuf[2]/U0/U_IOPAD  (.PAD(GPIO_OUT[2]), .D(
        \GPIO_OUT_obuf[2]/U0/DOUT ), .E(\GPIO_OUT_obuf[2]/U0/EOUT ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_190_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_31_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_190_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_190_rs_net_1 ));
    CFG4 #( .INIT(16'hF2F3) )  
        \CoreGPIO_0/xhdl1.GEN_BITS[9].APB_32.INTR_reg_126_0_o2_1_0[9]  
        (.A(\CoreGPIO_0/CONFIG_reg[9][6] ), .B(
        \CoreGPIO_0/edge_neg[9] ), .C(
        \CoreGPIO_0/INTR_reg_126_0_o2_0[9] ), .D(
        \CoreGPIO_0/CONFIG_reg[9][5] ), .Y(
        \CoreGPIO_0/INTR_reg_126_0_o2_1[9] ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_107  (.A(VCC), 
        .B(VCC), .C(VCC), .IPA(), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/FAB_RXVALID_net ), .IPC());
    SLE \reg_apb_wrp_0/reg16x8_0/mem_14_[7]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[7] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB7_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_14__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_247_i ), .ADn(VCC), .SLn(
        VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_14_rs[7] ));
    CFG2 #( .INIT(4'h8) )  
        \reg_apb_wrp_0/reg16x8_0/mem_6__1_sqmuxa_0_a3  (.A(
        \reg_apb_wrp_0/reg16x8_0/N_493 ), .B(
        \reg_apb_wrp_0/wr_enable_net_1 ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_6__1_sqmuxa ));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_8_[2]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[2] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB15_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_8__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_223_i ), .ADn(VCC), .SLn(
        VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_8_rs[2] ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_206_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_127_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_206_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_206_rs_net_1 ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_159  (.A(VCC), 
        .B(VCC), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/SPI0_SS3_F2H_SCP_net ), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/SPI0_SS1_F2H_SCP_net ), .IPC());
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_155  (.A(VCC), 
        .B(VCC), .C(VCC), .IPA(), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/MGPIO8A_F2H_GPIN_net ), .IPC());
    IO_DIFF \FIC_MSS_0/MDDR_DQS_1_PAD/U_ION  (.YIN(GND));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_69  (.A(GND), 
        .B(VCC), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[30] ), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[3] ), .IPC());
    IOTRI_OB_EB \FIC_MSS_0/MDDR_ODT_PAD/U_IOOUT  (.D(VCC), .E(VCC), 
        .DOUT(), .EOUT(\FIC_MSS_0/MDDR_ODT_PAD/EOUT ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[2].gpin2[2]  (.D(
        \CoreGPIO_0/gpin1[2] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB16_rgbr_net_1 ), .EN(VCC), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB6_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(\CoreGPIO_0/gpin2[2] )
        );
    IOBI_IB_OB_EB \FIC_MSS_0/MDDR_DQ_5_PAD/U_IOBI  (.D(VCC), .E(VCC), 
        .YIN(\FIC_MSS_0/MDDR_DQ_5_PAD/YIN ), .DOUT(), .EOUT(), .Y());
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_171_rs_RNIV2EH  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_70_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_171_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_8_rs[6] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_8_[6]_net_1 ));
    CFG4 #( .INIT(16'h7530) )  
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_1[2]  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_15_[2]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/mem_7_[2]_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/N_498 ), .D(
        \reg_apb_wrp_0/reg16x8_0/N_497 ), .Y(
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_1[2]_net_1 ));
    CFG2 #( .INIT(4'h8) )  
        \reg_apb_wrp_0/reg16x8_0/mem_8__1_sqmuxa_0_a3  (.A(
        \reg_apb_wrp_0/reg16x8_0/N_499 ), .B(
        \reg_apb_wrp_0/wr_enable_net_1 ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_8__1_sqmuxa ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_8  (.A(
        \FIC_MSS_0/FIC_MSS_0_FIC_0_APB_MASTER_PRDATA[6] ), .B(
        \FIC_MSS_0_FIC_0_APB_MASTER_PRDATA[13] ), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[6] ), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[13] ), .IPC());
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[0].REG_GEN.CONFIG_reg[0][7]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[7] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB11_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[0]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB1_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[0][7] ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[14].REG_GEN.CONFIG_reg[14][7]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[7] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB13_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[14]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB3_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[14][7] ));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_12_[2]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[2] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB10_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_12__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_226_i ), .ADn(VCC), .SLn(
        VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_12_rs[2] ));
    CFG2 #( .INIT(4'h6) )  \CoreGPIO_0/edge_both_2_sqmuxa_11_i_x2  (.A(
        \CoreGPIO_0/gpin2[4] ), .B(
        \CoreGPIO_0.xhdl1.GEN_BITS[4].gpin3[4] ), .Y(
        \CoreGPIO_0/N_143_i ));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/mem_12__RNI3NVT[6]  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_22_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_230_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_12_rs[6] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_12_[6]_net_1 ));
    CFG4 #( .INIT(16'hFFFE) )  
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_13[1]  (.A(
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_7[1]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_5[1]_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_6[1]_net_1 ), .D(
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_4[1]_net_1 ), .Y(
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_13[1]_net_1 ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[3].REG_GEN.CONFIG_reg[3][6]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[6] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB9_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[3]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_YR ), .ADn(VCC), .SLn(
        VCC), .SD(GND), .LAT(GND), .Q(\CoreGPIO_0/CONFIG_reg[3][6] ));
    CFG4 #( .INIT(16'hAA08) )  
        \CoreGPIO_0/xhdl1.GEN_BITS[1].APB_32.edge_both_23_iv_i_0[1]  (
        .A(\CoreGPIO_0/CONFIG_reg[1][3] ), .B(
        \CoreGPIO_0/edge_both[1] ), .C(
        \CoreAPB3_0_APBmslave3_PWDATA[1] ), .D(\CoreGPIO_0/N_142_i ), 
        .Y(\CoreGPIO_0/N_95 ));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_2_[6]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[6] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB14_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_2__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_150_i ), .ADn(VCC), .SLn(
        VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_2_rs[6] ));
    CFG2 #( .INIT(4'h7) )  \CoreGPIO_0/edge_both_2_sqmuxa_1_i  (.A(
        \CoreGPIO_0/N_248 ), .B(\CoreGPIO_0/CONFIG_reg[17][3] ), .Y(
        \CoreGPIO_0/edge_pos_2_sqmuxa_30_i_1 ));
    CFG3 #( .INIT(8'hF2) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_191  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_10_[0]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_491 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_191_i ));
    CFG4 #( .INIT(16'h1000) )  
        \CoreGPIO_0/xhdl1.GEN_BITS[20].REG_GEN.CONFIG_reg[20]2_0_a4_0_a2  
        (.A(\CoreAPB3_0_APBmslave3_PADDR[3] ), .B(
        \CoreAPB3_0_APBmslave3_PADDR[2] ), .C(\CoreGPIO_0/N_598 ), .D(
        \CoreGPIO_0/N_603 ), .Y(\CoreGPIO_0/CONFIG_reg[20]2 ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_124  (.A(VCC), 
        .B(GND), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/FAB_IDDIG_net ), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[6] ), .IPC());
    IOTRI_OB_EB \FIC_MSS_0/MDDR_BA_2_PAD/U_IOOUT  (.D(VCC), .E(VCC), 
        .DOUT(), .EOUT(\FIC_MSS_0/MDDR_BA_2_PAD/EOUT ));
    CFG3 #( .INIT(8'hB8) )  
        \CoreGPIO_0/xhdl1.GEN_BITS[0].APB_32.INTR_reg_9_0_m2_0[0]  (.A(
        \CoreGPIO_0/edge_neg[0] ), .B(\CoreGPIO_0/CONFIG_reg[0][5] ), 
        .C(\CoreGPIO_0/edge_pos[0] ), .Y(\CoreGPIO_0/N_175 ));
    RGB \FCCC_0/GL1_INST/U0_RGB1_RGB9  (.An(
        \FCCC_0/GL1_INST/U0_YNn_GSouth ), .ENn(GND), .YL(
        \FCCC_0/GL1_INST/U0_RGB1_RGB9_rgbl_net_1 ), .YR(
        \FCCC_0/GL1_INST/U0_RGB1_RGB9_rgbr_net_1 ));
    CFG2 #( .INIT(4'h2) )  
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_a3_11[3]  (.A(
        \reg_apb_wrp_0/reg16x8_0/N_492 ), .B(
        \reg_apb_wrp_0/reg16x8_0/mem_9_[3]_net_1 ), .Y(
        \reg_apb_wrp_0/reg16x8_0/N_414 ));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/mem_11__RNIHEPQ[6]  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_94_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_218_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_11_rs[6] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_11_[6]_net_1 ));
    CFG4 #( .INIT(16'h2000) )  
        \CoreGPIO_0/xhdl1.GEN_BITS[26].REG_GEN.CONFIG_reg[26]2_0_a4_0_a2  
        (.A(\CoreAPB3_0_APBmslave3_PADDR[3] ), .B(
        \CoreAPB3_0_APBmslave3_PADDR[2] ), .C(\CoreGPIO_0/N_598 ), .D(
        \CoreGPIO_0/N_610 ), .Y(\CoreGPIO_0/CONFIG_reg[26]2 ));
    CFG3 #( .INIT(8'hF2) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_250  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_15_[2]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_497 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_250_i ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_15  (.A(
        \FIC_MSS_0_FIC_0_APB_MASTER_PRDATA[20] ), .B(
        \FIC_MSS_0_FIC_0_APB_MASTER_PRDATA[27] ), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[20] ), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[27] ), .IPC());
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_39  (
        .A(\reg_apb_wrp_0/reg16x8_0/mem_6_[5]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_493 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_39_net_1 ));
    IOINFF_BYPASS \FIC_MSS_0/MMUART_0_RXD_PAD/U_IOINFF  (.A(
        \FIC_MSS_0/MMUART_0_RXD_PAD_Y ), .Y(
        \FIC_MSS_0/MMUART_0_RXD_PAD/YIN ));
    CFG3 #( .INIT(8'h20) )  
        \CoreGPIO_0/xhdl1.GEN_BITS[10].APB_32.edge_both_RNO[10]  (.A(
        \CoreGPIO_0/CONFIG_reg[10][3] ), .B(
        \CoreAPB3_0_APBmslave3_PWDATA[10] ), .C(
        \CoreGPIO_0/edge_pos[10] ), .Y(\CoreGPIO_0/edge_neg_149[10] ));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_9_[1]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[1] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB14_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_9__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_177_i ), .ADn(VCC), .SLn(
        VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_9_rs[1] ));
    CFG2 #( .INIT(4'h2) )  \CoreGPIO_0/edge_pos_2_sqmuxa_18_i_a2  (.A(
        \CoreGPIO_0/gpin2[3] ), .B(
        \CoreGPIO_0.xhdl1.GEN_BITS[3].gpin3[3] ), .Y(
        \CoreGPIO_0/N_687 ));
    INV_BA AFLSDF_INV_123 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_118_net_1 ), .Y(
        AFLSDF_INV_123_net_1));
    CFG3 #( .INIT(8'hF2) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_178  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_5_[3]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_490 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_178_i ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_130  (.A(VCC), 
        .B(GND), .C(VCC), .IPA(), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[12] ), .IPC());
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_204_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_125_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_204_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_204_rs_net_1 ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_236  (.A(VCC), 
        .B(VCC), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[34] ), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[46] ), .IPC());
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_79_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB16_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_9__1_sqmuxa ), .ALn(
        AFLSDF_INV_24_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(GND)
        , .Q(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_79_set_net_1 ));
    IOBI_IB_OB_EB \FIC_MSS_0/MDDR_DM_RDQS_0_PAD/U_IOBI  (.D(VCC), .E(
        VCC), .YIN(\FIC_MSS_0/MDDR_DM_RDQS_0_PAD/YIN ), .DOUT(), .EOUT(
        ), .Y());
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[31].REG_GEN.CONFIG_reg[31][1]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[1] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB11_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[31]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB1_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[31][1] ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_187_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_78_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_187_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_187_rs_net_1 ));
    CFG3 #( .INIT(8'hF2) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_252  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_15_[7]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_497 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_252_i ));
    sdf_IOPAD_TRI \GPIO_OUT_obuf[0]/U0/U_IOPAD  (.PAD(GPIO_OUT[0]), .D(
        \GPIO_OUT_obuf[0]/U0/DOUT ), .E(\GPIO_OUT_obuf[0]/U0/EOUT ));
    CFG4 #( .INIT(16'h8000) )  
        \CoreGPIO_0/xhdl1.GEN_BITS[7].REG_GEN.CONFIG_reg[7]2_0_a4_0_a2  
        (.A(\CoreAPB3_0_APBmslave3_PADDR[2] ), .B(
        \CoreAPB3_0_APBmslave3_PADDR[3] ), .C(\CoreGPIO_0/N_603 ), .D(
        \CoreGPIO_0/N_604 ), .Y(\CoreGPIO_0/CONFIG_reg[7]2 ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_109_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB4_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_13__1_sqmuxa ), .ALn(
        AFLSDF_INV_25_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(GND)
        , .Q(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_109_set_net_1 ));
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_126  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_3_[2]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_494 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_126_net_1 ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[0].APB_32.edge_both[0]  (.D(
        \CoreGPIO_0/N_97 ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB10_rgbr_net_1 ), .EN(
        \CoreGPIO_0/N_80 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB0_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/edge_both[0] ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_223  (.A(VCC), 
        .B(VCC), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[7] ), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[19] ), .IPC());
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_236_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_108_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_236_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_236_rs_net_1 ));
    RGB \FCCC_0/GL1_INST/U0_RGB1_RGB18  (.An(
        \FCCC_0/GL1_INST/U0_YNn_GSouth ), .ENn(GND), .YL(
        \FCCC_0/GL1_INST/U0_RGB1_RGB18_rgbl_net_1 ), .YR());
    CFG4 #( .INIT(16'h4657) )  
        \CoreGPIO_0/CONFIG_reg_o_2_31_am_1_1[1]  (.A(
        \CoreAPB3_0_APBmslave3_PADDR[4] ), .B(
        \CoreAPB3_0_APBmslave3_PADDR[3] ), .C(
        \CoreGPIO_0/CONFIG_reg_o_2_31_am_1_1_RNO[1]_net_1 ), .D(
        \CoreGPIO_0/CONFIG_reg_o_2_31_am_1_RNO_0[1]_net_1 ), .Y(
        \CoreGPIO_0/CONFIG_reg_o_2_31_am_1[1] ));
    CFG4 #( .INIT(16'hEAFA) )  \FIC_MSS_0/MSS_ADLIB_INST_RNO_4  (.A(
        \FIC_MSS_0/CoreAPB3_0_APBmslave5_PRDATA_m_0_0[5] ), .B(
        \CoreGPIO_0.PRDATA_iv_0_0_1[5] ), .C(
        CoreAPB3_0_APBmslave5_PSELx), .D(
        \FIC_MSS_0/CoreAPB3_0_APBmslave5_PRDATA_m_0_1_1[5] ), .Y(
        \FIC_MSS_0/FIC_MSS_0_FIC_0_APB_MASTER_PRDATA[5] ));
    CFG2 #( .INIT(4'h4) )  \CoreGPIO_0/PRDATA_0_iv_0_a2_0[24]  (.A(
        \CoreGPIO_0.N_247 ), .B(\CoreGPIO_0/INTR_reg[24] ), .Y(
        \CoreGPIO_0.N_538 ));
    CFG3 #( .INIT(8'hF2) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_153  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_3_[1]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_494 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_153_i ));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_6_[0]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[0] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB13_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_6__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_188_i ), .ADn(VCC), .SLn(
        VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_6_rs[0] ));
    IOTRI_OB_EB \FIC_MSS_0/MDDR_CKE_PAD/U_IOOUT  (.D(VCC), .E(VCC), 
        .DOUT(), .EOUT(\FIC_MSS_0/MDDR_CKE_PAD/EOUT ));
    CFG3 #( .INIT(8'h80) )  
        \CoreGPIO_0/xhdl1.GEN_BITS[0].APB_32.INTR_reg21_0_a2  (.A(
        CoreAPB3_0_APBmslave3_PENABLE), .B(CoreAPB3_0_APBmslave5_PSELx)
        , .C(CoreAPB3_0_APBmslave3_PWRITE), .Y(\CoreGPIO_0/INTR_reg21 )
        );
    IOTRI_OB_EB \FIC_MSS_0/MDDR_ADDR_11_PAD/U_IOOUT  (.D(VCC), .E(VCC), 
        .DOUT(), .EOUT(\FIC_MSS_0/MDDR_ADDR_11_PAD/EOUT ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_248_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_57_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_248_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_248_rs_net_1 ));
    CFG4 #( .INIT(16'h0F35) )  
        \CoreGPIO_0/CONFIG_reg_o_2_31_bm_1_RNO_2[2]  (.A(
        \CoreGPIO_0/CONFIG_reg[1][2] ), .B(
        \CoreGPIO_0/CONFIG_reg[17][2] ), .C(
        \CoreAPB3_0_APBmslave3_PADDR[6] ), .D(
        \CoreAPB3_0_APBmslave3_PADDR[5] ), .Y(
        \CoreGPIO_0/CONFIG_reg_o_2_18_1[2] ));
    CFG4 #( .INIT(16'h0001) )  
        \reg_apb_wrp_0/reg16x8_0/WRITE_GEN.mem_0__2_i_0_0_a2[5]  (.A(
        \CoreAPB3_0_APBmslave3_PADDR[3] ), .B(
        \CoreAPB3_0_APBmslave3_PADDR[2] ), .C(
        \CoreAPB3_0_APBmslave3_PADDR[0] ), .D(
        \CoreAPB3_0_APBmslave3_PADDR[1] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/N_496 ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_178_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_42_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_178_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_178_rs_net_1 ));
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_16  (
        .A(\reg_apb_wrp_0/reg16x8_0/mem_12_[0]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_495 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_16_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_0_[5]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[5] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB19_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_0__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_133_i ), .ADn(VCC), .SLn(
        VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_0_rs[5] ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[16].REG_GEN.CONFIG_reg[16][7]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[7] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB11_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[16]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB1_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[16][7] ));
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_68  (
        .A(\reg_apb_wrp_0/reg16x8_0/mem_8_[4]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_499 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_68_net_1 ));
    INV_BA AFLSDF_INV_34 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_47_net_1 ), .Y(
        AFLSDF_INV_34_net_1));
    CFG3 #( .INIT(8'hF2) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_249  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_15_[1]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_497 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_249_i ));
    CFG4 #( .INIT(16'hEFEE) )  
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_11[0]  (.A(
        \reg_apb_wrp_0/reg16x8_0/N_368 ), .B(
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_7[0]_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_0_[0]_net_1 ), .D(
        \reg_apb_wrp_0/reg16x8_0/N_496 ), .Y(
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_11[0]_net_1 ));
    CFG4 #( .INIT(16'h5410) )  \CoreGPIO_0/PRDATA_iv_0_0_1[5]  (.A(
        \CoreAPB3_0_APBmslave3_PADDR[7] ), .B(
        \CoreAPB3_0_APBmslave3_PADDR[2] ), .C(
        \CoreGPIO_0/CONFIG_reg_o_2_31_am[5]_net_1 ), .D(
        \CoreGPIO_0/CONFIG_reg_o_2_31_bm[5]_net_1 ), .Y(
        \CoreGPIO_0.PRDATA_iv_0_0_1[5] ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_49_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB6_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_7__1_sqmuxa ), .ALn(
        AFLSDF_INV_26_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(GND)
        , .Q(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_49_set_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_14_[6]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[6] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB13_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_14__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_246_i ), .ADn(VCC), .SLn(
        VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_14_rs[6] ));
    CFG4 #( .INIT(16'h7350) )  
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_6[3]  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_8_[3]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/mem_0_[3]_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/N_499 ), .D(
        \reg_apb_wrp_0/reg16x8_0/N_496 ), .Y(
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_6[3]_net_1 ));
    CFG4 #( .INIT(16'hB383) )  \CoreGPIO_0/CONFIG_reg_o_2_31_bm[2]  (
        .A(\CoreGPIO_0/CONFIG_reg_o_2_31_bm_RNO[2]_net_1 ), .B(
        \CoreGPIO_0/CONFIG_reg_o_2_31_bm_1[2] ), .C(
        \CoreAPB3_0_APBmslave3_PADDR[3] ), .D(
        \CoreGPIO_0/CONFIG_reg_o_2_31_bm_RNO_0[2]_net_1 ), .Y(
        \CoreGPIO_0/CONFIG_reg_o_2_31_bm[2]_net_1 ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_285  (.A(VCC), 
        .B(VCC), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PADDR_net[8] ), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[12] ), .IPC());
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_28  (
        .A(\reg_apb_wrp_0/reg16x8_0/mem_2_[1]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_501 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_28_net_1 ));
    CFG4 #( .INIT(16'hBBFB) )  \CoreGPIO_0/edge_neg_2_sqmuxa_25_i_0  (
        .A(\CoreGPIO_0/N_401 ), .B(\CoreGPIO_0/CONFIG_reg[0][3] ), .C(
        \CoreGPIO_0/INTR_reg21 ), .D(\CoreGPIO_0.N_247 ), .Y(
        \CoreGPIO_0/N_52 ));
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_44  (
        .A(\reg_apb_wrp_0/reg16x8_0/mem_5_[4]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_490 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_44_net_1 ));
    IOIN_IB \FIC_MSS_0/MDDR_DQS_TMATCH_0_IN_PAD/U_IOIN  (.YIN(
        \FIC_MSS_0/MDDR_DQS_TMATCH_0_IN_PAD/YIN ), .E(GND), .Y());
    CFG2 #( .INIT(4'h4) )  \CoreGPIO_0/PRDATA_0_iv_0_a2_0[20]  (.A(
        \CoreGPIO_0.N_247 ), .B(\CoreGPIO_0/INTR_reg[20] ), .Y(
        \CoreGPIO_0.N_546 ));
    CFG3 #( .INIT(8'hF2) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_151  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_2_[7]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_501 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_151_i ));
    CFG4 #( .INIT(16'h7350) )  
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_6[7]  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_8_[7]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/mem_0_[7]_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/N_499 ), .D(
        \reg_apb_wrp_0/reg16x8_0/N_496 ), .Y(
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_6[7]_net_1 ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[26].APB_32.INTR_reg[26]  (.D(
        \CoreGPIO_0/INTR_reg_347[26] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB16_rgbr_net_1 ), .EN(VCC), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB6_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0.xhdl1.GEN_BITS[26].APB_32.INTR_reg[26] ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_234_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_106_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_234_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_234_rs_net_1 ));
    CFG4 #( .INIT(16'hEFEE) )  
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_10[2]  (.A(
        \reg_apb_wrp_0/reg16x8_0/N_392 ), .B(
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_5[2]_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_4_[2]_net_1 ), .D(
        \reg_apb_wrp_0/reg16x8_0/N_504 ), .Y(
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_10[2]_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_228_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_20_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_228_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_228_rs_net_1 ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[24].APB_32.GPOUT_reg[24]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[24] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB9_rgbr_net_1 ), .EN(
        \CoreGPIO_0/GPOUT_reg_0_sqmuxa ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_YR ), .ADn(VCC), .SLn(
        VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0.xhdl1.GEN_BITS[24].APB_32.GPOUT_reg[24] ));
    RGB \FCCC_0/GL1_INST/U0_RGB1_RGB16  (.An(
        \FCCC_0/GL1_INST/U0_YNn_GSouth ), .ENn(GND), .YL(
        \FCCC_0/GL1_INST/U0_RGB1_RGB16_rgbl_net_1 ), .YR(
        \FCCC_0/GL1_INST/U0_RGB1_RGB16_rgbr_net_1 ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[11].APB_32.INTR_reg[11]  (.D(
        \CoreGPIO_0/INTR_reg_152[11] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB13_rgbr_net_1 ), .EN(VCC), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB3_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/INTR_reg[11] ));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_7_[4]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[4] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB8_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_7__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_158_i ), .ADn(VCC), .SLn(
        VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_7_rs[4] ));
    CFG4 #( .INIT(16'hBBFB) )  \CoreGPIO_0/edge_neg_2_sqmuxa_8_i_0  (
        .A(\CoreGPIO_0/N_397 ), .B(\CoreGPIO_0/CONFIG_reg[4][3] ), .C(
        \CoreGPIO_0/INTR_reg21 ), .D(\CoreGPIO_0.N_247 ), .Y(
        \CoreGPIO_0/N_58 ));
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_35  (
        .A(\reg_apb_wrp_0/reg16x8_0/mem_6_[3]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_493 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_35_net_1 ));
    INV_BA AFLSDF_INV_19 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_41_net_1 ), .Y(
        AFLSDF_INV_19_net_1));
    CFG4 #( .INIT(16'h0400) )  
        \CoreGPIO_0/xhdl1.GEN_BITS[8].REG_GEN.CONFIG_reg[8]2_0_a4_0_a2  
        (.A(\CoreAPB3_0_APBmslave3_PADDR[7] ), .B(\CoreGPIO_0/N_610 ), 
        .C(\CoreGPIO_0/N_243 ), .D(\CoreGPIO_0/INTR_reg21 ), .Y(
        \CoreGPIO_0/CONFIG_reg[8]2 ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_18_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB10_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_12__1_sqmuxa ), .ALn(
        AFLSDF_INV_27_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(GND)
        , .Q(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_18_set_net_1 ));
    IOTRI_OB_EB \FIC_MSS_0/MDDR_DQS_TMATCH_0_OUT_PAD/U_IOOUT  (.D(VCC), 
        .E(VCC), .DOUT(), .EOUT(
        \FIC_MSS_0/MDDR_DQS_TMATCH_0_OUT_PAD/EOUT ));
    sdf_IOPAD_TRI \FIC_MSS_0/MDDR_ADDR_14_PAD/U_IOPAD  (.PAD(
        MDDR_ADDR[14]), .D(\FIC_MSS_0/DRAM_ADDR_net_0[14] ), .E(
        \FIC_MSS_0/MDDR_ADDR_14_PAD/EOUT ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[15].APB_32.GPOUT_reg[15]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[15] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB9_rgbr_net_1 ), .EN(
        \CoreGPIO_0/GPOUT_reg_0_sqmuxa ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_YR ), .ADn(VCC), .SLn(
        VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0.xhdl1.GEN_BITS[15].APB_32.GPOUT_reg[15] ));
    CFG4 #( .INIT(16'hFF4F) )  \CoreGPIO_0/edge_both_2_sqmuxa_14_i_0  
        (.A(\CoreGPIO_0.N_247 ), .B(\CoreGPIO_0/INTR_reg21 ), .C(
        \CoreGPIO_0/CONFIG_reg[1][3] ), .D(\CoreGPIO_0/N_142_i ), .Y(
        \CoreGPIO_0/N_82 ));
    CFG3 #( .INIT(8'hF2) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_173  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_8_[7]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_499 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_173_i ));
    CFG4 #( .INIT(16'hFFFE) )  
        \CoreGPIO_0/xhdl1.GEN_BITS[0].APB_32.un5_PRDATA_o_0_a2_0_o2_sx  
        (.A(\CoreAPB3_0_APBmslave3_PADDR[2] ), .B(
        \CoreAPB3_0_APBmslave3_PADDR[4] ), .C(
        \CoreAPB3_0_APBmslave3_PADDR[5] ), .D(
        \CoreAPB3_0_APBmslave3_PADDR[3] ), .Y(
        \CoreGPIO_0/un5_PRDATA_o_0_a2_0_o2_sx ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_182  (.A(VCC), 
        .B(VCC), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/MGPIO27B_F2H_GPIN_net ), .IPB(), 
        .IPC());
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_170_rs_RNIMMRL  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_11_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_170_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_4_rs[7] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_4_[7]_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_95_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB16_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_11__1_sqmuxa ), .ALn(
        AFLSDF_INV_28_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(GND)
        , .Q(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_95_set_net_1 ));
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_6  (
        .A(\reg_apb_wrp_0/reg16x8_0/mem_4_[3]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_504 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_6_net_1 ));
    CFG2 #( .INIT(4'h2) )  
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_a3_5[0]  (.A(
        \reg_apb_wrp_0/reg16x8_0/N_495 ), .B(
        \reg_apb_wrp_0/reg16x8_0/mem_12_[0]_net_1 ), .Y(
        \reg_apb_wrp_0/reg16x8_0/N_360 ));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_31_set_RNIMA8B  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_31_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_190_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_6_rs[1] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_6_[1]_net_1 ));
    INV_BA AFLSDF_INV_17 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_71_net_1 ), .Y(
        AFLSDF_INV_17_net_1));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_146  (.A(VCC), 
        .B(VCC), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/MGPIO0A_F2H_GPIN_net ), .IPB(), .IPC(
        ));
    SLE \reg_apb_wrp_0/reg16x8_0/temp_data[4]  (.D(
        \reg_apb_wrp_0/reg16x8_0/N_19_i_0 ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB11_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/rd_enable_net_1 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB1_rgbl_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/temp_data[4]_net_1 ));
    CFG4 #( .INIT(16'h0800) )  
        \reg_apb_wrp_0/reg16x8_0/WRITE_GEN.mem_14__2_i_a2[4]  (.A(
        \CoreAPB3_0_APBmslave3_PADDR[3] ), .B(
        \CoreAPB3_0_APBmslave3_PADDR[2] ), .C(
        \CoreAPB3_0_APBmslave3_PADDR[0] ), .D(
        \CoreAPB3_0_APBmslave3_PADDR[1] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/N_503 ));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_133_rs_RNIRKPK  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_86_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_133_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_0_rs[5] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_0_[5]_net_1 ));
    CFG0 #( .INIT(1'h0) )  CFG0_GND_INST (.Y(CFG0_GND_INST_NET));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_167_rs_RNI9A1R  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_68_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_167_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_8_rs[4] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_8_[4]_net_1 ));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_35_set_RNI09DG  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_35_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_194_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_6_rs[3] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_6_[3]_net_1 ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_74  (.A(VCC), 
        .B(VCC), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[8] ), .IPB(), 
        .IPC());
    CFG2 #( .INIT(4'h8) )  
        \CoreGPIO_0/xhdl1.GEN_BITS[6].REG_GPOUT.un64_GPIO_OUT_i  (.A(
        \CoreGPIO_0.xhdl1.GEN_BITS[6].APB_32.GPOUT_reg[6] ), .B(
        \CoreGPIO_0/CONFIG_reg[6][0] ), .Y(\GPIO_OUT_net_2[6] ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[9].REG_GEN.CONFIG_reg[9][2]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[2] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB16_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[9]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB6_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[9][2] ));
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_2  (
        .A(\reg_apb_wrp_0/reg16x8_0/mem_4_[1]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_504 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_2_net_1 ));
    CFG4 #( .INIT(16'hAC0F) )  
        \CoreGPIO_0/CONFIG_reg_o_2_31_bm_1_1_RNO[5]  (.A(
        \CoreGPIO_0/CONFIG_reg[13][5] ), .B(
        \CoreGPIO_0/CONFIG_reg[29][5] ), .C(
        \CoreGPIO_0/CONFIG_reg_o_2_21_1[5] ), .D(
        \CoreAPB3_0_APBmslave3_PADDR[5] ), .Y(
        \CoreGPIO_0/CONFIG_reg_o_2_31_bm_1_1_RNO[5]_net_1 ));
    CFG4 #( .INIT(16'h330A) )  
        \CoreGPIO_0/xhdl1.GEN_BITS[28].APB_32.INTR_reg_373_0[28]  (.A(
        \CoreGPIO_0/INTR_reg[28] ), .B(
        \CoreGPIO_0/INTR_reg_373_0_o2_1[28] ), .C(
        \CoreAPB3_0_APBmslave3_PWDATA[28] ), .D(\CoreGPIO_0/N_248 ), 
        .Y(\CoreGPIO_0/INTR_reg_373[28] ));
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_11  (
        .A(\reg_apb_wrp_0/reg16x8_0/mem_4_[7]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_504 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_11_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_0_[7]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[7] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB2_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_0__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_135_i ), .ADn(VCC), .SLn(
        VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_0_rs[7] ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_59  (.A(VCC), 
        .B(GND), .C(VCC), .IPA(), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[20] ), .IPC());
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_234  (.A(VCC), 
        .B(VCC), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[32] ), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[44] ), .IPC());
    CFG3 #( .INIT(8'hF2) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_171  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_8_[6]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_499 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_171_i ));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/mem_14__RNIGAHT[0]  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_112_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_240_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_14_rs[0] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_14_[0]_net_1 ));
    CFG4 #( .INIT(16'hAC0F) )  
        \CoreGPIO_0/CONFIG_reg_o_2_31_bm_RNO_0[6]  (.A(
        \CoreGPIO_0/CONFIG_reg[15][6] ), .B(
        \CoreGPIO_0/CONFIG_reg[31][6] ), .C(
        \CoreGPIO_0/CONFIG_reg_o_2_28_1_1[6] ), .D(
        \CoreAPB3_0_APBmslave3_PADDR[5] ), .Y(
        \CoreGPIO_0/CONFIG_reg_o_2_31_bm_RNO_0[6]_net_1 ));
    IOBI_IB_OB_EB \FIC_MSS_0/MDDR_DQ_6_PAD/U_IOBI  (.D(VCC), .E(VCC), 
        .YIN(\FIC_MSS_0/MDDR_DQ_6_PAD/YIN ), .DOUT(), .EOUT(), .Y());
    IOINFF_BYPASS \FIC_MSS_0/MDDR_DQ_13_PAD/U_IOINFF  (.A(
        \FIC_MSS_0/MDDR_DQ_13_PAD_Y ), .Y(
        \FIC_MSS_0/MDDR_DQ_13_PAD/YIN ));
    INV_BA AFLSDF_INV_126 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_81_net_1 ), .Y(
        AFLSDF_INV_126_net_1));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[15].REG_GEN.CONFIG_reg[15][4]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[4] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB10_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[15]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB0_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[15][4] ));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_165_rs_RNI08GR  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_65_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_165_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_4_rs[4] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_4_[4]_net_1 ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_241  (.A(VCC), 
        .B(GND), .C(GND), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[53] ), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/F_WSTRB_net[1] ), .IPC(
        \FIC_MSS_0/MSS_ADLIB_INST/F_BREADY_net ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_49  (.A(GND), 
        .B(VCC), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[3] ), .IPB(), .IPC());
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[9].APB_32.GPOUT_reg[9]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[9] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB14_rgbr_net_1 ), .EN(
        \CoreGPIO_0/GPOUT_reg_0_sqmuxa ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB4_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0.xhdl1.GEN_BITS[9].APB_32.GPOUT_reg[9] ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_116  (.A(GND), 
        .B(VCC), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/FAB_RXVALIDH_net ), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/FAB_VSTATUS_net[5] ), .IPC());
    CFG4 #( .INIT(16'hAC0F) )  
        \CoreGPIO_0/CONFIG_reg_o_2_31_am_1_RNO_0[3]  (.A(
        \CoreGPIO_0/CONFIG_reg[8][3] ), .B(
        \CoreGPIO_0/CONFIG_reg[24][3] ), .C(
        \CoreGPIO_0/CONFIG_reg_o_2_3_1[3] ), .D(
        \CoreAPB3_0_APBmslave3_PADDR[5] ), .Y(
        \CoreGPIO_0/CONFIG_reg_o_2_31_am_1_RNO_0[3]_net_1 ));
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_37  (
        .A(\reg_apb_wrp_0/reg16x8_0/mem_6_[4]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_493 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_37_net_1 ));
    CFG4 #( .INIT(16'hAC0F) )  
        \CoreGPIO_0/CONFIG_reg_o_2_31_am_RNO[2]  (.A(
        \CoreGPIO_0/CONFIG_reg[10][2] ), .B(
        \CoreGPIO_0/CONFIG_reg[26][2] ), .C(
        \CoreGPIO_0/CONFIG_reg_o_2_10_1_1[2] ), .D(
        \CoreAPB3_0_APBmslave3_PADDR[5] ), .Y(
        \CoreGPIO_0/CONFIG_reg_o_2_31_am_RNO[2]_net_1 ));
    sdf_IOPAD_BI \FIC_MSS_0/MDDR_DQ_13_PAD/U_IOPAD  (.PAD(MDDR_DQ[13]), 
        .D(\FIC_MSS_0/DRAM_DQ_OUT_net_0[13] ), .E(
        \FIC_MSS_0/DRAM_DQ_OE_net_0[13] ), .Y(
        \FIC_MSS_0/MDDR_DQ_13_PAD_Y ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_147_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_32_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_147_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_147_rs_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_2_[3]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[3] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB8_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_2__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_147_i ), .ADn(VCC), .SLn(
        VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_2_rs[3] ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_143  (.A(VCC), 
        .B(VCC), .C(VCC), .IPA(), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/FAB_M3_RESET_N_net ), .IPC());
    CFG4 #( .INIT(16'hAC0F) )  
        \CoreGPIO_0/CONFIG_reg_o_2_31_am_RNO[3]  (.A(
        \CoreGPIO_0/CONFIG_reg[10][3] ), .B(
        \CoreGPIO_0/CONFIG_reg[26][3] ), .C(
        \CoreGPIO_0/CONFIG_reg_o_2_10_1_1[3] ), .D(
        \CoreAPB3_0_APBmslave3_PADDR[5] ), .Y(
        \CoreGPIO_0/CONFIG_reg_o_2_31_am_RNO[3]_net_1 ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_71  (.A(VCC), 
        .B(VCC), .C(VCC), .IPA(), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[5] ), .IPC());
    CFG3 #( .INIT(8'hF2) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_229  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_12_[5]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_495 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_229_i ));
    CFG4 #( .INIT(16'h2000) )  
        \CoreGPIO_0/xhdl1.GEN_BITS[14].REG_GEN.CONFIG_reg[14]2_0_a4_0_a2  
        (.A(\CoreAPB3_0_APBmslave3_PADDR[3] ), .B(
        \CoreAPB3_0_APBmslave3_PADDR[2] ), .C(\CoreGPIO_0/N_604 ), .D(
        \CoreGPIO_0/N_605 ), .Y(\CoreGPIO_0/CONFIG_reg[14]2 ));
    CFG4 #( .INIT(16'hF2F3) )  
        \CoreGPIO_0/xhdl1.GEN_BITS[22].APB_32.INTR_reg_295_0_o2_1_0[22]  
        (.A(\CoreGPIO_0/CONFIG_reg[22][6] ), .B(
        \CoreGPIO_0/edge_neg[22] ), .C(
        \CoreGPIO_0/INTR_reg_295_0_o2_0[22] ), .D(
        \CoreGPIO_0/CONFIG_reg[22][5] ), .Y(
        \CoreGPIO_0/INTR_reg_295_0_o2_1[22] ));
    CFG3 #( .INIT(8'hF2) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_167  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_8_[4]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_499 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_167_i ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[25].APB_32.GPOUT_reg[25]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[25] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB14_rgbr_net_1 ), .EN(
        \CoreGPIO_0/GPOUT_reg_0_sqmuxa ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB4_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0.xhdl1.GEN_BITS[25].APB_32.GPOUT_reg[25] ));
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_42  (
        .A(\reg_apb_wrp_0/reg16x8_0/mem_5_[3]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_490 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_42_net_1 ));
    IOTRI_OB_EB \GPIO_OUT_obuf[0]/U0/U_IOTRI  (.D(\GPIO_OUT_net_2[0] ), 
        .E(VCC), .DOUT(\GPIO_OUT_obuf[0]/U0/DOUT1 ), .EOUT(
        \GPIO_OUT_obuf[0]/U0/EOUT1 ));
    CFG3 #( .INIT(8'h20) )  
        \CoreGPIO_0/xhdl1.GEN_BITS[20].APB_32.edge_both_RNO[20]  (.A(
        \CoreGPIO_0/CONFIG_reg[20][3] ), .B(
        \CoreAPB3_0_APBmslave3_PWDATA[20] ), .C(
        \CoreGPIO_0/edge_neg[20] ), .Y(\CoreGPIO_0/edge_neg_289[20] ));
    IOTRI_OB_EB \FIC_MSS_0/MDDR_ADDR_6_PAD/U_IOOUT  (.D(VCC), .E(VCC), 
        .DOUT(), .EOUT(\FIC_MSS_0/MDDR_ADDR_6_PAD/EOUT ));
    CFG3 #( .INIT(8'hF2) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_234  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_13_[2]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_500 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_234_i ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_3  (.A(
        \FIC_MSS_0/FIC_MSS_0_FIC_0_APB_MASTER_PRDATA[1] ), .B(
        \FIC_MSS_0_FIC_0_APB_MASTER_PRDATA[8] ), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[1] ), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[8] ), .IPC());
    CFG4 #( .INIT(16'hEFEE) )  
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_8[1]  (.A(
        \reg_apb_wrp_0/reg16x8_0/N_374 ), .B(
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_1[1]_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_5_[1]_net_1 ), .D(
        \reg_apb_wrp_0/reg16x8_0/N_490 ), .Y(
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_8[1]_net_1 ));
    CFG3 #( .INIT(8'h7F) )  \FIC_MSS_0/MSS_ADLIB_INST_RNO_18  (.A(
        \CoreGPIO_0.xhdl1.GEN_BITS[4].gpin3[4] ), .B(
        \CoreGPIO_0.RDATA_32.un12_PRDATA_o ), .C(
        \CoreGPIO_0.xhdl1.GEN_BITS[4].REG_GEN.CONFIG_reg[4][1] ), .Y(
        \FIC_MSS_0/CoreAPB3_0_APBmslave5_PRDATA_m_0_1_0[4] ));
    CFG2 #( .INIT(4'h4) )  \CoreGPIO_0/PRDATA_0_iv_0_a2_0[8]  (.A(
        \CoreGPIO_0.N_247 ), .B(\CoreGPIO_0/INTR_reg[8] ), .Y(
        \CoreGPIO_0.N_570 ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_188_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_29_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_188_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_188_rs_net_1 ));
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_73  (
        .A(\reg_apb_wrp_0/reg16x8_0/mem_9_[1]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_492 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_73_net_1 ));
    INV_BA AFLSDF_INV_72 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_57_net_1 ), .Y(
        AFLSDF_INV_72_net_1));
    CFG2 #( .INIT(4'h7) )  \CoreGPIO_0/edge_both_2_sqmuxa_3_i  (.A(
        \CoreGPIO_0/N_248 ), .B(\CoreGPIO_0/CONFIG_reg[16][3] ), .Y(
        \CoreGPIO_0/edge_pos_2_sqmuxa_29_i_1 ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_211  (.A(VCC), 
        .B(GND), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[29] ), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/F_AWLOCK_HMASTLOCK0_net[1] ), .IPC());
    IP_INTERFACE \FCCC_0/CCC_INST/IP_INTERFACE_13  (.A(VCC), .B(VCC), 
        .C(VCC), .IPA(\FCCC_0/CCC_INST/NGMUX1_ARST_N_net ), .IPB(), 
        .IPC(\FCCC_0/CCC_INST/PADDR_net[3] ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[6].APB_32.edge_neg[6]  (.D(
        \CoreGPIO_0/N_113 ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB12_rgbr_net_1 ), .EN(
        \CoreGPIO_0/N_62 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB2_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/edge_neg[6] ));
    CFG4 #( .INIT(16'h0CAE) )  \CoreGPIO_0/PRDATA_iv_0_0_1[2]  (.A(
        \CoreGPIO_0/PRDATA_iv_0_0_a2_0_0[2]_net_1 ), .B(
        \CoreGPIO_0/INTR_reg[2] ), .C(\CoreGPIO_0.N_247 ), .D(
        \CoreGPIO_0.N_246 ), .Y(\CoreGPIO_0.PRDATA_iv_0_0_1[2] ));
    CFG3 #( .INIT(8'hF2) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_134  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_0_[6]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_496 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_134_i ));
    CFG4 #( .INIT(16'hF2F3) )  
        \CoreGPIO_0/xhdl1.GEN_BITS[7].APB_32.INTR_reg_100_0_o2_1_0[7]  
        (.A(\CoreGPIO_0/CONFIG_reg[7][6] ), .B(
        \CoreGPIO_0/edge_pos[7] ), .C(
        \CoreGPIO_0/INTR_reg_100_0_o2_0[7] ), .D(
        \CoreGPIO_0/CONFIG_reg[7][5] ), .Y(
        \CoreGPIO_0/INTR_reg_100_0_o2_1[7] ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_113  (.A(VCC), 
        .B(VCC), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/FAB_XDATAIN_net[5] ), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/FAB_VSTATUS_net[2] ), .IPC());
    CFG4 #( .INIT(16'h7350) )  
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_3[6]  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_11_[6]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/mem_3_[6]_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/N_505 ), .D(
        \reg_apb_wrp_0/reg16x8_0/N_494 ), .Y(
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_3[6]_net_1 ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[12].APB_32.INTR_reg[12]  (.D(
        \CoreGPIO_0/INTR_reg_165[12] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB13_rgbr_net_1 ), .EN(VCC), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB3_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/INTR_reg[12] ));
    CFG4 #( .INIT(16'h4657) )  
        \CoreGPIO_0/CONFIG_reg_o_2_31_bm_1_1[1]  (.A(
        \CoreAPB3_0_APBmslave3_PADDR[4] ), .B(
        \CoreAPB3_0_APBmslave3_PADDR[3] ), .C(
        \CoreGPIO_0/CONFIG_reg_o_2_31_bm_1_1_RNO[1]_net_1 ), .D(
        \CoreGPIO_0/CONFIG_reg_o_2_31_bm_1_RNO_0[1]_net_1 ), .Y(
        \CoreGPIO_0/CONFIG_reg_o_2_31_bm_1[1] ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[30].APB_32.edge_both[30]  (.D(
        \CoreGPIO_0/edge_neg_429[30] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB13_rgbr_net_1 ), .EN(
        \CoreGPIO_0/edge_neg_2_sqmuxa_6_i_1 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB3_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/edge_pos[30] ));
    CFG3 #( .INIT(8'h7F) )  \FIC_MSS_0/MSS_ADLIB_INST_RNO_28  (.A(
        \CoreGPIO_0.xhdl1.GEN_BITS[1].gpin3[1] ), .B(
        \CoreGPIO_0.RDATA_32.un12_PRDATA_o ), .C(
        \CoreGPIO_0.xhdl1.GEN_BITS[1].REG_GEN.CONFIG_reg[1][1] ), .Y(
        \FIC_MSS_0/CoreAPB3_0_APBmslave5_PRDATA_m_0_1_0[1] ));
    CFG2 #( .INIT(4'h1) )  
        \CoreGPIO_0/xhdl1.GEN_BITS[0].REG_GEN.CONFIG_reg[0]2_0_a4_0_a2_0  
        (.A(\CoreAPB3_0_APBmslave3_PADDR[5] ), .B(
        \CoreAPB3_0_APBmslave3_PADDR[4] ), .Y(\CoreGPIO_0/N_606 ));
    CFG4 #( .INIT(16'h0F35) )  
        \CoreGPIO_0/CONFIG_reg_o_2_31_bm_1_RNO_2[4]  (.A(
        \CoreGPIO_0/CONFIG_reg[1][4] ), .B(
        \CoreGPIO_0/CONFIG_reg[17][4] ), .C(
        \CoreAPB3_0_APBmslave3_PADDR[6] ), .D(
        \CoreAPB3_0_APBmslave3_PADDR[5] ), .Y(
        \CoreGPIO_0/CONFIG_reg_o_2_18_1[4] ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[22].REG_GEN.CONFIG_reg[22][5]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[5] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB12_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[22]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB2_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[22][5] ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_217_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_1_net_1 ), .EN(VCC), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_217_i ), .ADn(VCC), .SLn(
        VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_217_rs_net_1 ));
    CFG4 #( .INIT(16'hC5CA) )  
        \CoreGPIO_0/xhdl1.GEN_BITS[2].APB_32.INTR_reg_35_0_m2[2]  (.A(
        \CoreGPIO_0.xhdl1.GEN_BITS[2].gpin3[2] ), .B(
        \CoreGPIO_0/N_173 ), .C(\CoreGPIO_0/CONFIG_reg[2][6] ), .D(
        \CoreGPIO_0/CONFIG_reg[2][5] ), .Y(\CoreGPIO_0/N_178 ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_100  (.A(VCC), 
        .B(VCC), .C(VCC), .IPA(\FIC_MSS_0/MSS_ADLIB_INST/RCGF_net[0] ), 
        .IPB(\FIC_MSS_0/MSS_ADLIB_INST/RCGF_net[7] ), .IPC());
    CFG2 #( .INIT(4'h8) )  
        \reg_apb_wrp_0/reg16x8_0/mem_13__1_sqmuxa_0_a2_0_a3  (.A(
        \reg_apb_wrp_0/reg16x8_0/N_500 ), .B(
        \reg_apb_wrp_0/wr_enable_net_1 ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_13__1_sqmuxa ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_206  (.A(VCC), 
        .B(GND), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[24] ), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/F_AWLEN_HBURST0_net[2] ), .IPC());
    INV_BA AFLSDF_INV_124 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_58_net_1 ), .Y(
        AFLSDF_INV_124_net_1));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_220  (.A(VCC), 
        .B(VCC), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[4] ), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[16] ), .IPC());
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[18].APB_32.GPOUT_reg[18]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[18] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB16_rgbr_net_1 ), .EN(
        \CoreGPIO_0/GPOUT_reg_0_sqmuxa ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB6_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/GPOUT_reg[18] ));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_7_[2]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[2] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB6_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_7__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_208_i ), .ADn(VCC), .SLn(
        VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_7_rs[2] ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_125_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB7_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_7__1_sqmuxa ), .ALn(
        AFLSDF_INV_29_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(GND)
        , .Q(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_125_set_net_1 ));
    RGB \FCCC_0/GL1_INST/U0_RGB1_RGB6  (.An(\FCCC_0/GL1_INST/U0_YNn ), 
        .ENn(GND), .YL(\FCCC_0/GL1_INST/U0_RGB1_RGB6_rgbl_net_1 ), .YR(
        \FCCC_0/GL1_INST/U0_RGB1_RGB6_rgbr_net_1 ));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_88_set_RNICCUB  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_88_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_207_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_11_rs[0] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_11_[0]_net_1 ));
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_19  (
        .A(\reg_apb_wrp_0/reg16x8_0/mem_12_[3]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_495 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_19_net_1 ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_227  (.A(VCC), 
        .B(VCC), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[11] ), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[23] ), .IPC());
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_117  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_14_[5]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_503 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_117_net_1 ));
    CFG3 #( .INIT(8'h20) )  
        \CoreGPIO_0/xhdl1.GEN_BITS[25].APB_32.edge_both_RNO[25]  (.A(
        \CoreGPIO_0/CONFIG_reg[25][3] ), .B(
        \CoreAPB3_0_APBmslave3_PWDATA[25] ), .C(
        \CoreGPIO_0/edge_neg[25] ), .Y(\CoreGPIO_0/N_5911_i_0 ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_201_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_102_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_201_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_201_rs_net_1 ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_199  (.A(VCC), 
        .B(VCC), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[3] ), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[15] ), .IPC());
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_195  (.A(GND), 
        .B(VCC), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/F_AWID_HSEL0_net[3] ), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[11] ), .IPC());
    CFG3 #( .INIT(8'hF2) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_215  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_7_[6]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_498 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_215_i ));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_1_[4]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[4] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB14_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_1__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_140_i ), .ADn(VCC), .SLn(
        VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_1_rs[4] ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_248  (.A(VCC), 
        .B(GND), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[60] ), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/F_ARID_HSEL1_net[0] ), .IPC());
    CFG2 #( .INIT(4'h2) )  
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_a3_3[7]  (.A(
        \reg_apb_wrp_0/reg16x8_0/N_500 ), .B(
        \reg_apb_wrp_0/reg16x8_0/mem_13_[7]_net_1 ), .Y(
        \reg_apb_wrp_0/reg16x8_0/N_470 ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[3].APB_32.edge_both[3]  (.D(
        \CoreGPIO_0/edge_both_51_iv_i_0[3] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB9_rgbr_net_1 ), .EN(
        \CoreGPIO_0/edge_both_2_sqmuxa_12_i_1 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_YR ), .ADn(VCC), .SLn(
        VCC), .SD(GND), .LAT(GND), .Q(\CoreGPIO_0/edge_both[3] ));
    CFG4 #( .INIT(16'hFF4F) )  \CoreGPIO_0/edge_both_2_sqmuxa_23_i_0  
        (.A(\CoreGPIO_0.N_247 ), .B(\CoreGPIO_0/INTR_reg21 ), .C(
        \CoreGPIO_0/CONFIG_reg[5][3] ), .D(\CoreGPIO_0/N_139_i ), .Y(
        \CoreGPIO_0/N_76 ));
    CFG3 #( .INIT(8'hF2) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_188  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_6_[0]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_493 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_188_i ));
    CFG3 #( .INIT(8'h20) )  
        \CoreGPIO_0/xhdl1.GEN_BITS[18].APB_32.edge_both_RNO[18]  (.A(
        \CoreGPIO_0/CONFIG_reg[18][3] ), .B(
        \CoreAPB3_0_APBmslave3_PWDATA[18] ), .C(
        \CoreGPIO_0/edge_neg[18] ), .Y(\CoreGPIO_0/edge_neg_261[18] ));
    CFG2 #( .INIT(4'h7) )  \CoreGPIO_0/edge_both_2_sqmuxa_25_i  (.A(
        \CoreGPIO_0/N_248 ), .B(\CoreGPIO_0/CONFIG_reg[30][3] ), .Y(
        \CoreGPIO_0/edge_neg_2_sqmuxa_6_i_1 ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[2].REG_GEN.CONFIG_reg[2][1]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[1] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB16_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[2]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB6_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0.xhdl1.GEN_BITS[2].REG_GEN.CONFIG_reg[2][1] ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_269  (.A(VCC), 
        .B(GND), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[29] ), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/F_ARVALID_HWRITE1_net ), .IPC());
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[0].gpin3[0]  (.D(
        \CoreGPIO_0/gpin2[0] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB9_rgbr_net_1 ), .EN(VCC), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_YR ), .ADn(VCC), .SLn(
        VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0.xhdl1.GEN_BITS[0].gpin3[0] ));
    CFG4 #( .INIT(16'hAC0F) )  
        \CoreGPIO_0/CONFIG_reg_o_2_31_am_RNO[7]  (.A(
        \CoreGPIO_0/CONFIG_reg[10][7] ), .B(
        \CoreGPIO_0/CONFIG_reg[26][7] ), .C(
        \CoreGPIO_0/CONFIG_reg_o_2_10_1_1[7] ), .D(
        \CoreAPB3_0_APBmslave3_PADDR[5] ), .Y(
        \CoreGPIO_0/CONFIG_reg_o_2_31_am_RNO[7]_net_1 ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[30].REG_GEN.CONFIG_reg[30][4]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[4] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB14_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[30]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB4_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[30][4] ));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_180_rs_RNIRMOP  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_44_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_180_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_5_rs[4] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_5_[4]_net_1 ));
    INV_BA AFLSDF_INV_38 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_40_net_1 ), .Y(
        AFLSDF_INV_38_net_1));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/mem_4__RNI1LP21[1]  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_2_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_162_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_4_rs[1] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_4_[1]_net_1 ));
    IOBI_IB_OB_EB \FIC_MSS_0/MDDR_DQ_7_PAD/U_IOBI  (.D(VCC), .E(VCC), 
        .YIN(\FIC_MSS_0/MDDR_DQ_7_PAD/YIN ), .DOUT(), .EOUT(), .Y());
    CFG3 #( .INIT(8'hFD) )  \CoreGPIO_0/RDATA_32.un12_PRDATA_o_0_o2_1  
        (.A(\CoreAPB3_0_APBmslave3_PADDR[7] ), .B(
        \CoreAPB3_0_APBmslave3_PADDR[1] ), .C(
        \CoreAPB3_0_APBmslave3_PADDR[0] ), .Y(
        \CoreGPIO_0.RDATA_32.un12_PRDATA_o_0_o2_1 ));
    INV_BA AFLSDF_INV_49 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_123_net_1 ), .Y(
        AFLSDF_INV_49_net_1));
    CFG4 #( .INIT(16'h0F35) )  
        \CoreGPIO_0/CONFIG_reg_o_2_31_am_RNO_2[2]  (.A(
        \CoreGPIO_0/CONFIG_reg[6][2] ), .B(
        \CoreGPIO_0/CONFIG_reg[22][2] ), .C(
        \CoreAPB3_0_APBmslave3_PADDR[6] ), .D(
        \CoreAPB3_0_APBmslave3_PADDR[5] ), .Y(
        \CoreGPIO_0/CONFIG_reg_o_2_13_1_1[2] ));
    INV_BA AFLSDF_INV_120 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_13_net_1 ), .Y(
        AFLSDF_INV_120_net_1));
    CFG4 #( .INIT(16'h4000) )  
        \reg_apb_wrp_0/reg16x8_0/WRITE_GEN.mem_7__2_i_a2[6]  (.A(
        \CoreAPB3_0_APBmslave3_PADDR[3] ), .B(
        \CoreAPB3_0_APBmslave3_PADDR[2] ), .C(
        \CoreAPB3_0_APBmslave3_PADDR[0] ), .D(
        \CoreAPB3_0_APBmslave3_PADDR[1] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/N_498 ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[9].APB_32.INTR_reg[9]  (.D(
        \CoreGPIO_0/INTR_reg_126[9] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB14_rgbr_net_1 ), .EN(VCC), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB4_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/INTR_reg[9] ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[7].APB_32.INTR_reg[7]  (.D(
        \CoreGPIO_0/INTR_reg_100[7] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB11_rgbr_net_1 ), .EN(VCC), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB1_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/INTR_reg[7] ));
    CFG4 #( .INIT(16'h0010) )  
        \reg_apb_wrp_0/reg16x8_0/WRITE_GEN.mem_1__2_i_0_0_a2[5]  (.A(
        \CoreAPB3_0_APBmslave3_PADDR[3] ), .B(
        \CoreAPB3_0_APBmslave3_PADDR[2] ), .C(
        \CoreAPB3_0_APBmslave3_PADDR[0] ), .D(
        \CoreAPB3_0_APBmslave3_PADDR[1] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/N_502 ));
    INV_BA AFLSDF_INV_47 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_84_net_1 ), .Y(
        AFLSDF_INV_47_net_1));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_19  (.A(
        \FIC_MSS_0_FIC_0_APB_MASTER_PRDATA[24] ), .B(
        \FIC_MSS_0_FIC_0_APB_MASTER_PRDATA[31] ), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[24] ), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[31] ), .IPC());
    CFG3 #( .INIT(8'hF2) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_216  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_11_[5]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_505 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_216_i ));
    CFG4 #( .INIT(16'h1000) )  
        \CoreGPIO_0/xhdl1.GEN_BITS[28].REG_GEN.CONFIG_reg[28]2_0_a4_0_a2  
        (.A(\CoreAPB3_0_APBmslave3_PADDR[3] ), .B(
        \CoreAPB3_0_APBmslave3_PADDR[2] ), .C(\CoreGPIO_0/N_598 ), .D(
        \CoreGPIO_0/N_605 ), .Y(\CoreGPIO_0/CONFIG_reg[28]2 ));
    CFG4 #( .INIT(16'h330A) )  
        \CoreGPIO_0/xhdl1.GEN_BITS[7].APB_32.INTR_reg_100_0[7]  (.A(
        \CoreGPIO_0/INTR_reg[7] ), .B(
        \CoreGPIO_0/INTR_reg_100_0_o2_1[7] ), .C(
        \CoreAPB3_0_APBmslave3_PWDATA[7] ), .D(\CoreGPIO_0/N_248 ), .Y(
        \CoreGPIO_0/INTR_reg_100[7] ));
    CFG4 #( .INIT(16'h7350) )  
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_5[1]  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_14_[1]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/mem_6_[1]_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/N_503 ), .D(
        \reg_apb_wrp_0/reg16x8_0/N_493 ), .Y(
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_5[1]_net_1 ));
    CFG2 #( .INIT(4'h8) )  
        \CoreGPIO_0/xhdl1.GEN_BITS[3].REG_GPOUT.un34_GPIO_OUT_i  (.A(
        \CoreGPIO_0/GPOUT_reg[3] ), .B(\CoreGPIO_0/CONFIG_reg[3][0] ), 
        .Y(\GPIO_OUT_net_2[3] ));
    CFG2 #( .INIT(4'h2) )  \CoreGPIO_0/edge_pos_2_sqmuxa_5_i_a2  (.A(
        \CoreGPIO_0/gpin2[1] ), .B(
        \CoreGPIO_0.xhdl1.GEN_BITS[1].gpin3[1] ), .Y(
        \CoreGPIO_0/N_400 ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[23].REG_GEN.CONFIG_reg[23][4]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[4] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB10_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[23]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB0_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[23][4] ));
    RGB \FCCC_0/GL1_INST/U0_RGB1_RGB3  (.An(\FCCC_0/GL1_INST/U0_YNn ), 
        .ENn(GND), .YL(\FCCC_0/GL1_INST/U0_RGB1_RGB3_rgbl_net_1 ), .YR(
        ));
    INV_BA AFLSDF_INV_122 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_36_net_1 ), .Y(
        AFLSDF_INV_122_net_1));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_218  (.A(VCC), 
        .B(VCC), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[2] ), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[14] ), .IPC());
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/mem_12__RNICSF41[3]  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_19_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_227_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_12_rs[3] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_12_[3]_net_1 ));
    CFG4 #( .INIT(16'hAC0F) )  
        \CoreGPIO_0/CONFIG_reg_o_2_31_am_1_RNO_0[4]  (.A(
        \CoreGPIO_0/CONFIG_reg[8][4] ), .B(
        \CoreGPIO_0/CONFIG_reg[24][4] ), .C(
        \CoreGPIO_0/CONFIG_reg_o_2_3_1[4] ), .D(
        \CoreAPB3_0_APBmslave3_PADDR[5] ), .Y(
        \CoreGPIO_0/CONFIG_reg_o_2_31_am_1_RNO_0[4]_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_231_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_23_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_231_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_231_rs_net_1 ));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_set_RNIEHIN  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_161_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_4_rs[0] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_4_[0]_net_1 ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[27].APB_32.edge_both[27]  (.D(
        \CoreGPIO_0/N_5912_i_0 ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB9_rgbr_net_1 ), .EN(
        \CoreGPIO_0/N_161 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_YR ), .ADn(VCC), .SLn(
        VCC), .SD(GND), .LAT(GND), .Q(\CoreGPIO_0/edge_neg[27] ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_77_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB13_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_9__1_sqmuxa ), .ALn(
        AFLSDF_INV_30_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(GND)
        , .Q(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_77_set_net_1 ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[0].REG_GEN.CONFIG_reg[0][4]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[4] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB15_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[0]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB5_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[0][4] ));
    CFG2 #( .INIT(4'h4) )  \CoreGPIO_0/PRDATA_0_iv_0_a2_0[13]  (.A(
        \CoreGPIO_0.N_247 ), .B(\CoreGPIO_0/INTR_reg[13] ), .Y(
        \CoreGPIO_0.N_560 ));
    CFG2 #( .INIT(4'h2) )  
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_a3_13[0]  (.A(
        \reg_apb_wrp_0/reg16x8_0/N_499 ), .B(
        \reg_apb_wrp_0/reg16x8_0/mem_8_[0]_net_1 ), .Y(
        \reg_apb_wrp_0/reg16x8_0/N_368 ));
    CFG2 #( .INIT(4'h2) )  \CoreGPIO_0/edge_pos_2_sqmuxa_2_i_0_0_a2  (
        .A(\CoreGPIO_0/gpin2[6] ), .B(
        \CoreGPIO_0.xhdl1.GEN_BITS[6].gpin3[6] ), .Y(
        \CoreGPIO_0/N_689 ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_86_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB19_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_0__1_sqmuxa ), .ALn(
        AFLSDF_INV_31_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(GND)
        , .Q(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_86_set_net_1 ));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_58_set_RNIIPAE  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_58_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_253_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_15_rs[4] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_15_[4]_net_1 ));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/mem_7__RNI1ELO[2]  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_49_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_208_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_7_rs[2] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_7_[2]_net_1 ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[24].REG_GEN.CONFIG_reg[24][2]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[2] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB15_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[24]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB5_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[24][2] ));
    CFG4 #( .INIT(16'h7530) )  
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_0_1[5]  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_15_[5]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/mem_7_[5]_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/N_498 ), .D(
        \reg_apb_wrp_0/reg16x8_0/N_497 ), .Y(
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_0_1[5]_net_1 ));
    CFG4 #( .INIT(16'hF2F3) )  
        \CoreGPIO_0/xhdl1.GEN_BITS[28].APB_32.INTR_reg_373_0_o2_1_0[28]  
        (.A(\CoreGPIO_0/CONFIG_reg[28][6] ), .B(
        \CoreGPIO_0/edge_pos[28] ), .C(
        \CoreGPIO_0/INTR_reg_373_0_o2_0[28] ), .D(
        \CoreGPIO_0/CONFIG_reg[28][5] ), .Y(
        \CoreGPIO_0/INTR_reg_373_0_o2_1[28] ));
    CFG4 #( .INIT(16'hAA08) )  
        \CoreGPIO_0/xhdl1.GEN_BITS[5].APB_32.edge_both_79_iv_i_0[5]  (
        .A(\CoreGPIO_0/CONFIG_reg[5][3] ), .B(
        \CoreGPIO_0/edge_both[5] ), .C(
        \CoreAPB3_0_APBmslave3_PWDATA[5] ), .D(\CoreGPIO_0/N_139_i ), 
        .Y(\CoreGPIO_0/N_89 ));
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_15  (
        .A(\reg_apb_wrp_0/reg16x8_0/mem_5_[1]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_490 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_15_net_1 ));
    CFG4 #( .INIT(16'h8000) )  
        \CoreGPIO_0/xhdl1.GEN_BITS[23].REG_GEN.CONFIG_reg[23]2_0_a4_0_a2  
        (.A(\CoreAPB3_0_APBmslave3_PADDR[3] ), .B(
        \CoreAPB3_0_APBmslave3_PADDR[2] ), .C(\CoreGPIO_0/N_598 ), .D(
        \CoreGPIO_0/N_603 ), .Y(\CoreGPIO_0/CONFIG_reg[23]2 ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[15].REG_GEN.CONFIG_reg[15][3]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[3] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB10_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[15]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB0_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[15][3] ));
    CFG4 #( .INIT(16'h0F35) )  
        \CoreGPIO_0/CONFIG_reg_o_2_31_bm_1_RNO_1[4]  (.A(
        \CoreGPIO_0/CONFIG_reg[5][4] ), .B(
        \CoreGPIO_0/CONFIG_reg[21][4] ), .C(
        \CoreAPB3_0_APBmslave3_PADDR[6] ), .D(
        \CoreAPB3_0_APBmslave3_PADDR[5] ), .Y(
        \CoreGPIO_0/CONFIG_reg_o_2_21_1[4] ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[21].APB_32.GPOUT_reg[21]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[21] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB13_rgbr_net_1 ), .EN(
        \CoreGPIO_0/GPOUT_reg_0_sqmuxa ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB3_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0.xhdl1.GEN_BITS[21].APB_32.GPOUT_reg[21] ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_24  (.A(GND), 
        .B(VCC), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[0] ), .IPB(), .IPC());
    CFG3 #( .INIT(8'h20) )  
        \CoreGPIO_0/xhdl1.GEN_BITS[7].APB_32.edge_both_RNO[7]  (.A(
        \CoreGPIO_0/CONFIG_reg[7][3] ), .B(
        \CoreAPB3_0_APBmslave3_PWDATA[7] ), .C(
        \CoreGPIO_0/edge_pos[7] ), .Y(\CoreGPIO_0/N_83_i_0 ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_148_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_34_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_148_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_148_rs_net_1 ));
    CFG4 #( .INIT(16'hFFFE) )  
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_13[7]  (.A(
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_7[7]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_5[7]_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_6[7]_net_1 ), .D(
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_4[7]_net_1 ), .Y(
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_13[7]_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_55_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB18_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_3__1_sqmuxa ), .ALn(
        AFLSDF_INV_32_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(GND)
        , .Q(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_55_set_net_1 ));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_50_set_RNIP9UK  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_50_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_156_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_3_rs[4] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_3_[4]_net_1 ));
    CFG4 #( .INIT(16'hEAFA) )  \FIC_MSS_0/MSS_ADLIB_INST_RNO_3  (.A(
        \FIC_MSS_0/CoreAPB3_0_APBmslave5_PRDATA_m_0_1[4] ), .B(
        \CoreGPIO_0.PRDATA_iv_0_0_1[4] ), .C(
        CoreAPB3_0_APBmslave5_PSELx), .D(
        \FIC_MSS_0/CoreAPB3_0_APBmslave5_PRDATA_m_0_1_0[4] ), .Y(
        \FIC_MSS_0/FIC_MSS_0_FIC_0_APB_MASTER_PRDATA[4] ));
    CFG3 #( .INIT(8'hF2) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_142  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_1_[6]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_502 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_142_i ));
    sdf_IOPAD_TRI \FIC_MSS_0/MDDR_ADDR_12_PAD/U_IOPAD  (.PAD(
        MDDR_ADDR[12]), .D(\FIC_MSS_0/DRAM_ADDR_net_0[12] ), .E(
        \FIC_MSS_0/MDDR_ADDR_12_PAD/EOUT ));
    CFG4 #( .INIT(16'h0F35) )  
        \CoreGPIO_0/CONFIG_reg_o_2_31_am_1_RNO_2[6]  (.A(
        \CoreGPIO_0/CONFIG_reg[0][6] ), .B(
        \CoreGPIO_0/CONFIG_reg[16][6] ), .C(
        \CoreAPB3_0_APBmslave3_PADDR[6] ), .D(
        \CoreAPB3_0_APBmslave3_PADDR[5] ), .Y(
        \CoreGPIO_0/CONFIG_reg_o_2_3_1[6] ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[16].REG_GEN.CONFIG_reg[16][0]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[0] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB11_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[16]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB1_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[16][0] ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_204  (.A(VCC), 
        .B(GND), .C(GND), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[22] ), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/F_AWLEN_HBURST0_net[0] ), .IPC(
        \FIC_MSS_0/MSS_ADLIB_INST/F_AWVALID_HWRITE0_net ));
    CFG3 #( .INIT(8'hE2) )  \CoreGPIO_0/CONFIG_reg_o_2_31_ns[7]  (.A(
        \CoreGPIO_0/CONFIG_reg_o_2_31_am[7]_net_1 ), .B(
        \CoreAPB3_0_APBmslave3_PADDR[2] ), .C(
        \CoreGPIO_0/CONFIG_reg_o_2_31_bm[7]_net_1 ), .Y(
        \CoreGPIO_0.CONFIG_reg_o_2[7] ));
    CFG3 #( .INIT(8'hF2) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_183  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_9_[4]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_492 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_183_i ));
    CFG2 #( .INIT(4'h8) )  
        \reg_apb_wrp_0/reg16x8_0/mem_10__1_sqmuxa_0_a3  (.A(
        \reg_apb_wrp_0/reg16x8_0/N_491 ), .B(
        \reg_apb_wrp_0/wr_enable_net_1 ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_10__1_sqmuxa ));
    CFG4 #( .INIT(16'h5410) )  \CoreGPIO_0/PRDATA_iv_0_0_0_1[6]  (.A(
        \CoreAPB3_0_APBmslave3_PADDR[7] ), .B(
        \CoreAPB3_0_APBmslave3_PADDR[2] ), .C(
        \CoreGPIO_0/CONFIG_reg_o_2_31_am[6]_net_1 ), .D(
        \CoreGPIO_0/CONFIG_reg_o_2_31_bm[6]_net_1 ), .Y(
        \CoreGPIO_0.PRDATA_iv_0_0_0_0[6] ));
    INV_BA AFLSDF_INV_23 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_111_net_1 ), .Y(
        AFLSDF_INV_23_net_1));
    CFG2 #( .INIT(4'h2) )  
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_0_a3_11[5]  (.A(
        \reg_apb_wrp_0/reg16x8_0/N_492 ), .B(
        \reg_apb_wrp_0/reg16x8_0/mem_9_[5]_net_1 ), .Y(
        \reg_apb_wrp_0/reg16x8_0/N_350 ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_168  (.A(VCC), 
        .B(VCC), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/MMUART1_CTS_F2H_SCP_net ), .IPB(), 
        .IPC());
    INV_BA AFLSDF_INV_83 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_2_net_1 ), .Y(
        AFLSDF_INV_83_net_1));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_11_[3]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[3] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB16_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_11__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_212_i ), .ADn(VCC), .SLn(
        VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_11_rs[3] ));
    CFG4 #( .INIT(16'h2000) )  
        \CoreGPIO_0/xhdl1.GEN_BITS[5].REG_GEN.CONFIG_reg[5]2_0_a4_0_a2  
        (.A(\CoreAPB3_0_APBmslave3_PADDR[2] ), .B(
        \CoreAPB3_0_APBmslave3_PADDR[3] ), .C(\CoreGPIO_0/N_603 ), .D(
        \CoreGPIO_0/N_604 ), .Y(\CoreGPIO_0/CONFIG_reg[5]2 ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[0].APB_32.edge_neg[0]  (.D(
        \CoreGPIO_0/N_123 ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB9_rgbr_net_1 ), .EN(
        \CoreGPIO_0/N_52 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_YR ), .ADn(VCC), .SLn(
        VCC), .SD(GND), .LAT(GND), .Q(\CoreGPIO_0/edge_neg[0] ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_8_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB2_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_0__1_sqmuxa ), .ALn(
        AFLSDF_INV_33_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(GND)
        , .Q(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_8_set_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_47_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB14_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_1__1_sqmuxa ), .ALn(
        AFLSDF_INV_34_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(GND)
        , .Q(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_47_set_net_1 ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[25].REG_GEN.CONFIG_reg[25][6]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[6] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB15_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[25]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB5_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[25][6] ));
    CFG4 #( .INIT(16'hAC0F) )  
        \CoreGPIO_0/CONFIG_reg_o_2_31_bm_1_1_RNO[7]  (.A(
        \CoreGPIO_0/CONFIG_reg[13][7] ), .B(
        \CoreGPIO_0/CONFIG_reg[29][7] ), .C(
        \CoreGPIO_0/CONFIG_reg_o_2_21_1[7] ), .D(
        \CoreAPB3_0_APBmslave3_PADDR[5] ), .Y(
        \CoreGPIO_0/CONFIG_reg_o_2_31_bm_1_1_RNO[7]_net_1 ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_242  (.A(VCC), 
        .B(GND), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[54] ), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/F_WSTRB_net[2] ), .IPC());
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_67  (.A(GND), 
        .B(VCC), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[28] ), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[1] ), .IPC());
    CFG2 #( .INIT(4'h8) )  
        \reg_apb_wrp_0/reg16x8_0/mem_11__1_sqmuxa_0_a3  (.A(
        \reg_apb_wrp_0/reg16x8_0/N_505 ), .B(
        \reg_apb_wrp_0/wr_enable_net_1 ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_11__1_sqmuxa ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[21].REG_GEN.CONFIG_reg[21][5]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[5] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB13_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[21]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB3_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[21][5] ));
    INV_BA AFLSDF_INV_14 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_14_net_1 ), .Y(
        AFLSDF_INV_14_net_1));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_215_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_3_net_1 ), .EN(VCC), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_215_i ), .ADn(VCC), .SLn(
        VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_215_rs_net_1 ));
    CFG3 #( .INIT(8'hF2) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_197  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_10_[3]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_491 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_197_i ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[15].REG_GEN.CONFIG_reg[15][0]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[0] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB11_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[15]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB1_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[15][0] ));
    CFG3 #( .INIT(8'hF2) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_181  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_9_[3]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_492 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_181_i ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_128_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_81_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_128_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_128_rs_net_1 ));
    CFG2 #( .INIT(4'h2) )  
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_a3_5[6]  (.A(
        \reg_apb_wrp_0/reg16x8_0/N_495 ), .B(
        \reg_apb_wrp_0/reg16x8_0/mem_12_[6]_net_1 ), .Y(
        \reg_apb_wrp_0/reg16x8_0/N_452 ));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/mem_11__RNID3DK[5]  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_93_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_216_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_11_rs[5] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_11_[5]_net_1 ));
    INV_BA AFLSDF_INV_26 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_49_net_1 ), .Y(
        AFLSDF_INV_26_net_1));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[22].REG_GEN.CONFIG_reg[22][1]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[1] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB15_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[22]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB5_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[22][1] ));
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_63  (
        .A(\reg_apb_wrp_0/reg16x8_0/mem_15_[6]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_497 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_63_net_1 ));
    INV_BA AFLSDF_INV_86 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_60_net_1 ), .Y(
        AFLSDF_INV_86_net_1));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_212_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_91_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_212_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_212_rs_net_1 ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_21  (.A(
        \FIC_MSS_0_FIC_0_APB_MASTER_PRDATA[26] ), .B(GND), .C(VCC), 
        .IPA(\FIC_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[26] ), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_SIZE_net[0] ), .IPC());
    SLE \reg_apb_wrp_0/fsm[1]  (.D(\reg_apb_wrp_0/fsm_ns[1] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB12_rgbr_net_1 ), .EN(VCC), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB2_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/fsm[1]_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/temp_data[6]  (.D(
        \reg_apb_wrp_0/reg16x8_0/N_52_i_0 ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB12_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/rd_enable_net_1 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB2_rgbl_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/temp_data[6]_net_1 ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_147  (.A(VCC), 
        .B(VCC), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/I2C1_SDA_F2H_SCP_net ), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/MGPIO4A_F2H_GPIN_net ), .IPC());
    CFG4 #( .INIT(16'h0CAE) )  \CoreGPIO_0/PRDATA_0_iv_0_0_0[7]  (.A(
        \CoreGPIO_0/PRDATA_0_iv_0_0_a2_0_0[7]_net_1 ), .B(
        \CoreGPIO_0/INTR_reg[7] ), .C(\CoreGPIO_0.N_247 ), .D(
        \CoreGPIO_0.N_246 ), .Y(\CoreGPIO_0.PRDATA_0_iv_0_0_0[7] ));
    CFG4 #( .INIT(16'h0400) )  \CoreAPB3_0/iPSELS_raw23  (.A(
        \FIC_MSS_0_FIC_0_APB_MASTER_PADDR[31] ), .B(
        \FIC_MSS_0_FIC_0_APB_MASTER_PADDR[28] ), .C(
        \FIC_MSS_0_FIC_0_APB_MASTER_PADDR[30] ), .D(
        \FIC_MSS_0_FIC_0_APB_MASTER_PADDR[29] ), .Y(
        \CoreAPB3_0.iPSELS_raw23 ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[29].APB_32.INTR_reg[29]  (.D(
        \CoreGPIO_0/INTR_reg_386[29] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB11_rgbr_net_1 ), .EN(VCC), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB1_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/INTR_reg[29] ));
    CFG4 #( .INIT(16'hAC0F) )  
        \CoreGPIO_0/CONFIG_reg_o_2_31_bm_RNO[2]  (.A(
        \CoreGPIO_0/CONFIG_reg[11][2] ), .B(
        \CoreGPIO_0/CONFIG_reg[27][2] ), .C(
        \CoreGPIO_0/CONFIG_reg_o_2_25_1_1[2] ), .D(
        \CoreAPB3_0_APBmslave3_PADDR[5] ), .Y(
        \CoreGPIO_0/CONFIG_reg_o_2_31_bm_RNO[2]_net_1 ));
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_86  (
        .A(\reg_apb_wrp_0/reg16x8_0/mem_0_[5]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_496 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_86_net_1 ));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_66_set_RNI1G0Q  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_66_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_225_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_8_rs[3] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_8_[3]_net_1 ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_156  (.A(VCC), 
        .B(VCC), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/MGPIO9A_F2H_GPIN_net ), .IPB(), .IPC(
        ));
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_17  (
        .A(\reg_apb_wrp_0/reg16x8_0/mem_12_[1]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_495 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_17_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_15_[2]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[2] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB6_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_15__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_250_i ), .ADn(VCC), .SLn(
        VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_15_rs[2] ));
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_23  (
        .A(\reg_apb_wrp_0/reg16x8_0/mem_12_[7]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_495 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_23_net_1 ));
    CFG4 #( .INIT(16'hAC0F) )  
        \CoreGPIO_0/CONFIG_reg_o_2_31_bm_RNO[3]  (.A(
        \CoreGPIO_0/CONFIG_reg[11][3] ), .B(
        \CoreGPIO_0/CONFIG_reg[27][3] ), .C(
        \CoreGPIO_0/CONFIG_reg_o_2_25_1_1[3] ), .D(
        \CoreAPB3_0_APBmslave3_PADDR[5] ), .Y(
        \CoreGPIO_0/CONFIG_reg_o_2_31_bm_RNO[3]_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_169_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_69_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_169_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_169_rs_net_1 ));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/mem_6__RNI5OVQ[4]  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_37_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_196_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_6_rs[4] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_6_[4]_net_1 ));
    CFG4 #( .INIT(16'h0F35) )  
        \CoreGPIO_0/CONFIG_reg_o_2_31_bm_1_RNO_1[3]  (.A(
        \CoreGPIO_0/CONFIG_reg[5][3] ), .B(
        \CoreGPIO_0/CONFIG_reg[21][3] ), .C(
        \CoreAPB3_0_APBmslave3_PADDR[6] ), .D(
        \CoreAPB3_0_APBmslave3_PADDR[5] ), .Y(
        \CoreGPIO_0/CONFIG_reg_o_2_21_1[3] ));
    CFG4 #( .INIT(16'h7530) )  
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_7[7]  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_10_[7]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/mem_2_[7]_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/N_501 ), .D(
        \reg_apb_wrp_0/reg16x8_0/N_491 ), .Y(
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_7[7]_net_1 ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_75  (.A(VCC), 
        .B(VCC), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[9] ), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[16] ), .IPC());
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_38  (
        .A(\reg_apb_wrp_0/reg16x8_0/mem_2_[6]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_501 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_38_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_1_[2]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[2] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB15_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_1__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_138_i ), .ADn(VCC), .SLn(
        VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_1_rs[2] ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[16].REG_GEN.CONFIG_reg[16][3]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[3] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB11_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[16]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB1_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[16][3] ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_9  (.A(
        \FIC_MSS_0_FIC_0_APB_MASTER_PRDATA[7] ), .B(
        \FIC_MSS_0_FIC_0_APB_MASTER_PRDATA[14] ), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[7] ), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[14] ), .IPC());
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_212  (.A(VCC), 
        .B(GND), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[30] ), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/F_WID_HREADY01_net[0] ), .IPC());
    CFG4 #( .INIT(16'h0F35) )  
        \CoreGPIO_0/CONFIG_reg_o_2_31_bm_1_RNO_1[6]  (.A(
        \CoreGPIO_0/CONFIG_reg[5][6] ), .B(
        \CoreGPIO_0/CONFIG_reg[21][6] ), .C(
        \CoreAPB3_0_APBmslave3_PADDR[6] ), .D(
        \CoreAPB3_0_APBmslave3_PADDR[5] ), .Y(
        \CoreGPIO_0/CONFIG_reg_o_2_21_1[6] ));
    CFG4 #( .INIT(16'hEC00) )  \CoreAPB3_0/u_mux_p_to_b3/PRDATA[16]  (
        .A(\CoreGPIO_0.xhdl1.GEN_BITS[0].APB_32.GPOUT_reg9 ), .B(
        \CoreGPIO_0.N_554 ), .C(
        \CoreGPIO_0.xhdl1.GEN_BITS[16].APB_32.GPOUT_reg[16] ), .D(
        CoreAPB3_0_APBmslave5_PSELx), .Y(
        \FIC_MSS_0_FIC_0_APB_MASTER_PRDATA[16] ));
    CFG4 #( .INIT(16'hAC0F) )  
        \CoreGPIO_0/CONFIG_reg_o_2_31_am_RNO[5]  (.A(
        \CoreGPIO_0/CONFIG_reg[10][5] ), .B(
        \CoreGPIO_0/CONFIG_reg[26][5] ), .C(
        \CoreGPIO_0/CONFIG_reg_o_2_10_1_1[5] ), .D(
        \CoreAPB3_0_APBmslave3_PADDR[5] ), .Y(
        \CoreGPIO_0/CONFIG_reg_o_2_31_am_RNO[5]_net_1 ));
    CFG3 #( .INIT(8'h7F) )  \FIC_MSS_0/MSS_ADLIB_INST_RNO_15  (.A(
        \CoreGPIO_0.xhdl1.GEN_BITS[0].gpin3[0] ), .B(
        \CoreGPIO_0.RDATA_32.un12_PRDATA_o ), .C(
        \CoreGPIO_0.xhdl1.GEN_BITS[0].REG_GEN.CONFIG_reg[0][1] ), .Y(
        \FIC_MSS_0/CoreAPB3_0_APBmslave5_PRDATA_m_0_1[0] ));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_5_[4]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[4] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB6_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_5__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_180_i ), .ADn(VCC), .SLn(
        VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_5_rs[4] ));
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_96  (
        .A(\reg_apb_wrp_0/reg16x8_0/mem_10_[3]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_491 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_96_net_1 ));
    CFG4 #( .INIT(16'h0F35) )  
        \CoreGPIO_0/CONFIG_reg_o_2_31_bm_RNO_2[3]  (.A(
        \CoreGPIO_0/CONFIG_reg[7][3] ), .B(
        \CoreGPIO_0/CONFIG_reg[23][3] ), .C(
        \CoreAPB3_0_APBmslave3_PADDR[6] ), .D(
        \CoreAPB3_0_APBmslave3_PADDR[5] ), .Y(
        \CoreGPIO_0/CONFIG_reg_o_2_28_1_1[3] ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_164  (.A(VCC), 
        .B(VCC), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/MGPIO13A_F2H_GPIN_net ), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/MGPIO16A_F2H_GPIN_net ), .IPC());
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[2].APB_32.GPOUT_reg[2]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[2] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB16_rgbr_net_1 ), .EN(
        \CoreGPIO_0/GPOUT_reg_0_sqmuxa ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB6_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/GPOUT_reg[2] ));
    CFG4 #( .INIT(16'hB383) )  \CoreGPIO_0/CONFIG_reg_o_2_31_bm[3]  (
        .A(\CoreGPIO_0/CONFIG_reg_o_2_31_bm_RNO[3]_net_1 ), .B(
        \CoreGPIO_0/CONFIG_reg_o_2_31_bm_1[3] ), .C(
        \CoreAPB3_0_APBmslave3_PADDR[3] ), .D(
        \CoreGPIO_0/CONFIG_reg_o_2_31_bm_RNO_0[3]_net_1 ), .Y(
        \CONFIG_reg_o_2_31_bm[3] ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_153_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_124_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_153_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_153_rs_net_1 ));
    CFG2 #( .INIT(4'h7) )  \CoreGPIO_0/edge_both_2_sqmuxa_16_i  (.A(
        \CoreGPIO_0/N_248 ), .B(\CoreGPIO_0/CONFIG_reg[12][3] ), .Y(
        \CoreGPIO_0/N_188 ));
    CFG4 #( .INIT(16'hAA08) )  
        \CoreGPIO_0/xhdl1.GEN_BITS[3].APB_32.edge_pos_51_iv_i_0[3]  (
        .A(\CoreGPIO_0/CONFIG_reg[3][3] ), .B(\CoreGPIO_0/edge_pos[3] )
        , .C(\CoreAPB3_0_APBmslave3_PWDATA[3] ), .D(\CoreGPIO_0/N_687 )
        , .Y(\CoreGPIO_0/N_73 ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_176_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_40_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_176_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_176_rs_net_1 ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[1].APB_32.GPOUT_reg[1]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[1] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB16_rgbr_net_1 ), .EN(
        \CoreGPIO_0/GPOUT_reg_0_sqmuxa ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB6_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0.xhdl1.GEN_BITS[1].APB_32.GPOUT_reg[1] ));
    CFG4 #( .INIT(16'h7530) )  
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_1[1]  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_15_[1]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/mem_7_[1]_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/N_498 ), .D(
        \reg_apb_wrp_0/reg16x8_0/N_497 ), .Y(
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_1[1]_net_1 ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_117  (.A(VCC), 
        .B(VCC), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/FAB_RXACTIVE_net ), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/FAB_VSTATUS_net[6] ), .IPC());
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_251  (.A(VCC), 
        .B(GND), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[63] ), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/F_ARID_HSEL1_net[3] ), .IPC());
    CFG3 #( .INIT(8'hFE) )  
        \CoreGPIO_0/xhdl1.GEN_BITS[0].APB_32.un5_PRDATA_o_0_a2_0_o2_0  
        (.A(\CoreGPIO_0/N_243 ), .B(\CoreAPB3_0_APBmslave3_PADDR[4] ), 
        .C(\CoreGPIO_0.RDATA_32.un12_PRDATA_o_0_o2_1 ), .Y(
        \CoreGPIO_0.N_246 ));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_197_rs_RNIL735  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_96_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_197_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_10_rs[3] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_10_[3]_net_1 ));
    CFG4 #( .INIT(16'h330A) )  
        \CoreGPIO_0/xhdl1.GEN_BITS[13].APB_32.INTR_reg_178_0[13]  (.A(
        \CoreGPIO_0/INTR_reg[13] ), .B(
        \CoreGPIO_0/INTR_reg_178_0_o2_1[13] ), .C(
        \CoreAPB3_0_APBmslave3_PWDATA[13] ), .D(\CoreGPIO_0/N_248 ), 
        .Y(\CoreGPIO_0/INTR_reg_178[13] ));
    RGB \FCCC_0/GL1_INST/U0_RGB1_RGB10  (.An(
        \FCCC_0/GL1_INST/U0_YNn_GSouth ), .ENn(GND), .YL(
        \FCCC_0/GL1_INST/U0_RGB1_RGB10_rgbl_net_1 ), .YR(
        \FCCC_0/GL1_INST/U0_RGB1_RGB10_rgbr_net_1 ));
    CFG3 #( .INIT(8'hF2) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_207  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_11_[0]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_505 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_207_i ));
    CFG2 #( .INIT(4'h8) )  \FIC_MSS_0/MSS_ADLIB_INST_RNO_25  (.A(
        CoreAPB3_0_APBmslave5_PSELx), .B(
        \CoreGPIO_0.xhdl1.GEN_BITS[5].APB_32.INTR_reg[5] ), .Y(
        \FIC_MSS_0/CoreAPB3_0_APBmslave5_PRDATA_m_c_c_0[5] ));
    INV_BA AFLSDF_INV_129 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_32_net_1 ), .Y(
        AFLSDF_INV_129_net_1));
    CFG4 #( .INIT(16'h7350) )  
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_3[4]  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_11_[4]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/mem_3_[4]_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/N_505 ), .D(
        \reg_apb_wrp_0/reg16x8_0/N_494 ), .Y(
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_3[4]_net_1 ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[29].REG_GEN.CONFIG_reg[29][7]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[7] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB13_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[29]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB3_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[29][7] ));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_3_[5]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[5] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB10_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_3__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_157_i ), .ADn(VCC), .SLn(
        VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_3_rs[5] ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_153  (.A(VCC), 
        .B(VCC), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/CAN_RXBUS_F2H_SCP_net ), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/MGPIO7A_F2H_GPIN_net ), .IPC());
    CFG3 #( .INIT(8'hF2) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_201  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_10_[5]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_491 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_201_i ));
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_122  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_3_[0]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_494 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_122_net_1 ));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_131_rs_RNIEHEP  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_80_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_131_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_0_rs[0] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_0_[0]_net_1 ));
    sdf_IOPAD_BI \FIC_MSS_0/MDDR_DQ_8_PAD/U_IOPAD  (.PAD(MDDR_DQ[8]), 
        .D(\FIC_MSS_0/DRAM_DQ_OUT_net_0[8] ), .E(
        \FIC_MSS_0/DRAM_DQ_OE_net_0[8] ), .Y(
        \FIC_MSS_0/MDDR_DQ_8_PAD_Y ));
    CFG3 #( .INIT(8'h20) )  
        \CoreGPIO_0/xhdl1.GEN_BITS[14].APB_32.edge_both_RNO[14]  (.A(
        \CoreGPIO_0/CONFIG_reg[14][3] ), .B(
        \CoreAPB3_0_APBmslave3_PWDATA[14] ), .C(
        \CoreGPIO_0/edge_neg[14] ), .Y(\CoreGPIO_0/edge_neg_205[14] ));
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_3  (
        .A(\reg_apb_wrp_0/reg16x8_0/mem_7_[6]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_498 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_3_net_1 ));
    CFG3 #( .INIT(8'hF2) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_157  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_3_[5]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_494 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_157_i ));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_11_[5]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[5] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB19_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_11__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_216_i ), .ADn(VCC), .SLn(
        VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_11_rs[5] ));
    CFG3 #( .INIT(8'hF2) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_255  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_15_[6]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_497 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_255_i ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_263  (.A(VCC), 
        .B(VCC), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[11] ), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[23] ), .IPC());
    CFG4 #( .INIT(16'h0F35) )  
        \CoreGPIO_0/CONFIG_reg_o_2_31_bm_RNO_1[5]  (.A(
        \CoreGPIO_0/CONFIG_reg[3][5] ), .B(
        \CoreGPIO_0/CONFIG_reg[19][5] ), .C(
        \CoreAPB3_0_APBmslave3_PADDR[6] ), .D(
        \CoreAPB3_0_APBmslave3_PADDR[5] ), .Y(
        \CoreGPIO_0/CONFIG_reg_o_2_25_1_1[5] ));
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_81  (
        .A(\reg_apb_wrp_0/reg16x8_0/mem_0_[1]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_496 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_81_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_65_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB11_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_4__1_sqmuxa ), .ALn(
        AFLSDF_INV_35_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(GND)
        , .Q(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_65_set_net_1 ));
    INV_BA AFLSDF_INV_59 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_35_net_1 ), .Y(
        AFLSDF_INV_59_net_1));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[16].APB_32.GPOUT_reg[16]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[16] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB9_rgbr_net_1 ), .EN(
        \CoreGPIO_0/GPOUT_reg_0_sqmuxa ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_YR ), .ADn(VCC), .SLn(
        VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0.xhdl1.GEN_BITS[16].APB_32.GPOUT_reg[16] ));
    CFG4 #( .INIT(16'hBBFB) )  \CoreGPIO_0/edge_pos_2_sqmuxa_5_i_0  (
        .A(\CoreGPIO_0/N_400 ), .B(\CoreGPIO_0/CONFIG_reg[1][3] ), .C(
        \CoreGPIO_0/INTR_reg21 ), .D(\CoreGPIO_0.N_247 ), .Y(
        \CoreGPIO_0/N_66 ));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_11_[4]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[4] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB19_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_11__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_214_i ), .ADn(VCC), .SLn(
        VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_11_rs[4] ));
    SLE \reg_apb_wrp_0/wr_enable  (.D(\reg_apb_wrp_0/N_70 ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB12_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/N_45_i_0 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB2_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/wr_enable_net_1 ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[9].REG_GEN.CONFIG_reg[9][7]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[7] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB14_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[9]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB4_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[9][7] ));
    CFG4 #( .INIT(16'hEC00) )  \CoreAPB3_0/u_mux_p_to_b3/PRDATA[13]  (
        .A(\CoreGPIO_0.xhdl1.GEN_BITS[0].APB_32.GPOUT_reg9 ), .B(
        \CoreGPIO_0.N_560 ), .C(
        \CoreGPIO_0.xhdl1.GEN_BITS[13].APB_32.GPOUT_reg[13] ), .D(
        CoreAPB3_0_APBmslave5_PSELx), .Y(
        \FIC_MSS_0_FIC_0_APB_MASTER_PRDATA[13] ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_255_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_63_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_255_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_255_rs_net_1 ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[28].REG_GEN.CONFIG_reg[28][2]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[2] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB14_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[28]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB4_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[28][2] ));
    INV_BA AFLSDF_INV_57 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_76_net_1 ), .Y(
        AFLSDF_INV_57_net_1));
    INV_BA AFLSDF_INV_105 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_66_net_1 ), .Y(
        AFLSDF_INV_105_net_1));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[3].gpin3[3]  (.D(
        \CoreGPIO_0/gpin2[3] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB9_rgbr_net_1 ), .EN(VCC), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_YR ), .ADn(VCC), .SLn(
        VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0.xhdl1.GEN_BITS[3].gpin3[3] ));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_113_set_RNIJIQI  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_113_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_241_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_14_rs[1] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_14_[1]_net_1 ));
    CFG4 #( .INIT(16'hFFFE) )  
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_0_13[5]  (.A(
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_0_7[5]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_0_5[5]_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_0_6[5]_net_1 ), .D(
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_0_4[5]_net_1 ), .Y(
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_0_13[5]_net_1 ));
    CFG4 #( .INIT(16'h330A) )  
        \CoreGPIO_0/xhdl1.GEN_BITS[25].APB_32.INTR_reg_334_0[25]  (.A(
        \CoreGPIO_0/INTR_reg[25] ), .B(
        \CoreGPIO_0/INTR_reg_334_0_o2_1[25] ), .C(
        \CoreAPB3_0_APBmslave3_PWDATA[25] ), .D(\CoreGPIO_0/N_248 ), 
        .Y(\CoreGPIO_0/INTR_reg_334[25] ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_70_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB14_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_8__1_sqmuxa ), .ALn(
        AFLSDF_INV_36_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(GND)
        , .Q(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_70_set_net_1 ));
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_91  (
        .A(\reg_apb_wrp_0/reg16x8_0/mem_11_[3]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_505 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_91_net_1 ));
    INV_BA AFLSDF_INV_63 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_124_net_1 ), .Y(
        AFLSDF_INV_63_net_1));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_13_[0]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[0] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB10_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_13__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_232_i ), .ADn(VCC), .SLn(
        VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_13_rs[0] ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_252_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_60_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_252_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_252_rs_net_1 ));
    CFG3 #( .INIT(8'h40) )  \CoreGPIO_0/PRDATA_0_iv_0_a2[10]  (.A(
        \CoreGPIO_0.N_246 ), .B(\CoreGPIO_0/GPOUT_reg[10] ), .C(
        \CoreAPB3_0_APBmslave3_PADDR[5] ), .Y(\CoreGPIO_0.N_565 ));
    CFG4 #( .INIT(16'hAC0F) )  
        \CoreGPIO_0/CONFIG_reg_o_2_31_bm_RNO[7]  (.A(
        \CoreGPIO_0/CONFIG_reg[11][7] ), .B(
        \CoreGPIO_0/CONFIG_reg[27][7] ), .C(
        \CoreGPIO_0/CONFIG_reg_o_2_25_1_1[7] ), .D(
        \CoreAPB3_0_APBmslave3_PADDR[5] ), .Y(
        \CoreGPIO_0/CONFIG_reg_o_2_31_bm_RNO[7]_net_1 ));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_181_rs_RNI3SOU  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_75_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_181_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_9_rs[3] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_9_[3]_net_1 ));
    CFG4 #( .INIT(16'h4000) )  
        \CoreGPIO_0/xhdl1.GEN_BITS[13].REG_GEN.CONFIG_reg[13]2_0_a4_0_a2  
        (.A(\CoreAPB3_0_APBmslave3_PADDR[3] ), .B(
        \CoreAPB3_0_APBmslave3_PADDR[2] ), .C(\CoreGPIO_0/N_604 ), .D(
        \CoreGPIO_0/N_605 ), .Y(\CoreGPIO_0/CONFIG_reg[13]2 ));
    IP_INTERFACE \FCCC_0/CCC_INST/IP_INTERFACE_9  (.A(VCC), .B(GND), 
        .C(VCC), .IPA(\FCCC_0/CCC_INST/PLL_BYPASS_N_net ), .IPB(
        \FCCC_0/CCC_INST/NGMUX3_SEL_net ), .IPC(
        \FCCC_0/CCC_INST/PWDATA_net[7] ));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/mem_2__RNIN1DH[3]  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_32_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_147_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_2_rs[3] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_2_[3]_net_1 ));
    INV_BA AFLSDF_INV_30 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_77_net_1 ), .Y(
        AFLSDF_INV_30_net_1));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[7].REG_GEN.CONFIG_reg[7][2]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[2] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB11_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[7]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB1_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[7][2] ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_1_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB3_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_7__1_sqmuxa ), .ALn(
        AFLSDF_INV_37_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(GND)
        , .Q(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_1_set_net_1 ));
    CFG3 #( .INIT(8'hF2) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_177  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_9_[1]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_492 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_177_i ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[12].APB_32.edge_both[12]  (.D(
        \CoreGPIO_0/edge_neg_177[12] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB12_rgbr_net_1 ), .EN(
        \CoreGPIO_0/N_188 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB2_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/edge_neg[12] ));
    INV_BA AFLSDF_INV_92 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_48_net_1 ), .Y(
        AFLSDF_INV_92_net_1));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_3_[7]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[7] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB17_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_3__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_160_i ), .ADn(VCC), .SLn(
        VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_3_rs[7] ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_57  (.A(GND), 
        .B(GND), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[11] ), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[18] ), .IPC());
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_174_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_15_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_174_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_174_rs_net_1 ));
    INV_BA AFLSDF_INV_66 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_102_net_1 ), .Y(
        AFLSDF_INV_66_net_1));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_218_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_94_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_218_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_218_rs_net_1 ));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/mem_10__RNILCFV[2]  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_99_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_195_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_10_rs[2] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_10_[2]_net_1 ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[6].gpin2[6]  (.D(
        \CoreGPIO_0/gpin1[6] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB12_rgbr_net_1 ), .EN(VCC), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB2_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(\CoreGPIO_0/gpin2[6] )
        );
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_40_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB5_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_5__1_sqmuxa ), .ALn(
        AFLSDF_INV_38_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(GND)
        , .Q(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_40_set_net_1 ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[22].APB_32.GPOUT_reg[22]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[22] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB13_rgbr_net_1 ), .EN(
        \CoreGPIO_0/GPOUT_reg_0_sqmuxa ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB3_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0.xhdl1.GEN_BITS[22].APB_32.GPOUT_reg[22] ));
    CFG4 #( .INIT(16'hBBFB) )  \CoreGPIO_0/edge_pos_2_sqmuxa_4_i_0  (
        .A(\CoreGPIO_0/N_398 ), .B(\CoreGPIO_0/CONFIG_reg[4][3] ), .C(
        \CoreGPIO_0/INTR_reg21 ), .D(\CoreGPIO_0.N_247 ), .Y(
        \CoreGPIO_0/N_68 ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_68  (.A(GND), 
        .B(VCC), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[29] ), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[2] ), .IPC());
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[16].REG_GEN.CONFIG_reg[16][5]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[5] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB11_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[16]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB1_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[16][5] ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[22].REG_GEN.CONFIG_reg[22][4]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[4] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB14_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[22]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB4_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[22][4] ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_73_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB13_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_9__1_sqmuxa ), .ALn(
        AFLSDF_INV_39_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(GND)
        , .Q(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_73_set_net_1 ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[28].APB_32.INTR_reg[28]  (.D(
        \CoreGPIO_0/INTR_reg_373[28] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB13_rgbr_net_1 ), .EN(VCC), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB3_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/INTR_reg[28] ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_258  (.A(VCC), 
        .B(VCC), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[6] ), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[18] ), .IPC());
    INV_BA AFLSDF_INV_113 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_85_net_1 ), .Y(
        AFLSDF_INV_113_net_1));
    CFG4 #( .INIT(16'h7530) )  
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_4[3]  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_12_[3]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/mem_4_[3]_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/N_504 ), .D(
        \reg_apb_wrp_0/reg16x8_0/N_495 ), .Y(
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_4[3]_net_1 ));
    CFG4 #( .INIT(16'h0F35) )  
        \CoreGPIO_0/CONFIG_reg_o_2_31_am_1_RNO_2[1]  (.A(
        \CoreGPIO_0.xhdl1.GEN_BITS[0].REG_GEN.CONFIG_reg[0][1] ), .B(
        \CoreGPIO_0/CONFIG_reg[16][1] ), .C(
        \CoreAPB3_0_APBmslave3_PADDR[6] ), .D(
        \CoreAPB3_0_APBmslave3_PADDR[5] ), .Y(
        \CoreGPIO_0/CONFIG_reg_o_2_3_1[1] ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_91_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB17_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_11__1_sqmuxa ), .ALn(
        AFLSDF_INV_40_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(GND)
        , .Q(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_91_set_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_12_[3]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[3] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB2_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_12__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_227_i ), .ADn(VCC), .SLn(
        VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_12_rs[3] ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[15].REG_GEN.CONFIG_reg[15][7]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[7] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB10_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[15]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB0_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[15][7] ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_47  (.A(VCC), 
        .B(GND), .C(VCC), .IPA(), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[1] ), .IPC());
    INV_BA AFLSDF_INV_44 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_110_net_1 ), .Y(
        AFLSDF_INV_44_net_1));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_112_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB6_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_14__1_sqmuxa ), .ALn(
        AFLSDF_INV_41_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(GND)
        , .Q(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_112_set_net_1 ));
    CFG3 #( .INIT(8'hF2) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_149  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_2_[5]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_501 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_149_i ));
    sdf_IOPADP_BI \FIC_MSS_0/MDDR_DQS_1_PAD/U_IOPADP  (.PAD_P(
        MDDR_DQS[1]), .N2PIN_P(\FIC_MSS_0/MDDR_DQS_1_PAD/U2_N2P ), 
        .OIN_P(\FIC_MSS_0/DRAM_DQS_OUT_net_0[1] ), .EIN_P(
        \FIC_MSS_0/DRAM_DQS_OE_net_0[1] ), .IOUT_P(
        \FIC_MSS_0/MDDR_DQS_1_PAD_Y ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[3].APB_32.edge_neg[3]  (.D(
        \CoreGPIO_0/edge_neg_51_iv_i_1[3] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB9_rgbr_net_1 ), .EN(
        \CoreGPIO_0/N_81 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_YR ), .ADn(VCC), .SLn(
        VCC), .SD(GND), .LAT(GND), .Q(\CoreGPIO_0/edge_neg[3] ));
    RGB \FCCC_0/GL1_INST/U0_RGB1_RGB8  (.An(\FCCC_0/GL1_INST/U0_YNn ), 
        .ENn(GND), .YL(\FCCC_0/GL1_INST/U0_RGB1_RGB8_rgbl_net_1 ), .YR(
        \FCCC_0/GL1_INST/U0_RGB1_RGB8_rgbr_net_1 ));
    CFG4 #( .INIT(16'h4000) )  
        \CoreGPIO_0/xhdl1.GEN_BITS[25].REG_GEN.CONFIG_reg[25]2_0_a4_0_a2  
        (.A(\CoreAPB3_0_APBmslave3_PADDR[3] ), .B(
        \CoreAPB3_0_APBmslave3_PADDR[2] ), .C(\CoreGPIO_0/N_598 ), .D(
        \CoreGPIO_0/N_610 ), .Y(\CoreGPIO_0/CONFIG_reg[25]2 ));
    CFG4 #( .INIT(16'hCC0A) )  
        \CoreGPIO_0/xhdl1.GEN_BITS[5].APB_32.INTR_reg_74_0_0[5]  (.A(
        \CoreGPIO_0.xhdl1.GEN_BITS[5].APB_32.INTR_reg[5] ), .B(
        \CoreGPIO_0/N_1579_tz ), .C(\CoreAPB3_0_APBmslave3_PWDATA[5] ), 
        .D(\CoreGPIO_0/N_248 ), .Y(\CoreGPIO_0/INTR_reg_74[5] ));
    CFG4 #( .INIT(16'h330A) )  
        \CoreGPIO_0/xhdl1.GEN_BITS[24].APB_32.INTR_reg_321_0[24]  (.A(
        \CoreGPIO_0/INTR_reg[24] ), .B(
        \CoreGPIO_0/INTR_reg_321_0_o2_1[24] ), .C(
        \CoreAPB3_0_APBmslave3_PWDATA[24] ), .D(\CoreGPIO_0/N_248 ), 
        .Y(\CoreGPIO_0/INTR_reg_321[24] ));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_5_[2]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[2] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB6_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_5__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_176_i ), .ADn(VCC), .SLn(
        VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_5_rs[2] ));
    IOENFF_BYPASS \GPIO_OUT_obuf[4]/U0/U_IOENFF  (.A(
        \GPIO_OUT_obuf[4]/U0/EOUT1 ), .Y(\GPIO_OUT_obuf[4]/U0/EOUT ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_82_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB11_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_0__1_sqmuxa ), .ALn(
        AFLSDF_INV_42_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(GND)
        , .Q(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_82_set_net_1 ));
    CFG4 #( .INIT(16'hC5CA) )  
        \CoreGPIO_0/xhdl1.GEN_BITS[6].APB_32.INTR_reg_87_0_0_m2[6]  (
        .A(\CoreGPIO_0.xhdl1.GEN_BITS[6].gpin3[6] ), .B(
        \CoreGPIO_0/INTR_reg_87_0_0_m2_0[6] ), .C(
        \CoreGPIO_0/CONFIG_reg[6][6] ), .D(
        \CoreGPIO_0/CONFIG_reg[6][5] ), .Y(
        \CoreGPIO_0/INTR_reg_87_0_0_m2[6] ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_126_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB17_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_3__1_sqmuxa ), .ALn(
        AFLSDF_INV_43_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(GND)
        , .Q(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_126_set_net_1 ));
    sdf_IOPAD_TRI \FIC_MSS_0/MDDR_BA_2_PAD/U_IOPAD  (.PAD(MDDR_BA[2]), 
        .D(\FIC_MSS_0/DRAM_BA_net_0[2] ), .E(
        \FIC_MSS_0/MDDR_BA_2_PAD/EOUT ));
    CFG4 #( .INIT(16'h4000) )  
        \CoreGPIO_0/xhdl1.GEN_BITS[17].REG_GEN.CONFIG_reg[17]2_0_a4_0_a2  
        (.A(\CoreAPB3_0_APBmslave3_PADDR[3] ), .B(
        \CoreAPB3_0_APBmslave3_PADDR[2] ), .C(\CoreGPIO_0/N_598 ), .D(
        \CoreGPIO_0/N_606 ), .Y(\CoreGPIO_0/CONFIG_reg[17]2 ));
    CFG2 #( .INIT(4'h7) )  \CoreGPIO_0/edge_both_2_sqmuxa_10_i  (.A(
        \CoreGPIO_0/N_248 ), .B(\CoreGPIO_0/CONFIG_reg[18][3] ), .Y(
        \CoreGPIO_0/N_192 ));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_8_[6]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[6] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB12_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_8__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_171_i ), .ADn(VCC), .SLn(
        VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_8_rs[6] ));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/mem_12__RNI6V831[7]  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_23_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_231_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_12_rs[7] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_12_[7]_net_1 ));
    IOTRI_OB_EB \FIC_MSS_0/MDDR_BA_1_PAD/U_IOOUT  (.D(VCC), .E(VCC), 
        .DOUT(), .EOUT(\FIC_MSS_0/MDDR_BA_1_PAD/EOUT ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_186_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_27_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_186_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_186_rs_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_110_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB11_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_13__1_sqmuxa ), .ALn(
        AFLSDF_INV_44_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(GND)
        , .Q(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_110_set_net_1 ));
    CFG2 #( .INIT(4'h7) )  \CoreGPIO_0/edge_both_2_sqmuxa_2_i  (.A(
        \CoreGPIO_0/N_248 ), .B(\CoreGPIO_0/CONFIG_reg[13][3] ), .Y(
        \CoreGPIO_0/edge_pos_2_sqmuxa_9_i_1 ));
    INV_BA AFLSDF_INV_75 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_113_net_1 ), .Y(
        AFLSDF_INV_75_net_1));
    CFG4 #( .INIT(16'h135F) )  
        \CoreAPB3_0/u_mux_p_to_b3/PRDATA_0_iv_1[7]  (.A(
        \CoreAPB3_0_APBmslave3_PRDATA[7] ), .B(
        CoreAPB3_0_APBmslave5_PSELx), .C(CoreAPB3_0_APBmslave3_PSELx), 
        .D(\CoreGPIO_0.PRDATA_0_iv_0_0_0[7] ), .Y(
        \CoreAPB3_0/u_mux_p_to_b3/PRDATA_0_iv_1[7]_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_43_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB15_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_1__1_sqmuxa ), .ALn(
        AFLSDF_INV_45_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(GND)
        , .Q(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_43_set_net_1 ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[6].REG_GEN.CONFIG_reg[6][1]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[1] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB15_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[6]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB5_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0.xhdl1.GEN_BITS[6].REG_GEN.CONFIG_reg[6][1] ));
    CFG4 #( .INIT(16'hAC0F) )  
        \CoreGPIO_0/CONFIG_reg_o_2_31_am_1_1_RNO[6]  (.A(
        \CoreGPIO_0/CONFIG_reg[12][6] ), .B(
        \CoreGPIO_0/CONFIG_reg[28][6] ), .C(
        \CoreGPIO_0/CONFIG_reg_o_2_6_1[6] ), .D(
        \CoreAPB3_0_APBmslave3_PADDR[5] ), .Y(
        \CoreGPIO_0/CONFIG_reg_o_2_31_am_1_1_RNO[6]_net_1 ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[20].REG_GEN.CONFIG_reg[20][0]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[0] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB12_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[20]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB2_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[20][0] ));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_251_rs_RNI9R3P  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_61_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_251_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_15_rs[3] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_15_[3]_net_1 ));
    CFG2 #( .INIT(4'h4) )  \CoreGPIO_0/PRDATA_0_iv_0_a2_0[14]  (.A(
        \CoreGPIO_0.N_247 ), .B(\CoreGPIO_0/INTR_reg[14] ), .Y(
        \CoreGPIO_0.N_558 ));
    INV_BA AFLSDF_INV_18 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_80_net_1 ), .Y(
        AFLSDF_INV_18_net_1));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/mem_3__RNI159N[0]  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_122_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_152_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_3_rs[0] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_3_[0]_net_1 ));
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_89  (
        .A(\reg_apb_wrp_0/reg16x8_0/mem_11_[1]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_505 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_89_net_1 ));
    CFG3 #( .INIT(8'hF2) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_138  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_1_[2]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_502 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_138_i ));
    IP_INTERFACE \FCCC_0/CCC_INST/IP_INTERFACE_12  (.A(VCC), .B(VCC), 
        .C(VCC), .IPA(\FCCC_0/CCC_INST/NGMUX0_ARST_N_net ), .IPB(), 
        .IPC(\FCCC_0/CCC_INST/PADDR_net[2] ));
    CFG4 #( .INIT(16'h1000) )  
        \CoreGPIO_0/xhdl1.GEN_BITS[3].REG_INT.un34_intr_u_ns_1  (.A(
        \CoreGPIO_0/CONFIG_reg[3][6] ), .B(
        \CoreGPIO_0/CONFIG_reg[3][5] ), .C(\CoreGPIO_0/edge_both[3] ), 
        .D(\CoreGPIO_0/CONFIG_reg[3][7] ), .Y(
        \CoreGPIO_0/un34_intr_u_ns_1 ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_239  (.A(VCC), 
        .B(VCC), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[37] ), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[49] ), .IPC());
    CFG3 #( .INIT(8'hF2) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_140  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_1_[4]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_502 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_140_i ));
    SLE \reg_apb_wrp_0/reg16x8_0/data_out[4]  (.D(
        \reg_apb_wrp_0/reg16x8_0/temp_data[4]_net_1 ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB13_rgbr_net_1 ), .EN(VCC), .ALn(
        VCC), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreAPB3_0_APBmslave3_PRDATA[4] ));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_2_[1]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[1] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB2_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_2__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_145_i ), .ADn(VCC), .SLn(
        VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_2_rs[1] ));
    IOTRI_OB_EB \FIC_MSS_0/MDDR_ADDR_2_PAD/U_IOOUT  (.D(VCC), .E(VCC), 
        .DOUT(), .EOUT(\FIC_MSS_0/MDDR_ADDR_2_PAD/EOUT ));
    CFG4 #( .INIT(16'hEFEE) )  
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_0_9[5]  (.A(
        \reg_apb_wrp_0/reg16x8_0/N_350 ), .B(
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_0_3[5]_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_1_[5]_net_1 ), .D(
        \reg_apb_wrp_0/reg16x8_0/N_502 ), .Y(
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_0_9[5]_net_1 ));
    RGB \FCCC_0/GL1_INST/U0_RGB1_RGB1  (.An(\FCCC_0/GL1_INST/U0_YNn ), 
        .ENn(GND), .YL(\FCCC_0/GL1_INST/U0_RGB1_RGB1_rgbl_net_1 ), .YR(
        \FCCC_0/GL1_INST/U0_RGB1_RGB1_rgbr_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_101_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB9_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_10__1_sqmuxa ), .ALn(
        AFLSDF_INV_46_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(GND)
        , .Q(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_101_set_net_1 ));
    CFG4 #( .INIT(16'hC480) )  
        \CoreGPIO_0/xhdl1.GEN_BITS[5].APB_32.INTR_reg_74_0_0_RNO[5]  (
        .A(\CoreGPIO_0/CONFIG_reg[5][7] ), .B(
        \CoreGPIO_0/CONFIG_reg[5][3] ), .C(
        \CoreGPIO_0/INTR_reg_74_0_0_54_tz_1 ), .D(
        \CoreGPIO_0/INTR_reg_74_0_0_m2[5] ), .Y(\CoreGPIO_0/N_1579_tz )
        );
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[16].APB_32.INTR_reg[16]  (.D(
        \CoreGPIO_0/INTR_reg_217[16] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB10_rgbr_net_1 ), .EN(VCC), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB0_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/INTR_reg[16] ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[18].REG_GEN.CONFIG_reg[18][5]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[5] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB17_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[18]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB7_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[18][5] ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[5].REG_GEN.CONFIG_reg[5][1]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[1] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB13_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[5]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB3_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0.xhdl1.GEN_BITS[5].REG_GEN.CONFIG_reg[5][1] ));
    RGB \FCCC_0/GL1_INST/U0_RGB1_RGB5  (.An(\FCCC_0/GL1_INST/U0_YNn ), 
        .ENn(GND), .YL(\FCCC_0/GL1_INST/U0_RGB1_RGB5_rgbl_net_1 ), .YR(
        \FCCC_0/GL1_INST/U0_RGB1_RGB5_rgbr_net_1 ));
    CFG4 #( .INIT(16'h7350) )  
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_5[7]  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_14_[7]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/mem_6_[7]_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/N_503 ), .D(
        \reg_apb_wrp_0/reg16x8_0/N_493 ), .Y(
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_5[7]_net_1 ));
    CFG3 #( .INIT(8'hF2) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_145  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_2_[1]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_501 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_145_i ));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_9_[5]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[5] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB13_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_9__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_185_i ), .ADn(VCC), .SLn(
        VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_9_rs[5] ));
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_99  (
        .A(\reg_apb_wrp_0/reg16x8_0/mem_10_[2]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_491 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_99_net_1 ));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_242_rs_RNIMQ38  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_114_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_242_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_14_rs[2] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_14_[2]_net_1 ));
    CFG4 #( .INIT(16'hAC0F) )  
        \CoreGPIO_0/CONFIG_reg_o_2_31_bm_1_RNO_0[1]  (.A(
        \CoreGPIO_0/CONFIG_reg[9][1] ), .B(
        \CoreGPIO_0/CONFIG_reg[25][1] ), .C(
        \CoreGPIO_0/CONFIG_reg_o_2_18_1[1] ), .D(
        \CoreAPB3_0_APBmslave3_PADDR[5] ), .Y(
        \CoreGPIO_0/CONFIG_reg_o_2_31_bm_1_RNO_0[1]_net_1 ));
    IOIN_IB \GPIO_IN_ibuf[2]/U0/U_IOIN  (.YIN(\GPIO_IN_ibuf[2]/U0/YIN )
        , .E(GND), .Y(\GPIO_IN_c[2] ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_25  (.A(GND), 
        .B(VCC), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[1] ), .IPB(), .IPC());
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[22].REG_GEN.CONFIG_reg[22][0]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[0] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB14_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[22]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB4_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[22][0] ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_165_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_65_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_165_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_165_rs_net_1 ));
    CFG4 #( .INIT(16'hAC0F) )  
        \CoreGPIO_0/CONFIG_reg_o_2_31_am_RNO_0[0]  (.A(
        \CoreGPIO_0/CONFIG_reg[14][0] ), .B(
        \CoreGPIO_0/CONFIG_reg[30][0] ), .C(
        \CoreGPIO_0/CONFIG_reg_o_2_13_1_1[0] ), .D(
        \CoreAPB3_0_APBmslave3_PADDR[5] ), .Y(
        \CoreGPIO_0/CONFIG_reg_o_2_31_am_RNO_0[0]_net_1 ));
    CFG4 #( .INIT(16'hFFF8) )  \FIC_MSS_0/MSS_ADLIB_INST_RNO_10  (.A(
        CoreAPB3_0_APBmslave3_PSELx), .B(
        \CoreAPB3_0_APBmslave3_PRDATA[4] ), .C(
        \FIC_MSS_0/CoreAPB3_0_APBmslave5_PRDATA_m_c_c[4] ), .D(
        \FIC_MSS_0/CoreAPB3_0_APBmslave5_PRDATA_m_c_d[4] ), .Y(
        \FIC_MSS_0/CoreAPB3_0_APBmslave5_PRDATA_m_0_1[4] ));
    CFG2 #( .INIT(4'h2) )  
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_a3_3[6]  (.A(
        \reg_apb_wrp_0/reg16x8_0/N_500 ), .B(
        \reg_apb_wrp_0/reg16x8_0/mem_13_[6]_net_1 ), .Y(
        \reg_apb_wrp_0/reg16x8_0/N_450 ));
    INV_BA AFLSDF_INV_3 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_16_net_1 ), .Y(
        AFLSDF_INV_3_net_1));
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_18  (
        .A(\reg_apb_wrp_0/reg16x8_0/mem_12_[2]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_495 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_18_net_1 ));
    CFG3 #( .INIT(8'hDF) )  \CoreGPIO_0/edge_neg_2_sqmuxa_9_i_0  (.A(
        \CoreGPIO_0/CONFIG_reg[3][3] ), .B(\CoreGPIO_0/N_686 ), .C(
        \CoreGPIO_0/N_248 ), .Y(\CoreGPIO_0/N_81 ));
    IOOUTFF_BYPASS \GPIO_OUT_obuf[2]/U0/U_IOOUTFF  (.A(
        \GPIO_OUT_obuf[2]/U0/DOUT1 ), .Y(\GPIO_OUT_obuf[2]/U0/DOUT ));
    CFG4 #( .INIT(16'hA9FF) )  
        \CoreGPIO_0/xhdl1.GEN_BITS[27].APB_32.INTR_reg_360_0_o2_0_0[27]  
        (.A(\CoreGPIO_0/CONFIG_reg[27][7] ), .B(
        \CoreGPIO_0/CONFIG_reg[27][6] ), .C(
        \CoreGPIO_0/CONFIG_reg[27][5] ), .D(
        \CoreGPIO_0/CONFIG_reg[27][3] ), .Y(
        \CoreGPIO_0/INTR_reg_360_0_o2_0[27] ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_252  (.A(VCC), 
        .B(VCC), .C(GND), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[0] ), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[12] ), .IPC(
        \FIC_MSS_0/MSS_ADLIB_INST/F_ARSIZE_HSIZE1_net[0] ));
    CFG3 #( .INIT(8'hF2) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_230  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_12_[6]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_495 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_230_i ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_179  (.A(VCC), 
        .B(VCC), .C(VCC), .IPA(), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/MGPIO21B_F2H_GPIN_net ), .IPC());
    CFG4 #( .INIT(16'h0F35) )  
        \CoreGPIO_0/CONFIG_reg_o_2_31_am_RNO_2[6]  (.A(
        \CoreGPIO_0/CONFIG_reg[6][6] ), .B(
        \CoreGPIO_0/CONFIG_reg[22][6] ), .C(
        \CoreAPB3_0_APBmslave3_PADDR[6] ), .D(
        \CoreAPB3_0_APBmslave3_PADDR[5] ), .Y(
        \CoreGPIO_0/CONFIG_reg_o_2_13_1_1[6] ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_175  (.A(VCC), 
        .B(VCC), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/MMUART1_SCK_F2H_SCP_net ), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/MGPIO19B_F2H_GPIN_net ), .IPC());
    CFG4 #( .INIT(16'hAC0F) )  
        \CoreGPIO_0/CONFIG_reg_o_2_31_bm_RNO[5]  (.A(
        \CoreGPIO_0/CONFIG_reg[11][5] ), .B(
        \CoreGPIO_0/CONFIG_reg[27][5] ), .C(
        \CoreGPIO_0/CONFIG_reg_o_2_25_1_1[5] ), .D(
        \CoreAPB3_0_APBmslave3_PADDR[5] ), .Y(
        \CoreGPIO_0/CONFIG_reg_o_2_31_bm_RNO[5]_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_12_[5]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[5] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB10_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_12__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_229_i ), .ADn(VCC), .SLn(
        VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_12_rs[5] ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_82  (.A(VCC), 
        .B(VCC), .C(VCC), .IPA(), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[23] ), .IPC());
    IOINFF_BYPASS \FIC_MSS_0/MDDR_DQ_0_PAD/U_IOINFF  (.A(
        \FIC_MSS_0/MDDR_DQ_0_PAD_Y ), .Y(\FIC_MSS_0/MDDR_DQ_0_PAD/YIN )
        );
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[5].APB_32.edge_neg[5]  (.D(
        \CoreGPIO_0/N_115 ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB10_rgbr_net_1 ), .EN(
        \CoreGPIO_0/N_60 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB0_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/edge_neg[5] ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_140  (.A(VCC), 
        .B(VCC), .C(VCC), .IPA(\FIC_MSS_0/MSS_ADLIB_INST/RX_EV_net ), 
        .IPB(\FIC_MSS_0/MSS_ADLIB_INST/USER_MSS_GPIO_RESET_N_net ), 
        .IPC());
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_246  (.A(VCC), 
        .B(GND), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[58] ), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/F_WSTRB_net[6] ), .IPC());
    CFG4 #( .INIT(16'h0F35) )  
        \CoreGPIO_0/CONFIG_reg_o_2_31_am_RNO_2[7]  (.A(
        \CoreGPIO_0/CONFIG_reg[6][7] ), .B(
        \CoreGPIO_0/CONFIG_reg[22][7] ), .C(
        \CoreAPB3_0_APBmslave3_PADDR[6] ), .D(
        \CoreAPB3_0_APBmslave3_PADDR[5] ), .Y(
        \CoreGPIO_0/CONFIG_reg_o_2_13_1_1[7] ));
    CFG2 #( .INIT(4'h7) )  \CoreGPIO_0/edge_both_2_sqmuxa_9_i  (.A(
        \CoreGPIO_0/N_248 ), .B(\CoreGPIO_0/CONFIG_reg[19][3] ), .Y(
        \CoreGPIO_0/N_194 ));
    CFG3 #( .INIT(8'hF2) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_232  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_13_[0]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_500 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_232_i ));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_79_set_RNIJ8A81  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_79_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_189_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_9_rs[7] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_9_[7]_net_1 ));
    CFG3 #( .INIT(8'h4C) )  \FIC_MSS_0/MSS_ADLIB_INST_RNO_20  (.A(
        \CoreGPIO_0.xhdl1.GEN_BITS[0].APB_32.GPOUT_reg9 ), .B(
        \FIC_MSS_0/CoreAPB3_0_APBmslave5_PRDATA_m_0_1_0[6] ), .C(
        \CoreGPIO_0.xhdl1.GEN_BITS[6].APB_32.GPOUT_reg[6] ), .Y(
        \FIC_MSS_0/CoreAPB3_0_APBmslave5_PRDATA_m_0_1_1[6] ));
    CFG3 #( .INIT(8'hF2) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_129  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_0_[2]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_496 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_129_i ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_260  (.A(VCC), 
        .B(VCC), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[8] ), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[20] ), .IPC());
    SLE \reg_apb_wrp_0/reg16x8_0/mem_12_[4]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[4] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB5_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_12__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_228_i ), .ADn(VCC), .SLn(
        VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_12_rs[4] ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[23].REG_GEN.CONFIG_reg[23][3]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[3] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB10_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[23]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB0_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[23][3] ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_184_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_25_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_184_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_184_rs_net_1 ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_157  (.A(VCC), 
        .B(VCC), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/SPI0_SS2_F2H_SCP_net ), .IPB(), .IPC(
        ));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_175_rs_RNI0LC21  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_72_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_175_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_9_rs[0] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_9_[0]_net_1 ));
    CFG4 #( .INIT(16'h330A) )  
        \CoreGPIO_0/xhdl1.GEN_BITS[19].APB_32.INTR_reg_256_0[19]  (.A(
        \CoreGPIO_0/INTR_reg[19] ), .B(
        \CoreGPIO_0/INTR_reg_256_0_o2_1[19] ), .C(
        \CoreAPB3_0_APBmslave3_PWDATA[19] ), .D(\CoreGPIO_0/N_248 ), 
        .Y(\CoreGPIO_0/INTR_reg_256[19] ));
    INV_BA AFLSDF_INV_116 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_64_net_1 ), .Y(
        AFLSDF_INV_116_net_1));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_138  (.A(VCC), 
        .B(VCC), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/SMBALERT_NI1_net ), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/F2_DMAREADY_net[0] ), .IPC());
    CFG4 #( .INIT(16'hB383) )  \CoreGPIO_0/CONFIG_reg_o_2_31_bm[1]  (
        .A(\CoreGPIO_0/CONFIG_reg_o_2_31_bm_RNO[1]_net_1 ), .B(
        \CoreGPIO_0/CONFIG_reg_o_2_31_bm_1[1] ), .C(
        \CoreAPB3_0_APBmslave3_PADDR[3] ), .D(
        \CoreGPIO_0/CONFIG_reg_o_2_31_bm_RNO_0[1]_net_1 ), .Y(
        \CoreGPIO_0/CONFIG_reg_o_2_31_bm[1]_net_1 ));
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_85  (
        .A(\reg_apb_wrp_0/reg16x8_0/mem_0_[4]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_496 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_85_net_1 ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_196  (.A(VCC), 
        .B(VCC), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[0] ), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[12] ), .IPC());
    CFG3 #( .INIT(8'hF2) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_133  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_0_[5]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_496 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_133_i ));
    CFG3 #( .INIT(8'hB8) )  
        \CoreGPIO_0/xhdl1.GEN_BITS[6].APB_32.INTR_reg_87_0_0_m2_0[6]  
        (.A(\CoreGPIO_0/edge_neg[6] ), .B(
        \CoreGPIO_0/CONFIG_reg[6][5] ), .C(\CoreGPIO_0/edge_pos[6] ), 
        .Y(\CoreGPIO_0/INTR_reg_87_0_0_m2_0[6] ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[13].REG_GEN.CONFIG_reg[13][2]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[2] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB14_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[13]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB4_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[13][2] ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_267  (.A(VCC), 
        .B(GND), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[27] ), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/F_ARLOCK_HMASTLOCK1_net[1] ), .IPC());
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[0].REG_GEN.CONFIG_reg[0][5]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[5] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB11_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[0]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB1_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[0][5] ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_84_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB9_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_0__1_sqmuxa ), .ALn(
        AFLSDF_INV_47_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(GND)
        , .Q(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_84_set_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_9_[7]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[7] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB16_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_9__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_189_i ), .ADn(VCC), .SLn(
        VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_9_rs[7] ));
    IOBI_IB_OB_EB \FIC_MSS_0/MDDR_DQ_12_PAD/U_IOBI  (.D(VCC), .E(VCC), 
        .YIN(\FIC_MSS_0/MDDR_DQ_12_PAD/YIN ), .DOUT(), .EOUT(), .Y());
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_79  (.A(VCC), 
        .B(VCC), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[13] ), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[20] ), .IPC());
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_17  (.A(
        \FIC_MSS_0_FIC_0_APB_MASTER_PRDATA[22] ), .B(
        \FIC_MSS_0_FIC_0_APB_MASTER_PRDATA[29] ), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[22] ), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[29] ), .IPC());
    IOIN_IB \MSS_RESET_N_F2M_ibuf/U0/U_IOIN  (.YIN(
        \MSS_RESET_N_F2M_ibuf/U0/YIN ), .E(GND), .Y(
        MSS_RESET_N_F2M_ibuf));
    CFG4 #( .INIT(16'h7530) )  
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_1[6]  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_15_[6]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/mem_7_[6]_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/N_498 ), .D(
        \reg_apb_wrp_0/reg16x8_0/N_497 ), .Y(
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_1[6]_net_1 ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[4].APB_32.edge_pos[4]  (.D(
        \CoreGPIO_0/N_103 ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB12_rgbr_net_1 ), .EN(
        \CoreGPIO_0/N_68 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB2_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/edge_pos[4] ));
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_1  (
        .A(\reg_apb_wrp_0/reg16x8_0/mem_7_[7]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_498 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_1_net_1 ));
    CFG3 #( .INIT(8'hB8) )  
        \CoreGPIO_0/xhdl1.GEN_BITS[2].APB_32.INTR_reg_35_0_m2_0[2]  (
        .A(\CoreGPIO_0/edge_neg[2] ), .B(\CoreGPIO_0/CONFIG_reg[2][5] )
        , .C(\CoreGPIO_0/edge_pos[2] ), .Y(\CoreGPIO_0/N_173 ));
    IOOUTFF_BYPASS \GPIO_OUT_obuf[5]/U0/U_IOOUTFF  (.A(
        \GPIO_OUT_obuf[5]/U0/DOUT1 ), .Y(\GPIO_OUT_obuf[5]/U0/DOUT ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_58  (.A(VCC), 
        .B(GND), .C(VCC), .IPA(), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[19] ), .IPC());
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_95  (
        .A(\reg_apb_wrp_0/reg16x8_0/mem_11_[7]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_505 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_95_net_1 ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_110  (.A(VCC), 
        .B(VCC), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/FAB_XDATAIN_net[2] ), .IPB(), .IPC());
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_120  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_2_[7]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_501 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_120_net_1 ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_216  (.A(VCC), 
        .B(VCC), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[0] ), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[12] ), .IPC(
        \FIC_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[24] ));
    CFG4 #( .INIT(16'h4000) )  
        \CoreGPIO_0/xhdl1.GEN_BITS[29].REG_GEN.CONFIG_reg[29]2_0_a4_0_a2  
        (.A(\CoreAPB3_0_APBmslave3_PADDR[3] ), .B(
        \CoreAPB3_0_APBmslave3_PADDR[2] ), .C(\CoreGPIO_0/N_598 ), .D(
        \CoreGPIO_0/N_605 ), .Y(\CoreGPIO_0/CONFIG_reg[29]2 ));
    CFG4 #( .INIT(16'h0F35) )  
        \CoreGPIO_0/CONFIG_reg_o_2_31_am_RNO_1[7]  (.A(
        \CoreGPIO_0/CONFIG_reg[2][7] ), .B(
        \CoreGPIO_0/CONFIG_reg[18][7] ), .C(
        \CoreAPB3_0_APBmslave3_PADDR[6] ), .D(
        \CoreAPB3_0_APBmslave3_PADDR[5] ), .Y(
        \CoreGPIO_0/CONFIG_reg_o_2_10_1_1[7] ));
    sdf_IOPAD_BI \FIC_MSS_0/MDDR_DQ_15_PAD/U_IOPAD  (.PAD(MDDR_DQ[15]), 
        .D(\FIC_MSS_0/DRAM_DQ_OUT_net_0[15] ), .E(
        \FIC_MSS_0/DRAM_DQ_OE_net_0[15] ), .Y(
        \FIC_MSS_0/MDDR_DQ_15_PAD_Y ));
    CFG3 #( .INIT(8'h04) )  
        \CoreGPIO_0/xhdl1.GEN_BITS[2].REG_GEN.CONFIG_reg[2]2_0_a4_0_a2_1  
        (.A(\CoreAPB3_0_APBmslave3_PADDR[6] ), .B(
        \CoreGPIO_0/INTR_reg21 ), .C(\CoreAPB3_0_APBmslave3_PADDR[7] ), 
        .Y(\CoreGPIO_0/N_604 ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_7_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB8_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_8__1_sqmuxa ), .ALn(
        AFLSDF_INV_48_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(GND)
        , .Q(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_7_set_net_1 ));
    CFG3 #( .INIT(8'hF2) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_131  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_0_[0]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_496 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_131_i ));
    CFG4 #( .INIT(16'hC480) )  
        \CoreGPIO_0/xhdl1.GEN_BITS[4].APB_32.INTR_reg_61_0_0_RNO[4]  (
        .A(\CoreGPIO_0/CONFIG_reg[4][7] ), .B(
        \CoreGPIO_0/CONFIG_reg[4][3] ), .C(
        \CoreGPIO_0/INTR_reg_61_0_0_53_tz_1 ), .D(\CoreGPIO_0/N_179 ), 
        .Y(\CoreGPIO_0/N_1578_tz ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_209_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_89_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_209_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_209_rs_net_1 ));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_21_set_RNI99FV  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_21_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_229_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_12_rs[5] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_12_[5]_net_1 ));
    CFG4 #( .INIT(16'h330A) )  
        \CoreGPIO_0/xhdl1.GEN_BITS[10].APB_32.INTR_reg_139_0[10]  (.A(
        \CoreGPIO_0.xhdl1.GEN_BITS[10].APB_32.INTR_reg[10] ), .B(
        \CoreGPIO_0/INTR_reg_139_0_o2_1[10] ), .C(
        \CoreAPB3_0_APBmslave3_PWDATA[10] ), .D(\CoreGPIO_0/N_248 ), 
        .Y(\CoreGPIO_0/INTR_reg_139[10] ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_146_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_30_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_146_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_146_rs_net_1 ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[22].REG_GEN.CONFIG_reg[22][2]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[2] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB14_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[22]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB4_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[22][2] ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_123_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB8_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_6__1_sqmuxa ), .ALn(
        AFLSDF_INV_49_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(GND)
        , .Q(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_123_set_net_1 ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[14].REG_GEN.CONFIG_reg[14][6]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[6] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB13_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[14]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB3_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[14][6] ));
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_125  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_7_[0]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_498 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_125_net_1 ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_48  (.A(GND), 
        .B(VCC), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[2] ), .IPB(), .IPC());
    CFG4 #( .INIT(16'hA9FF) )  
        \CoreGPIO_0/xhdl1.GEN_BITS[17].APB_32.INTR_reg_230_0_o2_0_0[17]  
        (.A(\CoreGPIO_0/CONFIG_reg[17][7] ), .B(
        \CoreGPIO_0/CONFIG_reg[17][6] ), .C(
        \CoreGPIO_0/CONFIG_reg[17][5] ), .D(
        \CoreGPIO_0/CONFIG_reg[17][3] ), .Y(
        \CoreGPIO_0/INTR_reg_230_0_o2_0[17] ));
    INV_BA AFLSDF_INV_71 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_93_net_1 ), .Y(
        AFLSDF_INV_71_net_1));
    CFG3 #( .INIT(8'hF2) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_204  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_7_[0]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_498 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_204_i ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_193  (.A(GND), 
        .B(VCC), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/F_AWID_HSEL0_net[1] ), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[9] ), .IPC(
        \FIC_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[21] ));
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_33  (
        .A(\reg_apb_wrp_0/reg16x8_0/mem_6_[2]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_493 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_33_net_1 ));
    RGB \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB6  (.An(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_YNn_GSouth ), .ENn(GND), .YL()
        , .YR(\MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB6_rgbr_net_1 ));
    sdf_IOPAD_IN \GPIO_IN_ibuf[6]/U0/U_IOPAD  (.PAD(GPIO_IN[6]), .Y(
        \GPIO_IN_ibuf[6]/U0/YIN1 ));
    CFG4 #( .INIT(16'h0F35) )  
        \CoreGPIO_0/CONFIG_reg_o_2_31_bm_RNO_2[5]  (.A(
        \CoreGPIO_0/CONFIG_reg[7][5] ), .B(
        \CoreGPIO_0/CONFIG_reg[23][5] ), .C(
        \CoreAPB3_0_APBmslave3_PADDR[6] ), .D(
        \CoreAPB3_0_APBmslave3_PADDR[5] ), .Y(
        \CoreGPIO_0/CONFIG_reg_o_2_28_1_1[5] ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_171_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_70_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_171_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_171_rs_net_1 ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[27].REG_GEN.CONFIG_reg[27][1]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[1] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB10_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[27]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB0_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[27][1] ));
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_87  (
        .A(\reg_apb_wrp_0/reg16x8_0/mem_0_[6]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_496 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_87_net_1 ));
    INV_BA AFLSDF_INV_54 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_25_net_1 ), .Y(
        AFLSDF_INV_54_net_1));
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_70  (
        .A(\reg_apb_wrp_0/reg16x8_0/mem_8_[6]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_499 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_70_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_4_[0]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[0] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB17_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_4__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_161_i ), .ADn(VCC), .SLn(
        VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_4_rs[0] ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_134  (.A(VCC), 
        .B(VCC), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/I2C0_BCLK_net ), .IPB(), .IPC());
    CFG4 #( .INIT(16'hA9FF) )  
        \CoreGPIO_0/xhdl1.GEN_BITS[24].APB_32.INTR_reg_321_0_o2_0_0[24]  
        (.A(\CoreGPIO_0/CONFIG_reg[24][7] ), .B(
        \CoreGPIO_0/CONFIG_reg[24][6] ), .C(
        \CoreGPIO_0/CONFIG_reg[24][5] ), .D(
        \CoreGPIO_0/CONFIG_reg[24][3] ), .Y(
        \CoreGPIO_0/INTR_reg_321_0_o2_0[24] ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[30].REG_GEN.CONFIG_reg[30][7]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[7] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB12_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[30]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB2_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[30][7] ));
    CFG3 #( .INIT(8'hDF) )  \CoreGPIO_0/edge_neg_2_sqmuxa_i_0_0  (.A(
        \CoreGPIO_0/CONFIG_reg[6][3] ), .B(\CoreGPIO_0/N_688 ), .C(
        \CoreGPIO_0/N_248 ), .Y(\CoreGPIO_0/N_62 ));
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_104  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_13_[0]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_500 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_104_net_1 ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[10].REG_GEN.CONFIG_reg[10][1]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[1] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB16_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[10]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB6_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[10][1] ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_172_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_13_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_172_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_172_rs_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_8_[3]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[3] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB8_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_8__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_225_i ), .ADn(VCC), .SLn(
        VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_8_rs[3] ));
    CFG4 #( .INIT(16'hA9FF) )  
        \CoreGPIO_0/xhdl1.GEN_BITS[12].APB_32.INTR_reg_165_0_o2_0_0[12]  
        (.A(\CoreGPIO_0/CONFIG_reg[12][7] ), .B(
        \CoreGPIO_0/CONFIG_reg[12][6] ), .C(
        \CoreGPIO_0/CONFIG_reg[12][5] ), .D(
        \CoreGPIO_0/CONFIG_reg[12][3] ), .Y(
        \CoreGPIO_0/INTR_reg_165_0_o2_0[12] ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_157_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_52_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_157_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_157_rs_net_1 ));
    IOINFF_BYPASS \FIC_MSS_0/MDDR_DQ_4_PAD/U_IOINFF  (.A(
        \FIC_MSS_0/MDDR_DQ_4_PAD_Y ), .Y(\FIC_MSS_0/MDDR_DQ_4_PAD/YIN )
        );
    INV_BA AFLSDF_INV_114 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_104_net_1 ), .Y(
        AFLSDF_INV_114_net_1));
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_97  (
        .A(\reg_apb_wrp_0/reg16x8_0/mem_10_[0]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_491 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_97_net_1 ));
    RGB \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB3  (.An(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_YNn_GSouth ), .ENn(GND), .YL()
        , .YR(\MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB3_rgbr_net_1 ));
    CFG3 #( .INIT(8'hF2) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_187  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_9_[6]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_492 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_187_i ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_99_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB14_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_10__1_sqmuxa ), .ALn(
        AFLSDF_INV_50_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(GND)
        , .Q(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_99_set_net_1 ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_244  (.A(VCC), 
        .B(GND), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[56] ), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/F_WSTRB_net[4] ), .IPC());
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[26].REG_GEN.CONFIG_reg[26][2]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[2] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB16_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[26]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB6_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[26][2] ));
    INV_BA AFLSDF_INV_48 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_7_net_1 ), .Y(
        AFLSDF_INV_48_net_1));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_239_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_111_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_239_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_239_rs_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_51_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB3_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_7__1_sqmuxa ), .ALn(
        AFLSDF_INV_51_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(GND)
        , .Q(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_51_set_net_1 ));
    IOINFF_BYPASS \FIC_MSS_0/MDDR_DQ_5_PAD/U_IOINFF  (.A(
        \FIC_MSS_0/MDDR_DQ_5_PAD_Y ), .Y(\FIC_MSS_0/MDDR_DQ_5_PAD/YIN )
        );
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[4].REG_GEN.CONFIG_reg[4][2]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[2] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB14_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[4]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB4_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[4][2] ));
    sdf_IOPAD_TRI \FIC_MSS_0/MDDR_CS_N_PAD/U_IOPAD  (.PAD(MDDR_CS_N), 
        .D(\FIC_MSS_0/MSS_ADLIB_INST_DRAM_CSN ), .E(
        \FIC_MSS_0/MDDR_CS_N_PAD/EOUT ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_233  (.A(VCC), 
        .B(VCC), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[31] ), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[43] ), .IPC());
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_127_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB7_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_7__1_sqmuxa ), .ALn(
        AFLSDF_INV_52_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(GND)
        , .Q(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_127_set_net_1 ));
    CFG4 #( .INIT(16'h4657) )  
        \CoreGPIO_0/CONFIG_reg_o_2_31_am_1_1[7]  (.A(
        \CoreAPB3_0_APBmslave3_PADDR[4] ), .B(
        \CoreAPB3_0_APBmslave3_PADDR[3] ), .C(
        \CoreGPIO_0/CONFIG_reg_o_2_31_am_1_1_RNO[7]_net_1 ), .D(
        \CoreGPIO_0/CONFIG_reg_o_2_31_am_1_RNO_0[7]_net_1 ), .Y(
        \CoreGPIO_0/CONFIG_reg_o_2_31_am_1[7] ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[16].APB_32.edge_both[16]  (.D(
        \CoreGPIO_0/edge_neg_233[16] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB9_rgbr_net_1 ), .EN(
        \CoreGPIO_0/edge_pos_2_sqmuxa_29_i_1 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_YR ), .ADn(VCC), .SLn(
        VCC), .SD(GND), .LAT(GND), .Q(\CoreGPIO_0/edge_neg[16] ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[8].REG_GEN.CONFIG_reg[8][1]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[1] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB15_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[8]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB5_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[8][1] ));
    CFG4 #( .INIT(16'h0F35) )  
        \CoreGPIO_0/CONFIG_reg_o_2_31_am_RNO_1[2]  (.A(
        \CoreGPIO_0/CONFIG_reg[2][2] ), .B(
        \CoreGPIO_0/CONFIG_reg[18][2] ), .C(
        \CoreAPB3_0_APBmslave3_PADDR[6] ), .D(
        \CoreAPB3_0_APBmslave3_PADDR[5] ), .Y(
        \CoreGPIO_0/CONFIG_reg_o_2_10_1_1[2] ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[25].REG_GEN.CONFIG_reg[25][7]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[7] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB14_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[25]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB4_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[25][7] ));
    CFG4 #( .INIT(16'hC5CA) )  
        \CoreGPIO_0/xhdl1.GEN_BITS[4].APB_32.INTR_reg_61_0_m2[4]  (.A(
        \CoreGPIO_0.xhdl1.GEN_BITS[4].gpin3[4] ), .B(
        \CoreGPIO_0/N_172 ), .C(\CoreGPIO_0/CONFIG_reg[4][6] ), .D(
        \CoreGPIO_0/CONFIG_reg[4][5] ), .Y(\CoreGPIO_0/N_179 ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_209  (.A(VCC), 
        .B(GND), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[27] ), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/F_AWBURST_HTRANS0_net[1] ), .IPC());
    CFG4 #( .INIT(16'h0001) )  
        \reg_apb_wrp_0/reg16x8_0/temp_data_RNO[6]  (.A(
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_11[6]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_10[6]_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_9[6]_net_1 ), .D(
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_8[6]_net_1 ), .Y(
        \reg_apb_wrp_0/reg16x8_0/N_52_i_0 ));
    CFG4 #( .INIT(16'hB383) )  \CoreGPIO_0/CONFIG_reg_o_2_31_bm[6]  (
        .A(\CoreGPIO_0/CONFIG_reg_o_2_31_bm_RNO[6]_net_1 ), .B(
        \CoreGPIO_0/CONFIG_reg_o_2_31_bm_1[6] ), .C(
        \CoreAPB3_0_APBmslave3_PADDR[3] ), .D(
        \CoreGPIO_0/CONFIG_reg_o_2_31_bm_RNO_0[6]_net_1 ), .Y(
        \CoreGPIO_0/CONFIG_reg_o_2_31_bm[6]_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_144_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_26_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_144_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_144_rs_net_1 ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[4].APB_32.INTR_reg[4]  (.D(
        \CoreGPIO_0/INTR_reg_61[4] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB13_rgbr_net_1 ), .EN(VCC), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB3_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0.xhdl1.GEN_BITS[4].APB_32.INTR_reg[4] ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[30].REG_GEN.CONFIG_reg[30][6]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[6] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB12_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[30]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB2_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[30][6] ));
    CFG2 #( .INIT(4'h8) )  \CoreGPIO_0/PRDATA_iv_0_0_a2_0_0[0]  (.A(
        \CoreAPB3_0_APBmslave3_PADDR[5] ), .B(
        \CoreGPIO_0/GPOUT_reg[0] ), .Y(
        \CoreGPIO_0/PRDATA_iv_0_0_a2_0_0[0]_net_1 ));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_136_rs_RNID1TQ  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_10_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_136_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_1_rs[0] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_1_[0]_net_1 ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[17].REG_GEN.CONFIG_reg[17][7]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[7] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB14_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[17]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB4_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[17][7] ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_214  (.A(GND), 
        .B(GND), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/F_AWSIZE_HSIZE0_net[0] ), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/F_WID_HREADY01_net[2] ), .IPC());
    INV_BA AFLSDF_INV_110 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_54_net_1 ), .Y(
        AFLSDF_INV_110_net_1));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_189  (.A(VCC), 
        .B(VCC), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/I2C0_SDA_F2H_SCP_net ), .IPB(), .IPC(
        ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_185  (.A(VCC), 
        .B(VCC), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/MMUART0_RXD_F2H_SCP_net ), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/I2C0_SCL_F2H_SCP_net ), .IPC());
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_107_set_RNIQ3951  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_107_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_235_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_13_rs[3] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_13_[3]_net_1 ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[9].REG_GEN.CONFIG_reg[9][4]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[4] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB14_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[9]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB4_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[9][4] ));
    CFG4 #( .INIT(16'h7350) )  
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_5[6]  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_14_[6]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/mem_6_[6]_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/N_503 ), .D(
        \reg_apb_wrp_0/reg16x8_0/N_493 ), .Y(
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_5[6]_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_139_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_43_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_139_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_139_rs_net_1 ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[27].APB_32.INTR_reg[27]  (.D(
        \CoreGPIO_0/INTR_reg_360[27] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB10_rgbr_net_1 ), .EN(VCC), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB0_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/INTR_reg[27] ));
    INV_BA AFLSDF_INV_10 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_12_net_1 ), .Y(
        AFLSDF_INV_10_net_1));
    SLE \reg_apb_wrp_0/reg16x8_0/temp_data[7]  (.D(
        \reg_apb_wrp_0/reg16x8_0/N_86_i_0 ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB11_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/rd_enable_net_1 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB1_rgbl_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/temp_data[7]_net_1 ));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_221_rs_RNI43JO  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_5_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_221_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_8_rs[1] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_8_[1]_net_1 ));
    CFG4 #( .INIT(16'h1000) )  
        \reg_apb_wrp_0/reg16x8_0/WRITE_GEN.mem_3__2_i_a2[6]  (.A(
        \CoreAPB3_0_APBmslave3_PADDR[3] ), .B(
        \CoreAPB3_0_APBmslave3_PADDR[2] ), .C(
        \CoreAPB3_0_APBmslave3_PADDR[0] ), .D(
        \CoreAPB3_0_APBmslave3_PADDR[1] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/N_494 ));
    CFG3 #( .INIT(8'h4C) )  \FIC_MSS_0/MSS_ADLIB_INST_RNO_19  (.A(
        \CoreGPIO_0.xhdl1.GEN_BITS[0].APB_32.GPOUT_reg9 ), .B(
        \FIC_MSS_0/CoreAPB3_0_APBmslave5_PRDATA_m_0_1_0[5] ), .C(
        \CoreGPIO_0.xhdl1.GEN_BITS[5].APB_32.GPOUT_reg[5] ), .Y(
        \FIC_MSS_0/CoreAPB3_0_APBmslave5_PRDATA_m_0_1_1[5] ));
    CFG3 #( .INIT(8'hF2) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_166  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_4_[5]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_504 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_166_i ));
    CFG4 #( .INIT(16'h0F35) )  
        \CoreGPIO_0/CONFIG_reg_o_2_31_am_1_RNO_2[7]  (.A(
        \CoreGPIO_0/CONFIG_reg[0][7] ), .B(
        \CoreGPIO_0/CONFIG_reg[16][7] ), .C(
        \CoreAPB3_0_APBmslave3_PADDR[6] ), .D(
        \CoreAPB3_0_APBmslave3_PADDR[5] ), .Y(
        \CoreGPIO_0/CONFIG_reg_o_2_3_1[7] ));
    CFG4 #( .INIT(16'hAC0F) )  
        \CoreGPIO_0/CONFIG_reg_o_2_31_bm_RNO_0[2]  (.A(
        \CoreGPIO_0/CONFIG_reg[15][2] ), .B(
        \CoreGPIO_0/CONFIG_reg[31][2] ), .C(
        \CoreGPIO_0/CONFIG_reg_o_2_28_1_1[2] ), .D(
        \CoreAPB3_0_APBmslave3_PADDR[5] ), .Y(
        \CoreGPIO_0/CONFIG_reg_o_2_31_bm_RNO_0[2]_net_1 ));
    INV_BA AFLSDF_INV_112 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_17_net_1 ), .Y(
        AFLSDF_INV_112_net_1));
    CFG4 #( .INIT(16'hAA08) )  
        \CoreGPIO_0/xhdl1.GEN_BITS[5].APB_32.edge_pos_79_iv_i_0[5]  (
        .A(\CoreGPIO_0/CONFIG_reg[5][3] ), .B(\CoreGPIO_0/edge_pos[5] )
        , .C(\CoreAPB3_0_APBmslave3_PWDATA[5] ), .D(\CoreGPIO_0/N_406 )
        , .Y(\CoreGPIO_0/N_101 ));
    IO_DIFF \FIC_MSS_0/MDDR_CLK_PAD/U_ION  (.YIN(GND));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_7_[6]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[6] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB7_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_7__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_215_i ), .ADn(VCC), .SLn(
        VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_7_rs[6] ));
    CFG4 #( .INIT(16'h330A) )  
        \CoreGPIO_0/xhdl1.GEN_BITS[22].APB_32.INTR_reg_295_0[22]  (.A(
        \CoreGPIO_0/INTR_reg[22] ), .B(
        \CoreGPIO_0/INTR_reg_295_0_o2_1[22] ), .C(
        \CoreAPB3_0_APBmslave3_PWDATA[22] ), .D(\CoreGPIO_0/N_248 ), 
        .Y(\CoreGPIO_0/INTR_reg_295[22] ));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_14_[2]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[2] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB7_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_14__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_242_i ), .ADn(VCC), .SLn(
        VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_14_rs[2] ));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_158_rs_RNI2CFK  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_53_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_158_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_7_rs[4] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_7_[4]_net_1 ));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_8_set_RNI90TH  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_8_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_135_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_0_rs[7] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_0_[7]_net_1 ));
    CFG4 #( .INIT(16'h7530) )  
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_4[7]  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_12_[7]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/mem_4_[7]_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/N_504 ), .D(
        \reg_apb_wrp_0/reg16x8_0/N_495 ), .Y(
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_4[7]_net_1 ));
    IP_INTERFACE \FCCC_0/CCC_INST/IP_INTERFACE_17  (.A(VCC), .B(VCC), 
        .C(VCC), .IPA(), .IPB(\FCCC_0/CCC_INST/GPD3_ARST_N_net ), .IPC(
        \FCCC_0/CCC_INST/PADDR_net[7] ));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_233_rs_RNIKJMA1  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_105_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_233_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_13_rs[1] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_13_[1]_net_1 ));
    CFG3 #( .INIT(8'h7F) )  \FIC_MSS_0/MSS_ADLIB_INST_RNO_29  (.A(
        \CoreGPIO_0.xhdl1.GEN_BITS[5].gpin3[5] ), .B(
        \CoreGPIO_0.RDATA_32.un12_PRDATA_o ), .C(
        \CoreGPIO_0.xhdl1.GEN_BITS[5].REG_GEN.CONFIG_reg[5][1] ), .Y(
        \FIC_MSS_0/CoreAPB3_0_APBmslave5_PRDATA_m_0_1_0[5] ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_3_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB5_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_7__1_sqmuxa ), .ALn(
        AFLSDF_INV_53_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(GND)
        , .Q(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_3_set_net_1 ));
    CFG4 #( .INIT(16'hAC0F) )  
        \CoreGPIO_0/CONFIG_reg_o_2_31_bm_1_1_RNO[0]  (.A(
        \CoreGPIO_0/CONFIG_reg[13][0] ), .B(
        \CoreGPIO_0/CONFIG_reg[29][0] ), .C(
        \CoreGPIO_0/CONFIG_reg_o_2_21_1[0] ), .D(
        \CoreAPB3_0_APBmslave3_PADDR[5] ), .Y(
        \CoreGPIO_0/CONFIG_reg_o_2_31_bm_1_1_RNO[0]_net_1 ));
    INV_BA AFLSDF_INV_108 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_33_net_1 ), .Y(
        AFLSDF_INV_108_net_1));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_18  (.A(
        \FIC_MSS_0_FIC_0_APB_MASTER_PRDATA[23] ), .B(
        \FIC_MSS_0_FIC_0_APB_MASTER_PRDATA[30] ), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[23] ), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[30] ), .IPC());
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_54  (
        .A(\reg_apb_wrp_0/reg16x8_0/mem_7_[5]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_498 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_54_net_1 ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_32  (.A(GND), 
        .B(GND), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[8] ), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[15] ), .IPC());
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[4].gpin3[4]  (.D(
        \CoreGPIO_0/gpin2[4] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB13_rgbr_net_1 ), .EN(VCC), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB3_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0.xhdl1.GEN_BITS[4].gpin3[4] ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[29].APB_32.GPOUT_reg[29]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[29] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB11_rgbr_net_1 ), .EN(
        \CoreGPIO_0/GPOUT_reg_0_sqmuxa ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB1_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0.xhdl1.GEN_BITS[29].APB_32.GPOUT_reg[29] ));
    IOTRI_OB_EB \FIC_MSS_0/MDDR_CAS_N_PAD/U_IOOUT  (.D(VCC), .E(VCC), 
        .DOUT(), .EOUT(\FIC_MSS_0/MDDR_CAS_N_PAD/EOUT ));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_13_[1]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[1] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB9_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_13__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_233_i ), .ADn(VCC), .SLn(
        VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_13_rs[1] ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[7].REG_GEN.CONFIG_reg[7][7]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[7] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB10_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[7]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB0_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[7][7] ));
    sdf_IOPAD_BI \FIC_MSS_0/MDDR_DQ_12_PAD/U_IOPAD  (.PAD(MDDR_DQ[12]), 
        .D(\FIC_MSS_0/DRAM_DQ_OUT_net_0[12] ), .E(
        \FIC_MSS_0/DRAM_DQ_OE_net_0[12] ), .Y(
        \FIC_MSS_0/MDDR_DQ_12_PAD_Y ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_181_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_75_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_181_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_181_rs_net_1 ));
    CFG4 #( .INIT(16'hF2F3) )  
        \CoreGPIO_0/xhdl1.GEN_BITS[20].APB_32.INTR_reg_269_0_o2_1_0[20]  
        (.A(\CoreGPIO_0/CONFIG_reg[20][6] ), .B(
        \CoreGPIO_0/edge_neg[20] ), .C(
        \CoreGPIO_0/INTR_reg_269_0_o2_0[20] ), .D(
        \CoreGPIO_0/CONFIG_reg[20][5] ), .Y(
        \CoreGPIO_0/INTR_reg_269_0_o2_1[20] ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_25_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB10_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_5__1_sqmuxa ), .ALn(
        AFLSDF_INV_54_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(GND)
        , .Q(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_25_set_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_115_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB8_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_14__1_sqmuxa ), .ALn(
        AFLSDF_INV_55_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(GND)
        , .Q(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_115_set_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_13_[7]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[7] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB4_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_13__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_239_i ), .ADn(VCC), .SLn(
        VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_13_rs[7] ));
    CFG3 #( .INIT(8'h20) )  
        \CoreGPIO_0/xhdl1.GEN_BITS[16].APB_32.edge_both_RNO[16]  (.A(
        \CoreGPIO_0/CONFIG_reg[16][3] ), .B(
        \CoreAPB3_0_APBmslave3_PWDATA[16] ), .C(
        \CoreGPIO_0/edge_neg[16] ), .Y(\CoreGPIO_0/edge_neg_233[16] ));
    RCOSC_25_50MHZ #( .FREQUENCY(50.0) )  \OSC_0/I_RCOSC_25_50MHZ  (
        .CLKOUT(OSC_0_RCOSC_25_50MHZ_CCC_OUT_RCOSC_25_50MHZ_CCC));
    CFG3 #( .INIT(8'h7F) )  \FIC_MSS_0/MSS_ADLIB_INST_RNO_17  (.A(
        \CoreGPIO_0.xhdl1.GEN_BITS[2].gpin3[2] ), .B(
        \CoreGPIO_0.RDATA_32.un12_PRDATA_o ), .C(
        \CoreGPIO_0.xhdl1.GEN_BITS[2].REG_GEN.CONFIG_reg[2][1] ), .Y(
        \FIC_MSS_0/CoreAPB3_0_APBmslave5_PRDATA_m_0_1[2] ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_108  (.A(VCC), 
        .B(VCC), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/FAB_XDATAIN_net[0] ), .IPB(), .IPC());
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[28].APB_32.edge_both[28]  (.D(
        \CoreGPIO_0/N_87_i_0 ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB13_rgbr_net_1 ), .EN(
        \CoreGPIO_0/N_163 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB3_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/edge_pos[28] ));
    CFG2 #( .INIT(4'h7) )  \CoreGPIO_0/edge_both_2_sqmuxa_31_i  (.A(
        \CoreGPIO_0/N_248 ), .B(\CoreGPIO_0/CONFIG_reg[24][3] ), .Y(
        \CoreGPIO_0/N_155 ));
    CFG4 #( .INIT(16'h7350) )  
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_3[0]  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_11_[0]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/mem_3_[0]_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/N_505 ), .D(
        \reg_apb_wrp_0/reg16x8_0/N_494 ), .Y(
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_3[0]_net_1 ));
    CFG4 #( .INIT(16'h5410) )  \CoreGPIO_0/PRDATA_iv_0_0_0_1[0]  (.A(
        \CoreAPB3_0_APBmslave3_PADDR[7] ), .B(
        \CoreAPB3_0_APBmslave3_PADDR[2] ), .C(
        \CoreGPIO_0/CONFIG_reg_o_2_31_am[0]_net_1 ), .D(
        \CoreGPIO_0/CONFIG_reg_o_2_31_bm[0]_net_1 ), .Y(
        \CoreGPIO_0.PRDATA_iv_0_0_0_0[0] ));
    CFG4 #( .INIT(16'hAA08) )  
        \CoreGPIO_0/xhdl1.GEN_BITS[4].APB_32.edge_pos_65_iv_i_0[4]  (
        .A(\CoreGPIO_0/CONFIG_reg[4][3] ), .B(\CoreGPIO_0/edge_pos[4] )
        , .C(\CoreAPB3_0_APBmslave3_PWDATA[4] ), .D(\CoreGPIO_0/N_398 )
        , .Y(\CoreGPIO_0/N_103 ));
    IOTRI_OB_EB \FIC_MSS_0/MDDR_ADDR_1_PAD/U_IOOUT  (.D(VCC), .E(VCC), 
        .DOUT(), .EOUT(\FIC_MSS_0/MDDR_ADDR_1_PAD/EOUT ));
    RGB \FCCC_0/GL1_INST/U0_RGB1_RGB15  (.An(
        \FCCC_0/GL1_INST/U0_YNn_GSouth ), .ENn(GND), .YL(
        \FCCC_0/GL1_INST/U0_RGB1_RGB15_rgbl_net_1 ), .YR(
        \FCCC_0/GL1_INST/U0_RGB1_RGB15_rgbr_net_1 ));
    CFG4 #( .INIT(16'h2000) )  
        \CoreGPIO_0/xhdl1.GEN_BITS[22].REG_GEN.CONFIG_reg[22]2_0_a4_0_a2  
        (.A(\CoreAPB3_0_APBmslave3_PADDR[3] ), .B(
        \CoreAPB3_0_APBmslave3_PADDR[2] ), .C(\CoreGPIO_0/N_598 ), .D(
        \CoreGPIO_0/N_603 ), .Y(\CoreGPIO_0/CONFIG_reg[22]2 ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_182_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_46_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_182_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_182_rs_net_1 ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[1].REG_GEN.CONFIG_reg[1][1]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[1] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB16_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[1]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB6_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0.xhdl1.GEN_BITS[1].REG_GEN.CONFIG_reg[1][1] ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_199_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_101_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_199_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_199_rs_net_1 ));
    INV_BA AFLSDF_INV_95 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_106_net_1 ), .Y(
        AFLSDF_INV_95_net_1));
    sdf_IOPAD_IN \FIC_MSS_0/MDDR_DQS_TMATCH_0_IN_PAD/U_IOPAD  (.PAD(
        MDDR_DQS_TMATCH_0_IN), .Y(
        \FIC_MSS_0/MDDR_DQS_TMATCH_0_IN_PAD_Y ));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_6_[4]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[4] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB7_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_6__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_196_i ), .ADn(VCC), .SLn(
        VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_6_rs[4] ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_29  (.A(GND), 
        .B(GND), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[5] ), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[12] ), .IPC());
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_116  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_14_[4]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_503 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_116_net_1 ));
    RGB \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB2  (.An(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_YNn_GSouth ), .ENn(GND), .YL(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB2_rgbl_net_1 ), .YR(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB2_rgbr_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_61_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB5_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_15__1_sqmuxa ), .ALn(
        AFLSDF_INV_56_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(GND)
        , .Q(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_61_set_net_1 ));
    CFG4 #( .INIT(16'hA9FF) )  
        \CoreGPIO_0/xhdl1.GEN_BITS[10].APB_32.INTR_reg_139_0_o2_0_0[10]  
        (.A(\CoreGPIO_0/CONFIG_reg[10][7] ), .B(
        \CoreGPIO_0/CONFIG_reg[10][6] ), .C(
        \CoreGPIO_0/CONFIG_reg[10][5] ), .D(
        \CoreGPIO_0/CONFIG_reg[10][3] ), .Y(
        \CoreGPIO_0/INTR_reg_139_0_o2_0[10] ));
    CFG3 #( .INIT(8'h80) )  \FIC_MSS_0/MSS_ADLIB_INST_RNO_27  (.A(
        \CoreGPIO_0.xhdl1.GEN_BITS[3].gpin3[3] ), .B(
        CoreAPB3_0_APBmslave5_PSELx), .C(
        \CoreGPIO_0.xhdl1.GEN_BITS[3].REG_GEN.CONFIG_reg[3][1] ), .Y(
        \FIC_MSS_0/CoreAPB3_0_APBmslave5_PRDATA_m_c_c_1[3] ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[2].gpin1[2]  (.D(\GPIO_IN_c[2] ), 
        .CLK(\FCCC_0/GL1_INST/U0_RGB1_RGB17_rgbr_net_1 ), .EN(VCC), 
        .ALn(\MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB7_rgbr_net_1 ), 
        .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/gpin1[2] ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[19].APB_32.INTR_reg[19]  (.D(
        \CoreGPIO_0/INTR_reg_256[19] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB10_rgbr_net_1 ), .EN(VCC), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB0_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/INTR_reg[19] ));
    INV_BA AFLSDF_INV_29 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_125_net_1 ), .Y(
        AFLSDF_INV_29_net_1));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/mem_2__RNI4TJP[7]  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_120_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_151_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_2_rs[7] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_2_[7]_net_1 ));
    CFG4 #( .INIT(16'hFFFE) )  
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_13[4]  (.A(
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_7[4]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_5[4]_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_6[4]_net_1 ), .D(
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_4[4]_net_1 ), .Y(
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_13[4]_net_1 ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[21].REG_GEN.CONFIG_reg[21][6]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[6] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB13_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[21]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB3_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[21][6] ));
    INV_BA AFLSDF_INV_89 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_96_net_1 ), .Y(
        AFLSDF_INV_89_net_1));
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_60  (
        .A(\reg_apb_wrp_0/reg16x8_0/mem_15_[7]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_497 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_60_net_1 ));
    IOENFF_BYPASS \GPIO_OUT_obuf[6]/U0/U_IOENFF  (.A(
        \GPIO_OUT_obuf[6]/U0/EOUT1 ), .Y(\GPIO_OUT_obuf[6]/U0/EOUT ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_158_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_53_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_158_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_158_rs_net_1 ));
    CFG4 #( .INIT(16'hB383) )  \CoreGPIO_0/CONFIG_reg_o_2_31_am[7]  (
        .A(\CoreGPIO_0/CONFIG_reg_o_2_31_am_RNO[7]_net_1 ), .B(
        \CoreGPIO_0/CONFIG_reg_o_2_31_am_1[7] ), .C(
        \CoreAPB3_0_APBmslave3_PADDR[3] ), .D(
        \CoreGPIO_0/CONFIG_reg_o_2_31_am_RNO_0[7]_net_1 ), .Y(
        \CoreGPIO_0/CONFIG_reg_o_2_31_am[7]_net_1 ));
    INV_BA AFLSDF_INV_27 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_18_net_1 ), .Y(
        AFLSDF_INV_27_net_1));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_121  (.A(VCC), 
        .B(VCC), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/FAB_AVALID_net ), .IPB(), .IPC());
    CFG2 #( .INIT(4'h7) )  \CoreGPIO_0/edge_both_2_sqmuxa_7_i  (.A(
        \CoreGPIO_0/N_248 ), .B(\CoreGPIO_0/CONFIG_reg[21][3] ), .Y(
        \CoreGPIO_0/N_198 ));
    INV_BA AFLSDF_INV_87 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_63_net_1 ), .Y(
        AFLSDF_INV_87_net_1));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_0_[0]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[0] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB2_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_0__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_131_i ), .ADn(VCC), .SLn(
        VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_0_rs[0] ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_150  (.A(VCC), 
        .B(VCC), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/MGPIO2A_F2H_GPIN_net ), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/SPI0_SDI_F2H_SCP_net ), .IPC());
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_20  (
        .A(\reg_apb_wrp_0/reg16x8_0/mem_12_[4]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_495 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_20_net_1 ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_256  (.A(VCC), 
        .B(VCC), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[4] ), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[16] ), .IPC());
    CFG4 #( .INIT(16'hEFEE) )  
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_8[3]  (.A(
        \reg_apb_wrp_0/reg16x8_0/N_406 ), .B(
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_1[3]_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_5_[3]_net_1 ), .D(
        \reg_apb_wrp_0/reg16x8_0/N_490 ), .Y(
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_8[3]_net_1 ));
    CFG4 #( .INIT(16'hAC0F) )  
        \CoreGPIO_0/CONFIG_reg_o_2_31_am_1_1_RNO[1]  (.A(
        \CoreGPIO_0/CONFIG_reg[12][1] ), .B(
        \CoreGPIO_0/CONFIG_reg[28][1] ), .C(
        \CoreGPIO_0/CONFIG_reg_o_2_6_1[1] ), .D(
        \CoreAPB3_0_APBmslave3_PADDR[5] ), .Y(
        \CoreGPIO_0/CONFIG_reg_o_2_31_am_1_1_RNO[1]_net_1 ));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_54_set_RNISMNC  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_54_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_213_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_7_rs[5] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_7_[5]_net_1 ));
    INV_BA AFLSDF_INV_1 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_121_net_1 ), .Y(
        AFLSDF_INV_1_net_1));
    IOOUTFF_BYPASS \GPIO_OUT_obuf[1]/U0/U_IOOUTFF  (.A(
        \GPIO_OUT_obuf[1]/U0/DOUT1 ), .Y(\GPIO_OUT_obuf[1]/U0/DOUT ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[26].APB_32.edge_both[26]  (.D(
        \CoreGPIO_0/N_106_i_0 ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB17_rgbr_net_1 ), .EN(
        \CoreGPIO_0/N_159 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB7_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/edge_pos[26] ));
    CFG2 #( .INIT(4'h4) )  
        \CoreGPIO_0/xhdl1.GEN_BITS[4].REG_GEN.CONFIG_reg[4]2_0_a4_0_a2_0  
        (.A(\CoreAPB3_0_APBmslave3_PADDR[5] ), .B(
        \CoreAPB3_0_APBmslave3_PADDR[4] ), .Y(\CoreGPIO_0/N_603 ));
    CFG4 #( .INIT(16'hF2F3) )  
        \CoreGPIO_0/xhdl1.GEN_BITS[19].APB_32.INTR_reg_256_0_o2_1_0[19]  
        (.A(\CoreGPIO_0/CONFIG_reg[19][6] ), .B(
        \CoreGPIO_0/edge_neg[19] ), .C(
        \CoreGPIO_0/INTR_reg_256_0_o2_0[19] ), .D(
        \CoreGPIO_0/CONFIG_reg[19][5] ), .Y(
        \CoreGPIO_0/INTR_reg_256_0_o2_1[19] ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_197  (.A(VCC), 
        .B(VCC), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[1] ), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[13] ), .IPC());
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_104  (.A(VCC), 
        .B(VCC), .C(VCC), .IPA(\FIC_MSS_0/MSS_ADLIB_INST/RCGF_net[4] ), 
        .IPB(\FIC_MSS_0/MSS_ADLIB_INST/FAB_LINESTATE_net[0] ), .IPC());
    INV_BA AFLSDF_INV_127 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_68_net_1 ), .Y(
        AFLSDF_INV_127_net_1));
    INV_BA AFLSDF_INV_58 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_59_net_1 ), .Y(
        AFLSDF_INV_58_net_1));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[28].APB_32.GPOUT_reg[28]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[28] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB13_rgbr_net_1 ), .EN(
        \CoreGPIO_0/GPOUT_reg_0_sqmuxa ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB3_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0.xhdl1.GEN_BITS[28].APB_32.GPOUT_reg[28] ));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_15_[3]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[3] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB4_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_15__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_251_i ), .ADn(VCC), .SLn(
        VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_15_rs[3] ));
    CFG3 #( .INIT(8'hF2) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_243  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_14_[3]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_503 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_243_i ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[14].REG_GEN.CONFIG_reg[14][4]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[4] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB14_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[14]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB4_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[14][4] ));
    CFG4 #( .INIT(16'h4657) )  
        \CoreGPIO_0/CONFIG_reg_o_2_31_bm_1_1[7]  (.A(
        \CoreAPB3_0_APBmslave3_PADDR[4] ), .B(
        \CoreAPB3_0_APBmslave3_PADDR[3] ), .C(
        \CoreGPIO_0/CONFIG_reg_o_2_31_bm_1_1_RNO[7]_net_1 ), .D(
        \CoreGPIO_0/CONFIG_reg_o_2_31_bm_1_RNO_0[7]_net_1 ), .Y(
        \CoreGPIO_0/CONFIG_reg_o_2_31_bm_1[7] ));
    CFG4 #( .INIT(16'h7350) )  
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_5[2]  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_14_[2]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/mem_6_[2]_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/N_503 ), .D(
        \reg_apb_wrp_0/reg16x8_0/N_493 ), .Y(
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_5[2]_net_1 ));
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_13  (
        .A(\reg_apb_wrp_0/reg16x8_0/mem_5_[0]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_490 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_13_net_1 ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[18].REG_GEN.CONFIG_reg[18][6]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[6] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB17_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[18]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB7_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[18][6] ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[0].REG_GEN.CONFIG_reg[0][0]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[0] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB11_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[0]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB1_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[0][0] ));
    INV_BA AFLSDF_INV_119 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_10_net_1 ), .Y(
        AFLSDF_INV_119_net_1));
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_52  (
        .A(\reg_apb_wrp_0/reg16x8_0/mem_3_[5]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_494 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_52_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/data_out[6]  (.D(
        \reg_apb_wrp_0/reg16x8_0/temp_data[6]_net_1 ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB12_rgbr_net_1 ), .EN(VCC), .ALn(
        VCC), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreAPB3_0_APBmslave3_PRDATA[6] ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[30].REG_GEN.CONFIG_reg[30][5]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[5] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB12_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[30]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB2_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[30][5] ));
    CFG4 #( .INIT(16'hF2F3) )  
        \CoreGPIO_0/xhdl1.GEN_BITS[11].APB_32.INTR_reg_152_0_o2_1_0[11]  
        (.A(\CoreGPIO_0/CONFIG_reg[11][6] ), .B(
        \CoreGPIO_0/edge_neg[11] ), .C(
        \CoreGPIO_0/INTR_reg_152_0_o2_0[11] ), .D(
        \CoreGPIO_0/CONFIG_reg[11][5] ), .Y(
        \CoreGPIO_0/INTR_reg_152_0_o2_1[11] ));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_13_[6]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[6] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB11_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_13__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_238_i ), .ADn(VCC), .SLn(
        VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_13_rs[6] ));
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_88  (
        .A(\reg_apb_wrp_0/reg16x8_0/mem_11_[0]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_505 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_88_net_1 ));
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_46  (
        .A(\reg_apb_wrp_0/reg16x8_0/mem_5_[5]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_490 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_46_net_1 ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[19].REG_GEN.CONFIG_reg[19][1]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[1] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB10_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[19]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB0_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[19][1] ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[1].APB_32.edge_both[1]  (.D(
        \CoreGPIO_0/N_95 ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB16_rgbr_net_1 ), .EN(
        \CoreGPIO_0/N_82 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB6_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/edge_both[1] ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_76_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB13_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_9__1_sqmuxa ), .ALn(
        AFLSDF_INV_57_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(GND)
        , .Q(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_76_set_net_1 ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_230  (.A(VCC), 
        .B(VCC), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[28] ), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[40] ), .IPC());
    sdf_IOPAD_TRI \FIC_MSS_0/MDDR_ADDR_9_PAD/U_IOPAD  (.PAD(
        MDDR_ADDR[9]), .D(\FIC_MSS_0/DRAM_ADDR_net_0[9] ), .E(
        \FIC_MSS_0/MDDR_ADDR_9_PAD/EOUT ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_203  (.A(VCC), 
        .B(VCC), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[7] ), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[19] ), .IPC());
    RGB \FCCC_0/GL1_INST/U0_RGB1_RGB7  (.An(\FCCC_0/GL1_INST/U0_YNn ), 
        .ENn(GND), .YL(\FCCC_0/GL1_INST/U0_RGB1_RGB7_rgbl_net_1 ), .YR(
        \FCCC_0/GL1_INST/U0_RGB1_RGB7_rgbr_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_59_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB5_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_15__1_sqmuxa ), .ALn(
        AFLSDF_INV_58_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(GND)
        , .Q(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_59_set_net_1 ));
    IOENFF_BYPASS \GPIO_OUT_obuf[3]/U0/U_IOENFF  (.A(
        \GPIO_OUT_obuf[3]/U0/EOUT1 ), .Y(\GPIO_OUT_obuf[3]/U0/EOUT ));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_212_rs_RNI5DKN  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_91_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_212_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_11_rs[3] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_11_[3]_net_1 ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_237  (.A(VCC), 
        .B(VCC), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[35] ), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[47] ), .IPC());
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[17].REG_GEN.CONFIG_reg[17][0]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[0] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB16_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[17]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB6_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[17][0] ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[27].REG_GEN.CONFIG_reg[27][2]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[2] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB10_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[27]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB0_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[27][2] ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[22].REG_GEN.CONFIG_reg[22][3]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[3] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB12_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[22]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB2_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[22][3] ));
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_98  (
        .A(\reg_apb_wrp_0/reg16x8_0/mem_10_[1]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_491 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_98_net_1 ));
    INV_BA AFLSDF_INV_40 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_91_net_1 ), .Y(
        AFLSDF_INV_40_net_1));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_1_[6]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[6] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB16_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_1__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_142_i ), .ADn(VCC), .SLn(
        VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_1_rs[6] ));
    CFG2 #( .INIT(4'h4) )  \CoreGPIO_0/PRDATA_0_iv_0_a2_0[16]  (.A(
        \CoreGPIO_0.N_247 ), .B(\CoreGPIO_0/INTR_reg[16] ), .Y(
        \CoreGPIO_0.N_554 ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_35_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB8_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_6__1_sqmuxa ), .ALn(
        AFLSDF_INV_59_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(GND)
        , .Q(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_35_set_net_1 ));
    CFG4 #( .INIT(16'h330A) )  
        \CoreGPIO_0/xhdl1.GEN_BITS[18].APB_32.INTR_reg_243_0[18]  (.A(
        \CoreGPIO_0.xhdl1.GEN_BITS[18].APB_32.INTR_reg[18] ), .B(
        \CoreGPIO_0/INTR_reg_243_0_o2_1[18] ), .C(
        \CoreAPB3_0_APBmslave3_PWDATA[18] ), .D(\CoreGPIO_0/N_248 ), 
        .Y(\CoreGPIO_0/INTR_reg_243[18] ));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_7_[3]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[3] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB3_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_7__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_210_i ), .ADn(VCC), .SLn(
        VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_7_rs[3] ));
    CFG3 #( .INIT(8'h04) )  
        \CoreGPIO_0/xhdl1.GEN_BITS[6].APB_32.INTR_reg_87_0_0_RNO_0[6]  
        (.A(\CoreGPIO_0/CONFIG_reg[6][5] ), .B(
        \CoreGPIO_0/edge_both[6] ), .C(\CoreGPIO_0/CONFIG_reg[6][6] ), 
        .Y(\CoreGPIO_0/INTR_reg_87_0_0_55_tz_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_141_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_47_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_141_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_141_rs_net_1 ));
    CFG2 #( .INIT(4'h2) )  \CoreGPIO_0/edge_pos_2_sqmuxa_3_i_a2  (.A(
        \CoreGPIO_0/gpin2[5] ), .B(
        \CoreGPIO_0.xhdl1.GEN_BITS[5].gpin3[5] ), .Y(
        \CoreGPIO_0/N_406 ));
    CFG4 #( .INIT(16'hF2F3) )  
        \CoreGPIO_0/xhdl1.GEN_BITS[8].APB_32.INTR_reg_113_0_o2_1_0[8]  
        (.A(\CoreGPIO_0/CONFIG_reg[8][6] ), .B(
        \CoreGPIO_0/edge_pos[8] ), .C(
        \CoreGPIO_0/INTR_reg_113_0_o2_0[8] ), .D(
        \CoreGPIO_0/CONFIG_reg[8][5] ), .Y(
        \CoreGPIO_0/INTR_reg_113_0_o2_1[8] ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_46_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB8_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_5__1_sqmuxa ), .ALn(
        AFLSDF_INV_60_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(GND)
        , .Q(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_46_set_net_1 ));
    CFG3 #( .INIT(8'hF2) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_196  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_6_[4]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_493 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_196_i ));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_69_set_RNIDLDH  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_69_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_169_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_8_rs[5] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_8_[5]_net_1 ));
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_8  (
        .A(\reg_apb_wrp_0/reg16x8_0/mem_0_[7]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_496 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_8_net_1 ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_6  (.A(
        \FIC_MSS_0/FIC_MSS_0_FIC_0_APB_MASTER_PRDATA[4] ), .B(
        \FIC_MSS_0_FIC_0_APB_MASTER_PRDATA[11] ), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[4] ), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[11] ), .IPC());
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_142_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_45_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_142_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_142_rs_net_1 ));
    sdf_IOPAD_IN \GPIO_IN_ibuf[4]/U0/U_IOPAD  (.PAD(GPIO_IN[4]), .Y(
        \GPIO_IN_ibuf[4]/U0/YIN1 ));
    CFG4 #( .INIT(16'h4657) )  
        \CoreGPIO_0/CONFIG_reg_o_2_31_am_1_1[5]  (.A(
        \CoreAPB3_0_APBmslave3_PADDR[4] ), .B(
        \CoreAPB3_0_APBmslave3_PADDR[3] ), .C(
        \CoreGPIO_0/CONFIG_reg_o_2_31_am_1_1_RNO[5]_net_1 ), .D(
        \CoreGPIO_0/CONFIG_reg_o_2_31_am_1_RNO_0[5]_net_1 ), .Y(
        \CoreGPIO_0/CONFIG_reg_o_2_31_am_1[5] ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[29].REG_GEN.CONFIG_reg[29][0]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[0] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB14_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[29]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB4_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[29][0] ));
    CFG4 #( .INIT(16'h330A) )  
        \CoreGPIO_0/xhdl1.GEN_BITS[20].APB_32.INTR_reg_269_0[20]  (.A(
        \CoreGPIO_0/INTR_reg[20] ), .B(
        \CoreGPIO_0/INTR_reg_269_0_o2_1[20] ), .C(
        \CoreAPB3_0_APBmslave3_PWDATA[20] ), .D(\CoreGPIO_0/N_248 ), 
        .Y(\CoreGPIO_0/INTR_reg_269[20] ));
    CFG3 #( .INIT(8'hF2) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_219  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_8_[0]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_499 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_219_i ));
    CFG4 #( .INIT(16'hAC0F) )  
        \CoreGPIO_0/CONFIG_reg_o_2_31_bm_1_1_RNO[4]  (.A(
        \CoreGPIO_0/CONFIG_reg[13][4] ), .B(
        \CoreGPIO_0/CONFIG_reg[29][4] ), .C(
        \CoreGPIO_0/CONFIG_reg_o_2_21_1[4] ), .D(
        \CoreAPB3_0_APBmslave3_PADDR[5] ), .Y(
        \CoreGPIO_0/CONFIG_reg_o_2_31_bm_1_1_RNO[4]_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_6_[2]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[2] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB12_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_6__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_192_i ), .ADn(VCC), .SLn(
        VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_6_rs[2] ));
    INV_BA AFLSDF_INV_91 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_78_net_1 ), .Y(
        AFLSDF_INV_91_net_1));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[10].REG_GEN.CONFIG_reg[10][4]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[4] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB17_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[10]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB7_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[10][4] ));
    CFG4 #( .INIT(16'h4000) )  
        \CoreGPIO_0/xhdl1.GEN_BITS[9].REG_GEN.CONFIG_reg[9]2_0_a4_0_a2  
        (.A(\CoreAPB3_0_APBmslave3_PADDR[3] ), .B(
        \CoreAPB3_0_APBmslave3_PADDR[2] ), .C(\CoreGPIO_0/N_604 ), .D(
        \CoreGPIO_0/N_610 ), .Y(\CoreGPIO_0/CONFIG_reg[9]2 ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[12].REG_GEN.CONFIG_reg[12][7]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[7] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB12_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[12]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB2_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[12][7] ));
    CFG4 #( .INIT(16'h0F35) )  
        \CoreGPIO_0/CONFIG_reg_o_2_31_am_RNO_1[0]  (.A(
        \CoreGPIO_0/CONFIG_reg[2][0] ), .B(
        \CoreGPIO_0/CONFIG_reg[18][0] ), .C(
        \CoreAPB3_0_APBmslave3_PADDR[6] ), .D(
        \CoreAPB3_0_APBmslave3_PADDR[5] ), .Y(
        \CoreGPIO_0/CONFIG_reg_o_2_10_1_1[0] ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_135_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_8_net_1 ), .EN(VCC), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_135_i ), .ADn(VCC), .SLn(
        VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_135_rs_net_1 ));
    IOINFF_BYPASS \GPIO_IN_ibuf[6]/U0/U_IOINFF  (.A(
        \GPIO_IN_ibuf[6]/U0/YIN1 ), .Y(\GPIO_IN_ibuf[6]/U0/YIN ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_254  (.A(VCC), 
        .B(VCC), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[2] ), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[14] ), .IPC());
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[4].gpin2[4]  (.D(
        \CoreGPIO_0/gpin1[4] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB12_rgbr_net_1 ), .EN(VCC), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB2_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(\CoreGPIO_0/gpin2[4] )
        );
    CFG4 #( .INIT(16'hAC0F) )  
        \CoreGPIO_0/CONFIG_reg_o_2_31_am_RNO_0[4]  (.A(
        \CoreGPIO_0/CONFIG_reg[14][4] ), .B(
        \CoreGPIO_0/CONFIG_reg[30][4] ), .C(
        \CoreGPIO_0/CONFIG_reg_o_2_13_1_1[4] ), .D(
        \CoreAPB3_0_APBmslave3_PADDR[5] ), .Y(
        \CoreGPIO_0/CONFIG_reg_o_2_31_am_RNO_0[4]_net_1 ));
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_41  (
        .A(\reg_apb_wrp_0/reg16x8_0/mem_1_[4]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_502 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_41_net_1 ));
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_9  (
        .A(\reg_apb_wrp_0/reg16x8_0/mem_4_[6]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_504 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_9_net_1 ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[24].APB_32.INTR_reg[24]  (.D(
        \CoreGPIO_0/INTR_reg_321[24] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB10_rgbr_net_1 ), .EN(VCC), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB0_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/INTR_reg[24] ));
    CFG4 #( .INIT(16'hAC0F) )  
        \CoreGPIO_0/CONFIG_reg_o_2_31_am_1_RNO_0[2]  (.A(
        \CoreGPIO_0/CONFIG_reg[8][2] ), .B(
        \CoreGPIO_0/CONFIG_reg[24][2] ), .C(
        \CoreGPIO_0/CONFIG_reg_o_2_3_1[2] ), .D(
        \CoreAPB3_0_APBmslave3_PADDR[5] ), .Y(
        \CoreGPIO_0/CONFIG_reg_o_2_31_am_1_RNO_0[2]_net_1 ));
    INV_BA AFLSDF_INV_69 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_90_net_1 ), .Y(
        AFLSDF_INV_69_net_1));
    CFG3 #( .INIT(8'h20) )  
        \CoreGPIO_0/xhdl1.GEN_BITS[23].APB_32.edge_both_RNO[23]  (.A(
        \CoreGPIO_0/CONFIG_reg[23][3] ), .B(
        \CoreAPB3_0_APBmslave3_PWDATA[23] ), .C(
        \CoreGPIO_0/edge_neg[23] ), .Y(\CoreGPIO_0/N_96_i_0 ));
    CFG4 #( .INIT(16'h0F35) )  
        \CoreGPIO_0/CONFIG_reg_o_2_31_am_1_RNO_1[0]  (.A(
        \CoreGPIO_0/CONFIG_reg[4][0] ), .B(
        \CoreGPIO_0/CONFIG_reg[20][0] ), .C(
        \CoreAPB3_0_APBmslave3_PADDR[6] ), .D(
        \CoreAPB3_0_APBmslave3_PADDR[5] ), .Y(
        \CoreGPIO_0/CONFIG_reg_o_2_6_1[0] ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[3].REG_GEN.CONFIG_reg[3][1]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[1] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB10_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[3]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB0_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0.xhdl1.GEN_BITS[3].REG_GEN.CONFIG_reg[3][1] ));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_15_[5]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[5] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB7_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_15__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_254_i ), .ADn(VCC), .SLn(
        VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_15_rs[5] ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_97_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB1_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_10__1_sqmuxa ), .ALn(
        AFLSDF_INV_61_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(GND)
        , .Q(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_97_set_net_1 ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[18].APB_32.INTR_reg[18]  (.D(
        \CoreGPIO_0/INTR_reg_243[18] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB16_rgbr_net_1 ), .EN(VCC), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB6_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0.xhdl1.GEN_BITS[18].APB_32.INTR_reg[18] ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_176  (.A(VCC), 
        .B(VCC), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/MGPIO26B_F2H_GPIN_net ), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/MMUART0_CTS_F2H_SCP_net ), .IPC());
    CFG4 #( .INIT(16'h0F35) )  
        \CoreGPIO_0/CONFIG_reg_o_2_31_bm_RNO_2[1]  (.A(
        \CoreGPIO_0/CONFIG_reg[7][1] ), .B(
        \CoreGPIO_0/CONFIG_reg[23][1] ), .C(
        \CoreAPB3_0_APBmslave3_PADDR[6] ), .D(
        \CoreAPB3_0_APBmslave3_PADDR[5] ), .Y(
        \CoreGPIO_0/CONFIG_reg_o_2_28_1_1[1] ));
    CFG4 #( .INIT(16'h0F35) )  
        \CoreGPIO_0/CONFIG_reg_o_2_31_bm_RNO_1[3]  (.A(
        \CoreGPIO_0/CONFIG_reg[3][3] ), .B(
        \CoreGPIO_0/CONFIG_reg[19][3] ), .C(
        \CoreAPB3_0_APBmslave3_PADDR[6] ), .D(
        \CoreAPB3_0_APBmslave3_PADDR[5] ), .Y(
        \CoreGPIO_0/CONFIG_reg_o_2_25_1_1[3] ));
    CFG4 #( .INIT(16'hCC0A) )  
        \CoreGPIO_0/xhdl1.GEN_BITS[6].APB_32.INTR_reg_87_0_0[6]  (.A(
        \CoreGPIO_0.xhdl1.GEN_BITS[6].APB_32.INTR_reg[6] ), .B(
        \CoreGPIO_0/N_1580_tz ), .C(\CoreAPB3_0_APBmslave3_PWDATA[6] ), 
        .D(\CoreGPIO_0/N_248 ), .Y(\CoreGPIO_0/INTR_reg_87[6] ));
    CFG4 #( .INIT(16'hAC0F) )  
        \CoreGPIO_0/CONFIG_reg_o_2_31_am_RNO[0]  (.A(
        \CoreGPIO_0/CONFIG_reg[10][0] ), .B(
        \CoreGPIO_0/CONFIG_reg[26][0] ), .C(
        \CoreGPIO_0/CONFIG_reg_o_2_10_1_1[0] ), .D(
        \CoreAPB3_0_APBmslave3_PADDR[5] ), .Y(
        \CoreGPIO_0/CONFIG_reg_o_2_31_am_RNO[0]_net_1 ));
    INV_BA AFLSDF_INV_67 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_72_net_1 ), .Y(
        AFLSDF_INV_67_net_1));
    IP_INTERFACE \FCCC_0/CCC_INST/IP_INTERFACE_6  (.A(VCC), .B(VCC), 
        .C(VCC), .IPA(\FCCC_0/CCC_INST/CLK2_net ), .IPB(), .IPC(
        \FCCC_0/CCC_INST/PWDATA_net[4] ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[18].REG_GEN.CONFIG_reg[18][3]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[3] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB17_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[18]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB7_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[18][3] ));
    CFG3 #( .INIT(8'hF2) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_223  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_8_[2]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_499 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_223_i ));
    SLE \reg_apb_wrp_0/reg16x8_0/temp_data[5]  (.D(
        \reg_apb_wrp_0/reg16x8_0/N_25_i_0 ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB11_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/rd_enable_net_1 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB1_rgbl_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/temp_data[5]_net_1 ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_77  (.A(VCC), 
        .B(VCC), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[11] ), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[18] ), .IPC());
    CFG4 #( .INIT(16'h7530) )  
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_7[1]  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_10_[1]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/mem_2_[1]_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/N_501 ), .D(
        \reg_apb_wrp_0/reg16x8_0/N_491 ), .Y(
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_7[1]_net_1 ));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/mem_2__RNIK0IK[0]  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_26_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_144_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_2_rs[0] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_2_[0]_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_15_[4]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[4] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB6_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_15__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_253_i ), .ADn(VCC), .SLn(
        VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_15_rs[4] ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_92  (.A(VCC), 
        .B(VCC), .C(VCC), .IPA(\FIC_MSS_0/MSS_ADLIB_INST/RX_CLKPF_net )
        , .IPB(\FIC_MSS_0/MSS_ADLIB_INST/RX_ERRF_net ), .IPC());
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_86  (.A(VCC), 
        .B(VCC), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[27] ), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/RXDF_net[2] ), .IPC());
    CFG4 #( .INIT(16'hAA08) )  
        \CoreGPIO_0/xhdl1.GEN_BITS[4].APB_32.edge_neg_65_iv_i_0[4]  (
        .A(\CoreGPIO_0/CONFIG_reg[4][3] ), .B(\CoreGPIO_0/edge_neg[4] )
        , .C(\CoreAPB3_0_APBmslave3_PWDATA[4] ), .D(\CoreGPIO_0/N_397 )
        , .Y(\CoreGPIO_0/N_117 ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_88_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB17_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_11__1_sqmuxa ), .ALn(
        AFLSDF_INV_62_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(GND)
        , .Q(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_88_set_net_1 ));
    sdf_IOPAD_TRI \FIC_MSS_0/MDDR_ADDR_6_PAD/U_IOPAD  (.PAD(
        MDDR_ADDR[6]), .D(\FIC_MSS_0/DRAM_ADDR_net_0[6] ), .E(
        \FIC_MSS_0/MDDR_ADDR_6_PAD/EOUT ));
    CFG4 #( .INIT(16'hA9FF) )  
        \CoreGPIO_0/xhdl1.GEN_BITS[19].APB_32.INTR_reg_256_0_o2_0_0[19]  
        (.A(\CoreGPIO_0/CONFIG_reg[19][7] ), .B(
        \CoreGPIO_0/CONFIG_reg[19][6] ), .C(
        \CoreGPIO_0/CONFIG_reg[19][5] ), .D(
        \CoreGPIO_0/CONFIG_reg[19][3] ), .Y(
        \CoreGPIO_0/INTR_reg_256_0_o2_0[19] ));
    IOTRI_OB_EB \FIC_MSS_0/MDDR_ADDR_14_PAD/U_IOOUT  (.D(VCC), .E(VCC), 
        .DOUT(), .EOUT(\FIC_MSS_0/MDDR_ADDR_14_PAD/EOUT ));
    CFG3 #( .INIT(8'hF2) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_137  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_1_[1]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_502 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_137_i ));
    CFG4 #( .INIT(16'hAA08) )  
        \CoreGPIO_0/xhdl1.GEN_BITS[2].APB_32.edge_neg_37_iv_i_0[2]  (
        .A(\CoreGPIO_0/CONFIG_reg[2][3] ), .B(\CoreGPIO_0/edge_neg[2] )
        , .C(\CoreAPB3_0_APBmslave3_PWDATA[2] ), .D(\CoreGPIO_0/N_395 )
        , .Y(\CoreGPIO_0/N_119 ));
    CFG3 #( .INIT(8'hF2) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_235  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_13_[3]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_500 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_235_i ));
    CFG4 #( .INIT(16'h0F35) )  
        \CoreGPIO_0/CONFIG_reg_o_2_31_bm_1_RNO_1[5]  (.A(
        \CoreGPIO_0/CONFIG_reg[5][5] ), .B(
        \CoreGPIO_0/CONFIG_reg[21][5] ), .C(
        \CoreAPB3_0_APBmslave3_PADDR[6] ), .D(
        \CoreAPB3_0_APBmslave3_PADDR[5] ), .Y(
        \CoreGPIO_0/CONFIG_reg_o_2_21_1[5] ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[2].REG_GEN.CONFIG_reg[2][2]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[2] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB16_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[2]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB6_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[2][2] ));
    FLASH_FREEZE \flash_freeze_inst/INST_FLASH_FREEZE_IP  (
        .FF_TO_START(ff_to_start_net), .FF_DONE());
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_124_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB14_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_3__1_sqmuxa ), .ALn(
        AFLSDF_INV_63_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(GND)
        , .Q(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_124_set_net_1 ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[2].APB_32.edge_both[2]  (.D(
        \CoreGPIO_0/N_93 ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB17_rgbr_net_1 ), .EN(
        \CoreGPIO_0/N_86 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB7_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/edge_both[2] ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[17].REG_GEN.CONFIG_reg[17][1]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[1] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB16_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[17]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB6_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[17][1] ));
    CFG2 #( .INIT(4'h7) )  \CoreGPIO_0/edge_both_2_sqmuxa_13_i  (.A(
        \CoreGPIO_0/N_248 ), .B(\CoreGPIO_0/CONFIG_reg[29][3] ), .Y(
        \CoreGPIO_0/N_190 ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_271  (.A(VCC), 
        .B(VCC), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[31] ), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/FPGA_MDDR_ARESET_N_net ), .IPC());
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[20].REG_GEN.CONFIG_reg[20][3]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[3] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB12_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[20]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB2_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[20][3] ));
    CFG3 #( .INIT(8'hF2) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_156  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_3_[4]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_494 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_156_i ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[3].APB_32.INTR_reg[3]  (.D(
        \CoreGPIO_0/INTR_reg_48[3] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB10_rgbr_net_1 ), .EN(VCC), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB0_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0.xhdl1.GEN_BITS[3].APB_32.INTR_reg[3] ));
    CFG4 #( .INIT(16'hEFEE) )  
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_9[4]  (.A(
        \reg_apb_wrp_0/reg16x8_0/N_432 ), .B(
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_3[4]_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_1_[4]_net_1 ), .D(
        \reg_apb_wrp_0/reg16x8_0/N_502 ), .Y(
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_9[4]_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_10_[0]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[0] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB0_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_10__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_191_i ), .ADn(VCC), .SLn(
        VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_10_rs[0] ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_173  (.A(VCC), 
        .B(VCC), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/MMUART1_TXD_F2H_SCP_net ), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/MGPIO18B_F2H_GPIN_net ), .IPC());
    CFG3 #( .INIT(8'h7F) )  \FIC_MSS_0/MSS_ADLIB_INST_RNO_30  (.A(
        \CoreGPIO_0.xhdl1.GEN_BITS[6].gpin3[6] ), .B(
        \CoreGPIO_0.RDATA_32.un12_PRDATA_o ), .C(
        \CoreGPIO_0.xhdl1.GEN_BITS[6].REG_GEN.CONFIG_reg[6][1] ), .Y(
        \FIC_MSS_0/CoreAPB3_0_APBmslave5_PRDATA_m_0_1_0[6] ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[4].APB_32.edge_neg[4]  (.D(
        \CoreGPIO_0/N_117 ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB12_rgbr_net_1 ), .EN(
        \CoreGPIO_0/N_58 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB2_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/edge_neg[4] ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_195_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_99_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_195_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_195_rs_net_1 ));
    INV_BA AFLSDF_INV_4 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_89_net_1 ), .Y(
        AFLSDF_INV_4_net_1));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_69_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB18_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_8__1_sqmuxa ), .ALn(
        AFLSDF_INV_64_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(GND)
        , .Q(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_69_set_net_1 ));
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_108  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_13_[4]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_500 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_108_net_1 ));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/mem_10__RNIRVOI[4]  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_101_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_199_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_10_rs[4] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_10_[4]_net_1 ));
    CFG4 #( .INIT(16'h0F35) )  
        \CoreGPIO_0/CONFIG_reg_o_2_31_am_RNO_1[1]  (.A(
        \CoreGPIO_0.xhdl1.GEN_BITS[2].REG_GEN.CONFIG_reg[2][1] ), .B(
        \CoreGPIO_0/CONFIG_reg[18][1] ), .C(
        \CoreAPB3_0_APBmslave3_PADDR[6] ), .D(
        \CoreAPB3_0_APBmslave3_PADDR[5] ), .Y(
        \CoreGPIO_0/CONFIG_reg_o_2_10_1_1[1] ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[11].REG_GEN.CONFIG_reg[11][7]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[7] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB9_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[11]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_YR ), .ADn(VCC), .SLn(
        VCC), .SD(GND), .LAT(GND), .Q(\CoreGPIO_0/CONFIG_reg[11][7] ));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/mem_6__RNI8DDT[7]  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_123_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_202_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_6_rs[7] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_6_[7]_net_1 ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[19].APB_32.GPOUT_reg[19]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[19] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB10_rgbr_net_1 ), .EN(
        \CoreGPIO_0/GPOUT_reg_0_sqmuxa ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB0_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0.xhdl1.GEN_BITS[19].APB_32.GPOUT_reg[19] ));
    CFG3 #( .INIT(8'hF2) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_236  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_13_[4]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_500 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_236_i ));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/mem_3__RNI9T7Q[2]  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_126_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_154_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_3_rs[2] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_3_[2]_net_1 ));
    CFG3 #( .INIT(8'h20) )  
        \CoreGPIO_0/xhdl1.GEN_BITS[28].APB_32.edge_both_RNO[28]  (.A(
        \CoreGPIO_0/CONFIG_reg[28][3] ), .B(
        \CoreAPB3_0_APBmslave3_PWDATA[28] ), .C(
        \CoreGPIO_0/edge_pos[28] ), .Y(\CoreGPIO_0/N_87_i_0 ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[29].REG_GEN.CONFIG_reg[29][4]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[4] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB14_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[29]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB4_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[29][4] ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[4].REG_GEN.CONFIG_reg[4][7]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[7] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB12_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[4]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB2_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[4][7] ));
    RGB \FCCC_0/GL1_INST/U0_RGB1_RGB0  (.An(\FCCC_0/GL1_INST/U0_YNn ), 
        .ENn(GND), .YL(\FCCC_0/GL1_INST/U0_RGB1_RGB0_rgbl_net_1 ), .YR(
        ));
    SLE \reg_apb_wrp_0/reg16x8_0/temp_data[1]  (.D(
        \reg_apb_wrp_0/reg16x8_0/N_7_i_0 ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB12_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/rd_enable_net_1 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB2_rgbl_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/temp_data[1]_net_1 ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[27].REG_GEN.CONFIG_reg[27][0]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[0] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB9_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[27]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_YR ), .ADn(VCC), .SLn(
        VCC), .SD(GND), .LAT(GND), .Q(\CoreGPIO_0/CONFIG_reg[27][0] ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[21].REG_GEN.CONFIG_reg[21][3]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[3] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB13_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[21]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB3_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[21][3] ));
    CFG4 #( .INIT(16'h330A) )  
        \CoreGPIO_0/xhdl1.GEN_BITS[26].APB_32.INTR_reg_347_0[26]  (.A(
        \CoreGPIO_0.xhdl1.GEN_BITS[26].APB_32.INTR_reg[26] ), .B(
        \CoreGPIO_0/INTR_reg_347_0_o2_1[26] ), .C(
        \CoreAPB3_0_APBmslave3_PWDATA[26] ), .D(\CoreGPIO_0/N_248 ), 
        .Y(\CoreGPIO_0/INTR_reg_347[26] ));
    IO_DIFF \FIC_MSS_0/MDDR_CLK_PAD/U_IOP  (.YIN(GND));
    CFG2 #( .INIT(4'h7) )  \CoreGPIO_0/edge_both_2_sqmuxa_19_i  (.A(
        \CoreGPIO_0/N_248 ), .B(\CoreGPIO_0/CONFIG_reg[9][3] ), .Y(
        \CoreGPIO_0/N_182 ));
    sdf_IOPAD_TRI \FIC_MSS_0/MDDR_BA_1_PAD/U_IOPAD  (.PAD(MDDR_BA[1]), 
        .D(\FIC_MSS_0/DRAM_BA_net_0[1] ), .E(
        \FIC_MSS_0/MDDR_BA_1_PAD/EOUT ));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_5_[6]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[6] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB10_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_5__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_184_i ), .ADn(VCC), .SLn(
        VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_5_rs[6] ));
    CFG4 #( .INIT(16'h0F35) )  
        \CoreGPIO_0/CONFIG_reg_o_2_31_am_1_RNO_2[2]  (.A(
        \CoreGPIO_0/CONFIG_reg[0][2] ), .B(
        \CoreGPIO_0/CONFIG_reg[16][2] ), .C(
        \CoreAPB3_0_APBmslave3_PADDR[6] ), .D(
        \CoreAPB3_0_APBmslave3_PADDR[5] ), .Y(
        \CoreGPIO_0/CONFIG_reg_o_2_3_1[2] ));
    CFG4 #( .INIT(16'hEC00) )  \CoreAPB3_0/u_mux_p_to_b3/PRDATA[8]  (
        .A(\CoreGPIO_0.xhdl1.GEN_BITS[0].APB_32.GPOUT_reg9 ), .B(
        \CoreGPIO_0.N_570 ), .C(
        \CoreGPIO_0.xhdl1.GEN_BITS[8].APB_32.GPOUT_reg[8] ), .D(
        CoreAPB3_0_APBmslave5_PSELx), .Y(
        \FIC_MSS_0_FIC_0_APB_MASTER_PRDATA[8] ));
    sdf_IOPAD_IN \FIC_MSS_0/MMUART_0_RXD_PAD/U_IOPAD  (.PAD(
        MMUART_0_RXD), .Y(\FIC_MSS_0/MMUART_0_RXD_PAD_Y ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[30].APB_32.GPOUT_reg[30]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[30] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB13_rgbr_net_1 ), .EN(
        \CoreGPIO_0/GPOUT_reg_0_sqmuxa ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB3_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0.xhdl1.GEN_BITS[30].APB_32.GPOUT_reg[30] ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[2].APB_32.INTR_reg[2]  (.D(
        \CoreGPIO_0/INTR_reg_35[2] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB15_rgbr_net_1 ), .EN(VCC), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB5_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/INTR_reg[2] ));
    IOBI_IB_OB_EB \FIC_MSS_0/MDDR_DQ_10_PAD/U_IOBI  (.D(VCC), .E(VCC), 
        .YIN(\FIC_MSS_0/MDDR_DQ_10_PAD/YIN ), .DOUT(), .EOUT(), .Y());
    CFG3 #( .INIT(8'hF2) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_176  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_5_[2]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_490 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_176_i ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[11].REG_GEN.CONFIG_reg[11][6]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[6] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB9_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[11]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_YR ), .ADn(VCC), .SLn(
        VCC), .SD(GND), .LAT(GND), .Q(\CoreGPIO_0/CONFIG_reg[11][6] ));
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_49  (
        .A(\reg_apb_wrp_0/reg16x8_0/mem_7_[2]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_498 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_49_net_1 ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[3].APB_32.edge_pos[3]  (.D(
        \CoreGPIO_0/N_73 ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB9_rgbr_net_1 ), .EN(
        \CoreGPIO_0/N_79 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_YR ), .ADn(VCC), .SLn(
        VCC), .SD(GND), .LAT(GND), .Q(\CoreGPIO_0/edge_pos[3] ));
    CFG3 #( .INIT(8'hF2) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_248  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_15_[0]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_497 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_248_i ));
    CFG4 #( .INIT(16'h0F35) )  
        \CoreGPIO_0/CONFIG_reg_o_2_31_am_RNO_1[6]  (.A(
        \CoreGPIO_0/CONFIG_reg[2][6] ), .B(
        \CoreGPIO_0/CONFIG_reg[18][6] ), .C(
        \CoreAPB3_0_APBmslave3_PADDR[6] ), .D(
        \CoreAPB3_0_APBmslave3_PADDR[5] ), .Y(
        \CoreGPIO_0/CONFIG_reg_o_2_10_1_1[6] ));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_8_[1]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[1] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB4_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_8__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_221_i ), .ADn(VCC), .SLn(
        VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_8_rs[1] ));
    CFG2 #( .INIT(4'h6) )  
        \CoreGPIO_0/xhdl1.GEN_BITS[6].APB_32.edge_both_93_iv_i_0_i_x2[6]  
        (.A(\CoreGPIO_0/gpin2[6] ), .B(
        \CoreGPIO_0.xhdl1.GEN_BITS[6].gpin3[6] ), .Y(
        \CoreGPIO_0/N_252_i ));
    CFG4 #( .INIT(16'hC480) )  
        \CoreGPIO_0/xhdl1.GEN_BITS[1].APB_32.INTR_reg_22_0_0_RNO[1]  (
        .A(\CoreGPIO_0/CONFIG_reg[1][7] ), .B(
        \CoreGPIO_0/CONFIG_reg[1][3] ), .C(
        \CoreGPIO_0/INTR_reg_22_0_0_51_tz_1 ), .D(\CoreGPIO_0/N_177 ), 
        .Y(\CoreGPIO_0/N_1576_tz ));
    INV_BA AFLSDF_INV_24 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_79_net_1 ), .Y(
        AFLSDF_INV_24_net_1));
    CFG3 #( .INIT(8'hF2) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_200  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_6_[6]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_493 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_200_i ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[9].REG_GEN.CONFIG_reg[9][5]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[5] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB15_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[9]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB5_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[9][5] ));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_223_rs_RNIS0EV  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_64_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_223_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_8_rs[2] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_8_[2]_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_1_[3]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[3] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB15_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_1__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_139_i ), .ADn(VCC), .SLn(
        VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_1_rs[3] ));
    INV_BA AFLSDF_INV_84 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_29_net_1 ), .Y(
        AFLSDF_INV_84_net_1));
    CFG4 #( .INIT(16'h4657) )  
        \CoreGPIO_0/CONFIG_reg_o_2_31_am_1_1[0]  (.A(
        \CoreAPB3_0_APBmslave3_PADDR[4] ), .B(
        \CoreAPB3_0_APBmslave3_PADDR[3] ), .C(
        \CoreGPIO_0/CONFIG_reg_o_2_31_am_1_1_RNO[0]_net_1 ), .D(
        \CoreGPIO_0/CONFIG_reg_o_2_31_am_1_RNO_0[0]_net_1 ), .Y(
        \CoreGPIO_0/CONFIG_reg_o_2_31_am_1[0] ));
    CFG4 #( .INIT(16'hC5CA) )  
        \CoreGPIO_0/xhdl1.GEN_BITS[3].REG_INT.un34_intr_u_bm  (.A(
        \CoreGPIO_0.xhdl1.GEN_BITS[3].gpin3[3] ), .B(
        \CoreGPIO_0/N_4549 ), .C(\CoreGPIO_0/CONFIG_reg[3][6] ), .D(
        \CoreGPIO_0/CONFIG_reg[3][5] ), .Y(\CoreGPIO_0/un34_intr_u_bm )
        );
    SLE \reg_apb_wrp_0/reg16x8_0/mem_2_[5]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[5] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB15_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_2__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_149_i ), .ADn(VCC), .SLn(
        VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_2_rs[5] ));
    INV_BA AFLSDF_INV_50 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_99_net_1 ), .Y(
        AFLSDF_INV_50_net_1));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[25].APB_32.edge_both[25]  (.D(
        \CoreGPIO_0/N_5911_i_0 ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB14_rgbr_net_1 ), .EN(
        \CoreGPIO_0/N_157 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB4_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/edge_neg[25] ));
    CFG4 #( .INIT(16'hA9FF) )  
        \CoreGPIO_0/xhdl1.GEN_BITS[9].APB_32.INTR_reg_126_0_o2_0_0[9]  
        (.A(\CoreGPIO_0/CONFIG_reg[9][7] ), .B(
        \CoreGPIO_0/CONFIG_reg[9][6] ), .C(
        \CoreGPIO_0/CONFIG_reg[9][5] ), .D(
        \CoreGPIO_0/CONFIG_reg[9][3] ), .Y(
        \CoreGPIO_0/INTR_reg_126_0_o2_0[9] ));
    CFG4 #( .INIT(16'hFF4F) )  \CoreGPIO_0/edge_both_2_sqmuxa_i_0  (.A(
        \CoreGPIO_0.N_247 ), .B(\CoreGPIO_0/INTR_reg21 ), .C(
        \CoreGPIO_0/CONFIG_reg[2][3] ), .D(\CoreGPIO_0/N_144_i ), .Y(
        \CoreGPIO_0/N_86 ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_5  (.A(
        \FIC_MSS_0/FIC_MSS_0_FIC_0_APB_MASTER_PRDATA[3] ), .B(
        \FIC_MSS_0_FIC_0_APB_MASTER_PRDATA[10] ), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[3] ), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[10] ), .IPC());
    CFG3 #( .INIT(8'hF2) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_202  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_6_[7]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_493 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_202_i ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_200  (.A(VCC), 
        .B(VCC), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[4] ), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[16] ), .IPC());
    CFG4 #( .INIT(16'hEC00) )  \CoreAPB3_0/u_mux_p_to_b3/PRDATA[21]  (
        .A(\CoreGPIO_0.xhdl1.GEN_BITS[0].APB_32.GPOUT_reg9 ), .B(
        \CoreGPIO_0.N_544 ), .C(
        \CoreGPIO_0.xhdl1.GEN_BITS[21].APB_32.GPOUT_reg[21] ), .D(
        CoreAPB3_0_APBmslave5_PSELx), .Y(
        \FIC_MSS_0_FIC_0_APB_MASTER_PRDATA[21] ));
    CFG4 #( .INIT(16'hAC0F) )  
        \CoreGPIO_0/CONFIG_reg_o_2_31_bm_1_RNO_0[0]  (.A(
        \CoreGPIO_0/CONFIG_reg[9][0] ), .B(
        \CoreGPIO_0/CONFIG_reg[25][0] ), .C(
        \CoreGPIO_0/CONFIG_reg_o_2_18_1[0] ), .D(
        \CoreAPB3_0_APBmslave3_PADDR[5] ), .Y(
        \CoreGPIO_0/CONFIG_reg_o_2_31_bm_1_RNO_0[0]_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_116_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB9_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_14__1_sqmuxa ), .ALn(
        AFLSDF_INV_65_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(GND)
        , .Q(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_116_set_net_1 ));
    sdf_IOPAD_BI \FIC_MSS_0/MDDR_DQ_9_PAD/U_IOPAD  (.PAD(MDDR_DQ[9]), 
        .D(\FIC_MSS_0/DRAM_DQ_OUT_net_0[9] ), .E(
        \FIC_MSS_0/DRAM_DQ_OE_net_0[9] ), .Y(
        \FIC_MSS_0/MDDR_DQ_9_PAD_Y ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_102_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB11_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_10__1_sqmuxa ), .ALn(
        AFLSDF_INV_66_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(GND)
        , .Q(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_102_set_net_1 ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[7].REG_GEN.CONFIG_reg[7][4]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[4] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB10_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[7]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB0_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[7][4] ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_207  (.A(VCC), 
        .B(GND), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[25] ), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/F_AWLEN_HBURST0_net[3] ), .IPC());
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_278  (.A(VCC), 
        .B(VCC), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[2] ), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[5] ), .IPC());
    CFG4 #( .INIT(16'h4657) )  
        \CoreGPIO_0/CONFIG_reg_o_2_31_bm_1_1[5]  (.A(
        \CoreAPB3_0_APBmslave3_PADDR[4] ), .B(
        \CoreAPB3_0_APBmslave3_PADDR[3] ), .C(
        \CoreGPIO_0/CONFIG_reg_o_2_31_bm_1_1_RNO[5]_net_1 ), .D(
        \CoreGPIO_0/CONFIG_reg_o_2_31_bm_1_RNO_0[5]_net_1 ), .Y(
        \CoreGPIO_0/CONFIG_reg_o_2_31_bm_1[5] ));
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_103  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_10_[6]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_491 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_103_net_1 ));
    CFG4 #( .INIT(16'hAC0F) )  
        \CoreGPIO_0/CONFIG_reg_o_2_31_bm_RNO_0[1]  (.A(
        \CoreGPIO_0/CONFIG_reg[15][1] ), .B(
        \CoreGPIO_0/CONFIG_reg[31][1] ), .C(
        \CoreGPIO_0/CONFIG_reg_o_2_28_1_1[1] ), .D(
        \CoreAPB3_0_APBmslave3_PADDR[5] ), .Y(
        \CoreGPIO_0/CONFIG_reg_o_2_31_bm_RNO_0[1]_net_1 ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_4  (.A(
        \FIC_MSS_0/FIC_MSS_0_FIC_0_APB_MASTER_PRDATA[2] ), .B(
        \FIC_MSS_0_FIC_0_APB_MASTER_PRDATA[9] ), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[2] ), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[9] ), .IPC());
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_249  (.A(VCC), 
        .B(GND), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[61] ), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/F_ARID_HSEL1_net[1] ), .IPC());
    SLE \reg_apb_wrp_0/rd_enable  (.D(\reg_apb_wrp_0/N_76 ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB12_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/N_45_i_0 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB2_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/rd_enable_net_1 ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_0  (.A(
        \FIC_MSS_0/FIC_MSS_0_FIC_0_APB_MASTER_PREADY1_i_m_i_0 ), .B(
        VCC), .C(VCC), .IPA(\FIC_MSS_0/MSS_ADLIB_INST/F_HM0_READY_net )
        , .IPB(), .IPC());
    sdf_IOPAD_BI \FIC_MSS_0/MDDR_DM_RDQS_1_PAD/U_IOPAD  (.PAD(
        MDDR_DM_RDQS[1]), .D(\FIC_MSS_0/DRAM_DM_RDQS_OUT_net_0[1] ), 
        .E(\FIC_MSS_0/DM_OE_net_0[1] ), .Y(
        \FIC_MSS_0/MDDR_DM_RDQS_1_PAD_Y ));
    CFG4 #( .INIT(16'hF2F3) )  
        \CoreGPIO_0/xhdl1.GEN_BITS[10].APB_32.INTR_reg_139_0_o2_1_0[10]  
        (.A(\CoreGPIO_0/CONFIG_reg[10][6] ), .B(
        \CoreGPIO_0/edge_pos[10] ), .C(
        \CoreGPIO_0/INTR_reg_139_0_o2_0[10] ), .D(
        \CoreGPIO_0/CONFIG_reg[10][5] ), .Y(
        \CoreGPIO_0/INTR_reg_139_0_o2_1[10] ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_72_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB14_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_9__1_sqmuxa ), .ALn(
        AFLSDF_INV_67_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(GND)
        , .Q(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_72_set_net_1 ));
    RGB \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB7  (.An(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_YNn_GSouth ), .ENn(GND), .YL()
        , .YR(\MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB7_rgbr_net_1 ));
    CFG2 #( .INIT(4'h4) )  \CoreGPIO_0/PRDATA_0_iv_0_a2_0[31]  (.A(
        \CoreGPIO_0.N_247 ), .B(\CoreGPIO_0/INTR_reg[31] ), .Y(
        \CoreGPIO_0.N_524 ));
    CFG4 #( .INIT(16'hEFEE) )  
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_9[0]  (.A(
        \reg_apb_wrp_0/reg16x8_0/N_366 ), .B(
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_3[0]_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_1_[0]_net_1 ), .D(
        \reg_apb_wrp_0/reg16x8_0/N_502 ), .Y(
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_9[0]_net_1 ));
    CFG2 #( .INIT(4'h8) )  
        \reg_apb_wrp_0/reg16x8_0/mem_15__1_sqmuxa_0_a3  (.A(
        \reg_apb_wrp_0/reg16x8_0/N_497 ), .B(
        \reg_apb_wrp_0/wr_enable_net_1 ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_15__1_sqmuxa ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_100_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB11_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_10__1_sqmuxa ), .ALn(
        AFLSDF_INV_68_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(GND)
        , .Q(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_100_set_net_1 ));
    sdf_IOPAD_BI \FIC_MSS_0/MDDR_DQ_7_PAD/U_IOPAD  (.PAD(MDDR_DQ[7]), 
        .D(\FIC_MSS_0/DRAM_DQ_OUT_net_0[7] ), .E(
        \FIC_MSS_0/DRAM_DQ_OE_net_0[7] ), .Y(
        \FIC_MSS_0/MDDR_DQ_7_PAD_Y ));
    CFG4 #( .INIT(16'h0F35) )  
        \CoreGPIO_0/CONFIG_reg_o_2_31_am_RNO_2[4]  (.A(
        \CoreGPIO_0/CONFIG_reg[6][4] ), .B(
        \CoreGPIO_0/CONFIG_reg[22][4] ), .C(
        \CoreAPB3_0_APBmslave3_PADDR[6] ), .D(
        \CoreAPB3_0_APBmslave3_PADDR[5] ), .Y(
        \CoreGPIO_0/CONFIG_reg_o_2_13_1_1[4] ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_90_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB16_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_11__1_sqmuxa ), .ALn(
        AFLSDF_INV_69_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(GND)
        , .Q(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_90_set_net_1 ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_186  (.A(VCC), 
        .B(VCC), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/MGPIO29B_F2H_GPIN_net ), .IPB(), 
        .IPC());
    CFG4 #( .INIT(16'hB383) )  \CoreGPIO_0/CONFIG_reg_o_2_31_am[5]  (
        .A(\CoreGPIO_0/CONFIG_reg_o_2_31_am_RNO[5]_net_1 ), .B(
        \CoreGPIO_0/CONFIG_reg_o_2_31_am_1[5] ), .C(
        \CoreAPB3_0_APBmslave3_PADDR[3] ), .D(
        \CoreGPIO_0/CONFIG_reg_o_2_31_am_RNO_0[5]_net_1 ), .Y(
        \CoreGPIO_0/CONFIG_reg_o_2_31_am[5]_net_1 ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_225  (.A(VCC), 
        .B(VCC), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[9] ), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[21] ), .IPC());
    CFG4 #( .INIT(16'h0400) )  
        \CoreGPIO_0/xhdl1.GEN_BITS[4].REG_GEN.CONFIG_reg[4]2_0_a4_0_a2  
        (.A(\CoreAPB3_0_APBmslave3_PADDR[7] ), .B(\CoreGPIO_0/N_603 ), 
        .C(\CoreGPIO_0/N_243 ), .D(\CoreGPIO_0/INTR_reg21 ), .Y(
        \CoreGPIO_0/CONFIG_reg[4]2 ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[29].REG_GEN.CONFIG_reg[29][6]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[6] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB13_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[29]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB3_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[29][6] ));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_117_set_RNIVIV7  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_117_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_245_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_14_rs[5] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_14_[5]_net_1 ));
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_101  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_10_[4]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_491 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_101_net_1 ));
    CFG2 #( .INIT(4'h2) )  
        \CoreGPIO_0/xhdl1.GEN_BITS[8].REG_GEN.CONFIG_reg[8]2_0_a4_0_a2_0  
        (.A(\CoreAPB3_0_APBmslave3_PADDR[5] ), .B(
        \CoreAPB3_0_APBmslave3_PADDR[4] ), .Y(\CoreGPIO_0/N_610 ));
    CFG3 #( .INIT(8'hF2) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_162  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_4_[1]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_504 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_162_i ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_78  (.A(VCC), 
        .B(VCC), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[12] ), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[19] ), .IPC());
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_45  (
        .A(\reg_apb_wrp_0/reg16x8_0/mem_1_[6]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_502 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_45_net_1 ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[0].REG_GEN.CONFIG_reg[0][3]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[3] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB11_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[0]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB1_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[0][3] ));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_2_[7]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[7] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB12_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_2__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_151_i ), .ADn(VCC), .SLn(
        VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_2_rs[7] ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_42_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB5_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_5__1_sqmuxa ), .ALn(
        AFLSDF_INV_70_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(GND)
        , .Q(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_42_set_net_1 ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[11].REG_GEN.CONFIG_reg[11][1]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[1] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB10_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[11]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB0_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[11][1] ));
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_30  (
        .A(\reg_apb_wrp_0/reg16x8_0/mem_2_[2]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_501 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_30_net_1 ));
    CFG2 #( .INIT(4'h7) )  \CoreGPIO_0/edge_both_2_sqmuxa_24_i  (.A(
        \CoreGPIO_0/N_248 ), .B(\CoreGPIO_0/CONFIG_reg[31][3] ), .Y(
        \CoreGPIO_0/edge_pos_2_sqmuxa_19_i_1 ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_219  (.A(VCC), 
        .B(VCC), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[3] ), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[15] ), .IPC());
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[26].REG_GEN.CONFIG_reg[26][1]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[1] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB16_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[26]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB6_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[26][1] ));
    CFG2 #( .INIT(4'h8) )  
        \CoreGPIO_0/xhdl1.GEN_BITS[1].REG_GPOUT.un14_GPIO_OUT_i  (.A(
        \CoreGPIO_0.xhdl1.GEN_BITS[1].APB_32.GPOUT_reg[1] ), .B(
        \CoreGPIO_0/CONFIG_reg[1][0] ), .Y(\GPIO_OUT_net_2[1] ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[5].APB_32.edge_both[5]  (.D(
        \CoreGPIO_0/N_89 ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB10_rgbr_net_1 ), .EN(
        \CoreGPIO_0/N_76 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB0_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/edge_both[5] ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[31].REG_GEN.CONFIG_reg[31][3]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[3] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB10_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[31]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB0_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[31][3] ));
    CFG4 #( .INIT(16'hEC00) )  \CoreAPB3_0/u_mux_p_to_b3/PRDATA[28]  (
        .A(\CoreGPIO_0.xhdl1.GEN_BITS[0].APB_32.GPOUT_reg9 ), .B(
        \CoreGPIO_0.N_530 ), .C(
        \CoreGPIO_0.xhdl1.GEN_BITS[28].APB_32.GPOUT_reg[28] ), .D(
        CoreAPB3_0_APBmslave5_PSELx), .Y(
        \FIC_MSS_0_FIC_0_APB_MASTER_PRDATA[28] ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_122  (.A(VCC), 
        .B(VCC), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/FAB_SESSEND_net ), .IPB(), .IPC());
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_281  (.A(VCC), 
        .B(VCC), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PADDR_net[4] ), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[8] ), .IPC());
    CFG3 #( .INIT(8'h04) )  
        \CoreGPIO_0/xhdl1.GEN_BITS[0].APB_32.INTR_reg_9_0_0_RNO_0[0]  
        (.A(\CoreGPIO_0/CONFIG_reg[0][5] ), .B(
        \CoreGPIO_0/edge_both[0] ), .C(\CoreGPIO_0/CONFIG_reg[0][6] ), 
        .Y(\CoreGPIO_0/INTR_reg_9_0_0_50_tz_1 ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[26].REG_GEN.CONFIG_reg[26][7]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[7] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB17_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[26]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB7_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[26][7] ));
    CFG3 #( .INIT(8'hFE) )  
        \CoreGPIO_0/xhdl1.GEN_BITS[0].APB_32.un5_PRDATA_o_0_a2_0_o2  (
        .A(\CoreAPB3_0_APBmslave3_PADDR[6] ), .B(
        \CoreGPIO_0.RDATA_32.un12_PRDATA_o_0_o2_1 ), .C(
        \CoreGPIO_0/un5_PRDATA_o_0_a2_0_o2_sx ), .Y(\CoreGPIO_0.N_247 )
        );
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_93_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB19_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_11__1_sqmuxa ), .ALn(
        AFLSDF_INV_71_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(GND)
        , .Q(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_93_set_net_1 ));
    CFG3 #( .INIT(8'hF2) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_228  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_12_[4]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_495 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_228_i ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[10].REG_GEN.CONFIG_reg[10][0]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[0] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB16_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[10]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB6_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[10][0] ));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_74_set_RNI8B5V  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_74_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_179_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_9_rs[2] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_9_[2]_net_1 ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_36  (.A(GND), 
        .B(VCC), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[19] ), .IPB(), .IPC());
    CFG4 #( .INIT(16'hA9FF) )  
        \CoreGPIO_0/xhdl1.GEN_BITS[21].APB_32.INTR_reg_282_0_o2_0_0[21]  
        (.A(\CoreGPIO_0/CONFIG_reg[21][7] ), .B(
        \CoreGPIO_0/CONFIG_reg[21][6] ), .C(
        \CoreGPIO_0/CONFIG_reg[21][5] ), .D(
        \CoreGPIO_0/CONFIG_reg[21][3] ), .Y(
        \CoreGPIO_0/INTR_reg_282_0_o2_0[21] ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[29].REG_GEN.CONFIG_reg[29][1]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[1] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB13_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[29]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB3_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[29][1] ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_27  (.A(GND), 
        .B(GND), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[3] ), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[10] ), .IPC());
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_183  (.A(VCC), 
        .B(VCC), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/MMUART0_TXD_F2H_SCP_net ), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/MMUART0_RI_F2H_SCP_net ), .IPC());
    CFG4 #( .INIT(16'hEC00) )  \CoreAPB3_0/u_mux_p_to_b3/PRDATA[24]  (
        .A(\CoreGPIO_0.xhdl1.GEN_BITS[0].APB_32.GPOUT_reg9 ), .B(
        \CoreGPIO_0.N_538 ), .C(
        \CoreGPIO_0.xhdl1.GEN_BITS[24].APB_32.GPOUT_reg[24] ), .D(
        CoreAPB3_0_APBmslave5_PSELx), .Y(
        \FIC_MSS_0_FIC_0_APB_MASTER_PRDATA[24] ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_57_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB7_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_15__1_sqmuxa ), .ALn(
        AFLSDF_INV_72_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(GND)
        , .Q(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_57_set_net_1 ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[29].REG_GEN.CONFIG_reg[29][3]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[3] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB13_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[29]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB3_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[29][3] ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[31].REG_GEN.CONFIG_reg[31][6]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[6] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB10_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[31]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB0_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[31][6] ));
    CFG4 #( .INIT(16'hAC0F) )  
        \CoreGPIO_0/CONFIG_reg_o_2_31_bm_RNO[0]  (.A(
        \CoreGPIO_0/CONFIG_reg[11][0] ), .B(
        \CoreGPIO_0/CONFIG_reg[27][0] ), .C(
        \CoreGPIO_0/CONFIG_reg_o_2_25_1_1[0] ), .D(
        \CoreAPB3_0_APBmslave3_PADDR[5] ), .Y(
        \CoreGPIO_0/CONFIG_reg_o_2_31_bm_RNO[0]_net_1 ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[20].APB_32.edge_both[20]  (.D(
        \CoreGPIO_0/edge_neg_289[20] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB11_rgbr_net_1 ), .EN(
        \CoreGPIO_0/N_196 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB1_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/edge_neg[20] ));
    CFG2 #( .INIT(4'h2) )  \CoreGPIO_0/edge_pos_2_sqmuxa_4_i_a2  (.A(
        \CoreGPIO_0/gpin2[4] ), .B(
        \CoreGPIO_0.xhdl1.GEN_BITS[4].gpin3[4] ), .Y(
        \CoreGPIO_0/N_398 ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[24].REG_GEN.CONFIG_reg[24][7]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[7] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB11_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[24]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB1_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[24][7] ));
    CFG4 #( .INIT(16'hAC0F) )  
        \CoreGPIO_0/CONFIG_reg_o_2_31_am_RNO[6]  (.A(
        \CoreGPIO_0/CONFIG_reg[10][6] ), .B(
        \CoreGPIO_0/CONFIG_reg[26][6] ), .C(
        \CoreGPIO_0/CONFIG_reg_o_2_10_1_1[6] ), .D(
        \CoreAPB3_0_APBmslave3_PADDR[5] ), .Y(
        \CoreGPIO_0/CONFIG_reg_o_2_31_am_RNO[6]_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_156_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_50_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_156_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_156_rs_net_1 ));
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_83  (
        .A(\reg_apb_wrp_0/reg16x8_0/mem_3_[6]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_494 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_83_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/temp_data[2]  (.D(
        \reg_apb_wrp_0/reg16x8_0/N_9_i_0 ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB12_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/rd_enable_net_1 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB2_rgbl_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/temp_data[2]_net_1 ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_148  (.A(VCC), 
        .B(VCC), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/MGPIO1A_F2H_GPIN_net ), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/CAN_TX_EBL_F2H_SCP_net ), .IPC());
    CFG4 #( .INIT(16'hAC0F) )  
        \CoreGPIO_0/CONFIG_reg_o_2_31_am_1_1_RNO[2]  (.A(
        \CoreGPIO_0/CONFIG_reg[12][2] ), .B(
        \CoreGPIO_0/CONFIG_reg[28][2] ), .C(
        \CoreGPIO_0/CONFIG_reg_o_2_6_1[2] ), .D(
        \CoreAPB3_0_APBmslave3_PADDR[5] ), .Y(
        \CoreGPIO_0/CONFIG_reg_o_2_31_am_1_1_RNO[2]_net_1 ));
    INV_BA AFLSDF_INV_5 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_75_net_1 ), .Y(
        AFLSDF_INV_5_net_1));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_272  (.A(GND), 
        .B(GND), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/F_ARLEN_HBURST1_net[0] ), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/F_RMW_AXI_net ), .IPC());
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_21_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB10_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_12__1_sqmuxa ), .ALn(
        AFLSDF_INV_73_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(GND)
        , .Q(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_21_set_net_1 ));
    CFG4 #( .INIT(16'h7350) )  
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_3[2]  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_11_[2]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/mem_3_[2]_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/N_505 ), .D(
        \reg_apb_wrp_0/reg16x8_0/N_494 ), .Y(
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_3[2]_net_1 ));
    IOTRI_OB_EB \FIC_MSS_0/MDDR_ADDR_15_PAD/U_IOOUT  (.D(VCC), .E(VCC), 
        .DOUT(), .EOUT(\FIC_MSS_0/MDDR_ADDR_15_PAD/EOUT ));
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_47  (
        .A(\reg_apb_wrp_0/reg16x8_0/mem_1_[5]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_502 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_47_net_1 ));
    CFG4 #( .INIT(16'h330A) )  
        \CoreGPIO_0/xhdl1.GEN_BITS[31].APB_32.INTR_reg_412_0[31]  (.A(
        \CoreGPIO_0/INTR_reg[31] ), .B(
        \CoreGPIO_0/INTR_reg_412_0_o2_1[31] ), .C(
        \CoreAPB3_0_APBmslave3_PWDATA[31] ), .D(\CoreGPIO_0/N_248 ), 
        .Y(\CoreGPIO_0/INTR_reg_412[31] ));
    CFG2 #( .INIT(4'h7) )  \CoreGPIO_0/edge_both_2_sqmuxa_26_i  (.A(
        \CoreGPIO_0/N_248 ), .B(\CoreGPIO_0/CONFIG_reg[23][3] ), .Y(
        \CoreGPIO_0/edge_pos_2_sqmuxa_26_i_1 ));
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_112  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_14_[0]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_503 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_112_net_1 ));
    INV_BA AFLSDF_INV_64 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_69_net_1 ), .Y(
        AFLSDF_INV_64_net_1));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_163_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_4_net_1 ), .EN(VCC), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_163_i ), .ADn(VCC), .SLn(
        VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_163_rs_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_3_[0]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[0] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB14_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_3__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_152_i ), .ADn(VCC), .SLn(
        VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_3_rs[0] ));
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_93  (
        .A(\reg_apb_wrp_0/reg16x8_0/mem_11_[5]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_505 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_93_net_1 ));
    CFG3 #( .INIT(8'hDF) )  \CoreGPIO_0/edge_pos_2_sqmuxa_18_i_0  (.A(
        \CoreGPIO_0/CONFIG_reg[3][3] ), .B(\CoreGPIO_0/N_687 ), .C(
        \CoreGPIO_0/N_248 ), .Y(\CoreGPIO_0/N_79 ));
    IP_INTERFACE \FCCC_0/CCC_INST/IP_INTERFACE_3  (.A(GND), .B(GND), 
        .C(VCC), .IPA(\FCCC_0/CCC_INST/PRESET_N_net ), .IPB(
        \FCCC_0/CCC_INST/NGMUX1_SEL_net ), .IPC(
        \FCCC_0/CCC_INST/PWDATA_net[1] ));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_140_rs_RNIGALR  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_41_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_140_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_1_rs[4] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_1_[4]_net_1 ));
    CFG4 #( .INIT(16'h0F35) )  
        \CoreGPIO_0/CONFIG_reg_o_2_31_am_1_RNO_2[4]  (.A(
        \CoreGPIO_0/CONFIG_reg[0][4] ), .B(
        \CoreGPIO_0/CONFIG_reg[16][4] ), .C(
        \CoreAPB3_0_APBmslave3_PADDR[6] ), .D(
        \CoreAPB3_0_APBmslave3_PADDR[5] ), .Y(
        \CoreGPIO_0/CONFIG_reg_o_2_3_1[4] ));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_5_[3]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[3] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB5_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_5__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_178_i ), .ADn(VCC), .SLn(
        VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_5_rs[3] ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_177  (.A(VCC), 
        .B(VCC), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/MMUART1_RXD_F2H_SCP_net ), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/MGPIO20B_F2H_GPIN_net ), .IPC());
    sdf_IOPADP_BI \FIC_MSS_0/MDDR_DQS_0_PAD/U_IOPADP  (.PAD_P(
        MDDR_DQS[0]), .N2PIN_P(\FIC_MSS_0/MDDR_DQS_0_PAD/U2_N2P ), 
        .OIN_P(\FIC_MSS_0/DRAM_DQS_OUT_net_0[0] ), .EIN_P(
        \FIC_MSS_0/DRAM_DQS_OE_net_0[0] ), .IOUT_P(
        \FIC_MSS_0/MDDR_DQS_0_PAD_Y ));
    CFG4 #( .INIT(16'h7350) )  
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_0_6[5]  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_8_[5]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/mem_0_[5]_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/N_499 ), .D(
        \reg_apb_wrp_0/reg16x8_0/N_496 ), .Y(
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_0_6[5]_net_1 ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[29].REG_GEN.CONFIG_reg[29][2]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[2] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB14_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[29]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB4_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[29][2] ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[17].APB_32.INTR_reg[17]  (.D(
        \CoreGPIO_0/INTR_reg_230[17] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB14_rgbr_net_1 ), .EN(VCC), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB4_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/INTR_reg[17] ));
    IOINFF_BYPASS \GPIO_IN_ibuf[0]/U0/U_IOINFF  (.A(
        \GPIO_IN_ibuf[0]/U0/YIN1 ), .Y(\GPIO_IN_ibuf[0]/U0/YIN ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[18].REG_GEN.CONFIG_reg[18][4]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[4] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB17_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[18]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB7_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[18][4] ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_74_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB15_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_9__1_sqmuxa ), .ALn(
        AFLSDF_INV_74_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(GND)
        , .Q(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_74_set_net_1 ));
    CFG3 #( .INIT(8'h20) )  
        \CoreGPIO_0/xhdl1.GEN_BITS[21].APB_32.edge_both_RNO[21]  (.A(
        \CoreGPIO_0/CONFIG_reg[21][3] ), .B(
        \CoreAPB3_0_APBmslave3_PWDATA[21] ), .C(
        \CoreGPIO_0/edge_neg[21] ), .Y(\CoreGPIO_0/edge_neg_303[21] ));
    CFG4 #( .INIT(16'hEC00) )  \CoreAPB3_0/u_mux_p_to_b3/PRDATA[20]  (
        .A(\CoreGPIO_0.xhdl1.GEN_BITS[0].APB_32.GPOUT_reg9 ), .B(
        \CoreGPIO_0.N_546 ), .C(
        \CoreGPIO_0.xhdl1.GEN_BITS[20].APB_32.GPOUT_reg[20] ), .D(
        CoreAPB3_0_APBmslave5_PSELx), .Y(
        \FIC_MSS_0_FIC_0_APB_MASTER_PRDATA[20] ));
    INV_BA AFLSDF_INV_73 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_21_net_1 ), .Y(
        AFLSDF_INV_73_net_1));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/mem_15__RNIHSDR[0]  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_57_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_248_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_15_rs[0] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_15_[0]_net_1 ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_118  (.A(VCC), 
        .B(VCC), .C(VCC), .IPA(), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/FAB_VSTATUS_net[7] ), .IPC());
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_1  (.A(GND), 
        .B(VCC), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/F_HM0_RESP_net ), .IPB(), .IPC());
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_161  (.A(VCC), 
        .B(VCC), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/SPI1_SDI_F2H_SCP_net ), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/SPI1_SS1_F2H_SCP_net ), .IPC());
    CFG3 #( .INIT(8'h01) )  \reg_apb_wrp_0/reg16x8_0/temp_data_RNO[1]  
        (.A(\reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_8[1]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_13[1]_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_9[1]_net_1 ), .Y(
        \reg_apb_wrp_0/reg16x8_0/N_7_i_0 ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_113_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB6_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_14__1_sqmuxa ), .ALn(
        AFLSDF_INV_75_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(GND)
        , .Q(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_113_set_net_1 ));
    IOTRI_OB_EB \GPIO_OUT_obuf[2]/U0/U_IOTRI  (.D(\GPIO_OUT_net_2[2] ), 
        .E(VCC), .DOUT(\GPIO_OUT_obuf[2]/U0/DOUT1 ), .EOUT(
        \GPIO_OUT_obuf[2]/U0/EOUT1 ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[30].REG_GEN.CONFIG_reg[30][2]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[2] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB14_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[30]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB4_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[30][2] ));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_159_rs_RNI4GOJ  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_83_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_159_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_3_rs[6] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_3_[6]_net_1 ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[9].APB_32.edge_both[9]  (.D(
        \CoreGPIO_0/edge_neg_135[9] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB14_rgbr_net_1 ), .EN(
        \CoreGPIO_0/N_182 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB4_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/edge_neg[9] ));
    CFG4 #( .INIT(16'h4657) )  
        \CoreGPIO_0/CONFIG_reg_o_2_31_bm_1_1[0]  (.A(
        \CoreAPB3_0_APBmslave3_PADDR[4] ), .B(
        \CoreAPB3_0_APBmslave3_PADDR[3] ), .C(
        \CoreGPIO_0/CONFIG_reg_o_2_31_bm_1_1_RNO[0]_net_1 ), .D(
        \CoreGPIO_0/CONFIG_reg_o_2_31_bm_1_RNO_0[0]_net_1 ), .Y(
        \CoreGPIO_0/CONFIG_reg_o_2_31_bm_1[0] ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_170_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_11_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_170_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_170_rs_net_1 ));
    CFG2 #( .INIT(4'h6) )  \CoreGPIO_0/edge_both_2_sqmuxa_i_x2  (.A(
        \CoreGPIO_0/gpin2[2] ), .B(
        \CoreGPIO_0.xhdl1.GEN_BITS[2].gpin3[2] ), .Y(
        \CoreGPIO_0/N_144_i ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_144  (.A(
        FCCC_0_LOCK), .B(VCC), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/FAB_PLL_LOCK_net ), .IPB(), .IPC());
    IP_INTERFACE \FCCC_0/CCC_INST/IP_INTERFACE_2  (.A(VCC), .B(GND), 
        .C(VCC), .IPA(\FCCC_0/CCC_INST/PCLK_net ), .IPB(
        \FCCC_0/CCC_INST/NGMUX0_SEL_net ), .IPC(
        \FCCC_0/CCC_INST/PWDATA_net[0] ));
    IOBI_IB_OB_EB \FIC_MSS_0/MDDR_DQ_9_PAD/U_IOBI  (.D(VCC), .E(VCC), 
        .YIN(\FIC_MSS_0/MDDR_DQ_9_PAD/YIN ), .DOUT(), .EOUT(), .Y());
    RGB \FCCC_0/GL1_INST/U0_RGB1_RGB14  (.An(
        \FCCC_0/GL1_INST/U0_YNn_GSouth ), .ENn(GND), .YL(
        \FCCC_0/GL1_INST/U0_RGB1_RGB14_rgbl_net_1 ), .YR(
        \FCCC_0/GL1_INST/U0_RGB1_RGB14_rgbr_net_1 ));
    INV_BA AFLSDF_INV_76 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_44_net_1 ), .Y(
        AFLSDF_INV_76_net_1));
    CFG2 #( .INIT(4'hD) )  \CoreGPIO_0/edge_neg_2_sqmuxa_8_i_o4_0_o2  
        (.A(\CoreGPIO_0/INTR_reg21 ), .B(\CoreGPIO_0.N_247 ), .Y(
        \CoreGPIO_0/N_248 ));
    CFG4 #( .INIT(16'h7530) )  
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_4[1]  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_12_[1]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/mem_4_[1]_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/N_504 ), .D(
        \reg_apb_wrp_0/reg16x8_0/N_495 ), .Y(
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_4[1]_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_44_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB5_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_5__1_sqmuxa ), .ALn(
        AFLSDF_INV_76_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(GND)
        , .Q(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_44_set_net_1 ));
    sdf_IOPAD_BI \FIC_MSS_0/MDDR_DQ_0_PAD/U_IOPAD  (.PAD(MDDR_DQ[0]), 
        .D(\FIC_MSS_0/DRAM_DQ_OUT_net_0[0] ), .E(
        \FIC_MSS_0/DRAM_DQ_OE_net_0[0] ), .Y(
        \FIC_MSS_0/MDDR_DQ_0_PAD_Y ));
    CFG4 #( .INIT(16'h0CAE) )  \CoreGPIO_0/PRDATA_iv_0_0_1[0]  (.A(
        \CoreGPIO_0/PRDATA_iv_0_0_a2_0_0[0]_net_1 ), .B(
        \CoreGPIO_0/INTR_reg[0] ), .C(\CoreGPIO_0.N_247 ), .D(
        \CoreGPIO_0.N_246 ), .Y(\CoreGPIO_0.PRDATA_iv_0_0_1[0] ));
    IP_INTERFACE \FCCC_0/CCC_INST/IP_INTERFACE_5  (.A(VCC), .B(VCC), 
        .C(VCC), .IPA(), .IPB(\FCCC_0/CCC_INST/NGMUX1_HOLD_N_net ), 
        .IPC(\FCCC_0/CCC_INST/PWDATA_net[3] ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_154_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_126_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_154_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_154_rs_net_1 ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_83  (.A(VCC), 
        .B(VCC), .C(VCC), .IPA(), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[24] ), .IPC());
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_15_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB11_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_5__1_sqmuxa ), .ALn(
        AFLSDF_INV_77_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(GND)
        , .Q(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_15_set_net_1 ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[0].REG_GEN.CONFIG_reg[0][6]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[6] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB11_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[0]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB1_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[0][6] ));
    CFG4 #( .INIT(16'hAC0F) )  
        \CoreGPIO_0/CONFIG_reg_o_2_31_am_RNO_0[5]  (.A(
        \CoreGPIO_0/CONFIG_reg[14][5] ), .B(
        \CoreGPIO_0/CONFIG_reg[30][5] ), .C(
        \CoreGPIO_0/CONFIG_reg_o_2_13_1_1[5] ), .D(
        \CoreAPB3_0_APBmslave3_PADDR[5] ), .Y(
        \CoreGPIO_0/CONFIG_reg_o_2_31_am_RNO_0[5]_net_1 ));
    INV_BA AFLSDF_INV_28 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_95_net_1 ), .Y(
        AFLSDF_INV_28_net_1));
    CFG4 #( .INIT(16'hA9FF) )  
        \CoreGPIO_0/xhdl1.GEN_BITS[26].APB_32.INTR_reg_347_0_o2_0_0[26]  
        (.A(\CoreGPIO_0/CONFIG_reg[26][7] ), .B(
        \CoreGPIO_0/CONFIG_reg[26][6] ), .C(
        \CoreGPIO_0/CONFIG_reg[26][5] ), .D(
        \CoreGPIO_0/CONFIG_reg[26][3] ), .Y(
        \CoreGPIO_0/INTR_reg_347_0_o2_0[26] ));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_62_set_RNIFAJG  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_62_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_254_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_15_rs[5] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_15_[5]_net_1 ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[6].REG_GEN.CONFIG_reg[6][2]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[2] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB14_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[6]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB4_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[6][2] ));
    INV_BA AFLSDF_INV_88 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_39_net_1 ), .Y(
        AFLSDF_INV_88_net_1));
    CFG4 #( .INIT(16'h7350) )  
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_3[7]  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_11_[7]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/mem_3_[7]_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/N_505 ), .D(
        \reg_apb_wrp_0/reg16x8_0/N_494 ), .Y(
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_3[7]_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_14_[3]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[3] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB7_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_14__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_243_i ), .ADn(VCC), .SLn(
        VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_14_rs[3] ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[5].gpin1[5]  (.D(\GPIO_IN_c[5] ), 
        .CLK(\FCCC_0/GL1_INST/U0_RGB1_RGB10_rgbr_net_1 ), .EN(VCC), 
        .ALn(\MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB0_rgbr_net_1 ), 
        .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/gpin1[5] ));
    CFG4 #( .INIT(16'h8000) )  
        \CoreGPIO_0/xhdl1.GEN_BITS[19].REG_GEN.CONFIG_reg[19]2_0_a4_0_a2  
        (.A(\CoreAPB3_0_APBmslave3_PADDR[3] ), .B(
        \CoreAPB3_0_APBmslave3_PADDR[2] ), .C(\CoreGPIO_0/N_598 ), .D(
        \CoreGPIO_0/N_606 ), .Y(\CoreGPIO_0/CONFIG_reg[19]2 ));
    CFG3 #( .INIT(8'hDF) )  \CoreGPIO_0/edge_pos_2_sqmuxa_2_i_0_0  (.A(
        \CoreGPIO_0/CONFIG_reg[6][3] ), .B(\CoreGPIO_0/N_689 ), .C(
        \CoreGPIO_0/N_248 ), .Y(\CoreGPIO_0/N_72 ));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_178_rs_RNIV1V51  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_42_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_178_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_5_rs[3] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_5_[3]_net_1 ));
    CFG3 #( .INIT(8'hF2) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_186  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_5_[7]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_490 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_186_i ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_243  (.A(VCC), 
        .B(GND), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[55] ), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/F_WSTRB_net[3] ), .IPC());
    CFG4 #( .INIT(16'hC5CA) )  
        \CoreGPIO_0/xhdl1.GEN_BITS[0].APB_32.INTR_reg_9_0_0_m2[0]  (.A(
        \CoreGPIO_0.xhdl1.GEN_BITS[0].gpin3[0] ), .B(
        \CoreGPIO_0/N_175 ), .C(\CoreGPIO_0/CONFIG_reg[0][6] ), .D(
        \CoreGPIO_0/CONFIG_reg[0][5] ), .Y(
        \CoreGPIO_0/INTR_reg_9_0_0_m2[0] ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_117_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB8_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_14__1_sqmuxa ), .ALn(
        AFLSDF_INV_78_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(GND)
        , .Q(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_117_set_net_1 ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_114  (.A(VCC), 
        .B(VCC), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/FAB_XDATAIN_net[6] ), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/FAB_VSTATUS_net[3] ), .IPC());
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_67_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB16_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_4__1_sqmuxa ), .ALn(
        AFLSDF_INV_79_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(GND)
        , .Q(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_67_set_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_240_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_112_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_240_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_240_rs_net_1 ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[28].REG_GEN.CONFIG_reg[28][1]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[1] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB14_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[28]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB4_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[28][1] ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[20].REG_GEN.CONFIG_reg[20][4]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[4] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB14_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[20]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB4_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[20][4] ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[5].REG_GEN.CONFIG_reg[5][2]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[2] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB14_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[5]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB4_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[5][2] ));
    CFG4 #( .INIT(16'h5410) )  \FIC_MSS_0/MSS_ADLIB_INST_RNO_14  (.A(
        \CoreAPB3_0_APBmslave3_PADDR[7] ), .B(
        \CoreAPB3_0_APBmslave3_PADDR[2] ), .C(
        \CONFIG_reg_o_2_31_am[3] ), .D(\CONFIG_reg_o_2_31_bm[3] ), .Y(
        \FIC_MSS_0/CoreAPB3_0_APBmslave5_PRDATA_m_0_1[3] ));
    sdf_IOPAD_BI \FIC_MSS_0/MDDR_DQ_11_PAD/U_IOPAD  (.PAD(MDDR_DQ[11]), 
        .D(\FIC_MSS_0/DRAM_DQ_OUT_net_0[11] ), .E(
        \FIC_MSS_0/DRAM_DQ_OE_net_0[11] ), .Y(
        \FIC_MSS_0/MDDR_DQ_11_PAD_Y ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[26].REG_GEN.CONFIG_reg[26][4]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[4] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB17_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[26]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB7_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[26][4] ));
    CFG4 #( .INIT(16'hCC0A) )  
        \CoreGPIO_0/xhdl1.GEN_BITS[0].APB_32.INTR_reg_9_0_0[0]  (.A(
        \CoreGPIO_0/INTR_reg[0] ), .B(\CoreGPIO_0/N_1575_tz ), .C(
        \CoreAPB3_0_APBmslave3_PWDATA[0] ), .D(\CoreGPIO_0/N_248 ), .Y(
        \CoreGPIO_0/INTR_reg_9[0] ));
    CFG4 #( .INIT(16'h0F35) )  
        \CoreGPIO_0/CONFIG_reg_o_2_31_bm_1_RNO_2[3]  (.A(
        \CoreGPIO_0/CONFIG_reg[1][3] ), .B(
        \CoreGPIO_0/CONFIG_reg[17][3] ), .C(
        \CoreAPB3_0_APBmslave3_PADDR[6] ), .D(
        \CoreAPB3_0_APBmslave3_PADDR[5] ), .Y(
        \CoreGPIO_0/CONFIG_reg_o_2_18_1[3] ));
    CFG3 #( .INIT(8'hF2) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_192  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_6_[2]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_493 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_192_i ));
    CFG2 #( .INIT(4'h7) )  \CoreGPIO_0/edge_both_2_sqmuxa_18_i  (.A(
        \CoreGPIO_0/N_248 ), .B(\CoreGPIO_0/CONFIG_reg[10][3] ), .Y(
        \CoreGPIO_0/N_184 ));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_7_[1]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[1] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB7_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_7__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_206_i ), .ADn(VCC), .SLn(
        VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_7_rs[1] ));
    CFG4 #( .INIT(16'h0F35) )  
        \CoreGPIO_0/CONFIG_reg_o_2_31_am_1_RNO_1[4]  (.A(
        \CoreGPIO_0/CONFIG_reg[4][4] ), .B(
        \CoreGPIO_0/CONFIG_reg[20][4] ), .C(
        \CoreAPB3_0_APBmslave3_PADDR[6] ), .D(
        \CoreAPB3_0_APBmslave3_PADDR[5] ), .Y(
        \CoreGPIO_0/CONFIG_reg_o_2_6_1[4] ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[2].REG_GEN.CONFIG_reg[2][7]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[7] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB17_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[2]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB7_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[2][7] ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_31_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB6_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_6__1_sqmuxa ), .ALn(
        AFLSDF_INV_80_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(GND)
        , .Q(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_31_set_net_1 ));
    CFG4 #( .INIT(16'hFF4F) )  \CoreGPIO_0/edge_both_2_sqmuxa_11_i_0  
        (.A(\CoreGPIO_0.N_247 ), .B(\CoreGPIO_0/INTR_reg21 ), .C(
        \CoreGPIO_0/CONFIG_reg[4][3] ), .D(\CoreGPIO_0/N_143_i ), .Y(
        \CoreGPIO_0/N_84 ));
    CFG3 #( .INIT(8'hF2) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_169  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_8_[5]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_499 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_169_i ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_213  (.A(VCC), 
        .B(GND), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[31] ), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/F_WID_HREADY01_net[1] ), .IPC());
    CFG2 #( .INIT(4'h4) )  \CoreGPIO_0/edge_neg_2_sqmuxa_7_i_a2  (.A(
        \CoreGPIO_0/gpin2[5] ), .B(
        \CoreGPIO_0.xhdl1.GEN_BITS[5].gpin3[5] ), .Y(
        \CoreGPIO_0/N_405 ));
    CFG4 #( .INIT(16'h0040) )  \FIC_MSS_0/MSS_ADLIB_INST_RNO_24  (.A(
        \xhdl1.GEN_BITS[0].APB_32.un5_PRDATA_o_0_a2_0_o2_x ), .B(
        CoreAPB3_0_APBmslave5_PSELx), .C(
        \CoreGPIO_0.xhdl1.GEN_BITS[4].APB_32.INTR_reg[4] ), .D(
        \CoreGPIO_0.RDATA_32.un12_PRDATA_o_0_o2_1 ), .Y(
        \FIC_MSS_0/CoreAPB3_0_APBmslave5_PRDATA_m_c_d[4] ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[27].REG_GEN.CONFIG_reg[27][4]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[4] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB10_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[27]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB0_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[27][4] ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_28  (.A(GND), 
        .B(GND), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[4] ), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[11] ), .IPC());
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_220_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_95_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_220_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_220_rs_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_50_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB10_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_3__1_sqmuxa ), .ALn(
        AFLSDF_INV_81_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(GND)
        , .Q(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_50_set_net_1 ));
    CFG4 #( .INIT(16'hFFFE) )  
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_13[3]  (.A(
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_7[3]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_5[3]_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_6[3]_net_1 ), .D(
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_4[3]_net_1 ), .Y(
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_13[3]_net_1 ));
    CFG2 #( .INIT(4'h7) )  \CoreGPIO_0/edge_both_2_sqmuxa_20_i  (.A(
        \CoreGPIO_0/N_248 ), .B(\CoreGPIO_0/CONFIG_reg[8][3] ), .Y(
        \CoreGPIO_0/edge_neg_2_sqmuxa_4_i_1 ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[9].REG_GEN.CONFIG_reg[9][0]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[0] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB16_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[9]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB6_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[9][0] ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[4].REG_GEN.CONFIG_reg[4][4]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[4] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB14_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[4]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB4_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[4][4] ));
    INV_BA AFLSDF_INV_117 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_98_net_1 ), .Y(
        AFLSDF_INV_117_net_1));
    IO_DIFF \FIC_MSS_0/MDDR_DQS_0_PAD/U_ION  (.YIN(GND));
    CFG4 #( .INIT(16'hEC00) )  \CoreAPB3_0/u_mux_p_to_b3/PRDATA[22]  (
        .A(\CoreGPIO_0.xhdl1.GEN_BITS[0].APB_32.GPOUT_reg9 ), .B(
        \CoreGPIO_0.N_542 ), .C(
        \CoreGPIO_0.xhdl1.GEN_BITS[22].APB_32.GPOUT_reg[22] ), .D(
        CoreAPB3_0_APBmslave5_PSELx), .Y(
        \FIC_MSS_0_FIC_0_APB_MASTER_PRDATA[22] ));
    CFG4 #( .INIT(16'h8F88) )  \FIC_MSS_0/MSS_ADLIB_INST_RNO_8  (.A(
        \CoreAPB3_0_APBmslave3_PRDATA[1] ), .B(
        CoreAPB3_0_APBmslave3_PSELx), .C(\CoreGPIO_0.N_247 ), .D(
        \FIC_MSS_0/CoreAPB3_0_APBmslave5_PRDATA_m_c_c_0[1] ), .Y(
        \FIC_MSS_0/CoreAPB3_0_APBmslave5_PRDATA_m_0_0[1] ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[11].REG_GEN.CONFIG_reg[11][3]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[3] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB9_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[11]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_YR ), .ADn(VCC), .SLn(
        VCC), .SD(GND), .LAT(GND), .Q(\CoreGPIO_0/CONFIG_reg[11][3] ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_282  (.A(VCC), 
        .B(VCC), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PADDR_net[5] ), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[9] ), .IPC());
    CFG3 #( .INIT(8'h20) )  
        \CoreGPIO_0/xhdl1.GEN_BITS[26].APB_32.edge_both_RNO[26]  (.A(
        \CoreGPIO_0/CONFIG_reg[26][3] ), .B(
        \CoreAPB3_0_APBmslave3_PWDATA[26] ), .C(
        \CoreGPIO_0/edge_pos[26] ), .Y(\CoreGPIO_0/N_106_i_0 ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[0].gpin1[0]  (.D(\GPIO_IN_c[0] ), 
        .CLK(\FCCC_0/GL1_INST/U0_RGB1_RGB9_rgbr_net_1 ), .EN(VCC), 
        .ALn(\MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_YR ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(GND), .Q(\CoreGPIO_0/gpin1[0] ));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_9_[0]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[0] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB13_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_9__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_175_i ), .ADn(VCC), .SLn(
        VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_9_rs[0] ));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_10_[1]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[1] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB1_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_10__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_193_i ), .ADn(VCC), .SLn(
        VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_10_rs[1] ));
    IOTRI_OB_EB \FIC_MSS_0/MDDR_BA_0_PAD/U_IOOUT  (.D(VCC), .E(VCC), 
        .DOUT(), .EOUT(\FIC_MSS_0/MDDR_BA_0_PAD/EOUT ));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_198_rs_RNIA7I5  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_39_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_198_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_6_rs[5] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_6_[5]_net_1 ));
    CFG3 #( .INIT(8'hB8) )  
        \CoreGPIO_0/xhdl1.GEN_BITS[4].APB_32.INTR_reg_61_0_m2_0[4]  (
        .A(\CoreGPIO_0/edge_neg[4] ), .B(\CoreGPIO_0/CONFIG_reg[4][5] )
        , .C(\CoreGPIO_0/edge_pos[4] ), .Y(\CoreGPIO_0/N_172 ));
    CFG2 #( .INIT(4'h8) )  \CoreGPIO_0/PRDATA_iv_0_0_a2_0_0[2]  (.A(
        \CoreAPB3_0_APBmslave3_PADDR[5] ), .B(
        \CoreGPIO_0/GPOUT_reg[2] ), .Y(
        \CoreGPIO_0/PRDATA_iv_0_0_a2_0_0[2]_net_1 ));
    CFG3 #( .INIT(8'hF2) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_160  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_3_[7]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_494 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_160_i ));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/mem_8__RNICUH51[0]  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_7_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_219_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_8_rs[0] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_8_[0]_net_1 ));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_182_rs_RNI06B41  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_46_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_182_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_5_rs[5] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_5_[5]_net_1 ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[5].APB_32.edge_pos[5]  (.D(
        \CoreGPIO_0/N_101 ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB10_rgbr_net_1 ), .EN(
        \CoreGPIO_0/N_70 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB0_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/edge_pos[5] ));
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_10  (
        .A(\reg_apb_wrp_0/reg16x8_0/mem_1_[0]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_502 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_10_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_10_[7]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[7] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB12_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_10__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_205_i ), .ADn(VCC), .SLn(
        VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_10_rs[7] ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_259  (.A(VCC), 
        .B(VCC), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[7] ), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[19] ), .IPC());
    IOBI_IB_OB_EB \FIC_MSS_0/MDDR_DQ_1_PAD/U_IOBI  (.D(VCC), .E(VCC), 
        .YIN(\FIC_MSS_0/MDDR_DQ_1_PAD/YIN ), .DOUT(), .EOUT(), .Y());
    CFG3 #( .INIT(8'h20) )  
        \CoreGPIO_0/xhdl1.GEN_BITS[30].APB_32.edge_both_RNO[30]  (.A(
        \CoreGPIO_0/CONFIG_reg[30][3] ), .B(
        \CoreAPB3_0_APBmslave3_PWDATA[30] ), .C(
        \CoreGPIO_0/edge_pos[30] ), .Y(\CoreGPIO_0/edge_neg_429[30] ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_96  (.A(VCC), 
        .B(VCC), .C(VCC), .IPA(\FIC_MSS_0/MSS_ADLIB_INST/CRSF_net ), 
        .IPB(), .IPC());
    CFG4 #( .INIT(16'hEFEE) )  
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_10[6]  (.A(
        \reg_apb_wrp_0/reg16x8_0/N_452 ), .B(
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_5[6]_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_4_[6]_net_1 ), .D(
        \reg_apb_wrp_0/reg16x8_0/N_504 ), .Y(
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_10[6]_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_14_[5]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[5] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB7_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_14__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_245_i ), .ADn(VCC), .SLn(
        VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_14_rs[5] ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[11].REG_GEN.CONFIG_reg[11][0]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[0] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB9_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[11]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_YR ), .ADn(VCC), .SLn(
        VCC), .SD(GND), .LAT(GND), .Q(\CoreGPIO_0/CONFIG_reg[11][0] ));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_81_set_RNIM74H  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_81_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_128_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_0_rs[1] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_0_[1]_net_1 ));
    CFG4 #( .INIT(16'h0F35) )  
        \CoreGPIO_0/CONFIG_reg_o_2_31_am_1_RNO_1[3]  (.A(
        \CoreGPIO_0/CONFIG_reg[4][3] ), .B(
        \CoreGPIO_0/CONFIG_reg[20][3] ), .C(
        \CoreAPB3_0_APBmslave3_PADDR[6] ), .D(
        \CoreAPB3_0_APBmslave3_PADDR[5] ), .Y(
        \CoreGPIO_0/CONFIG_reg_o_2_6_1[3] ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_180_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_44_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_180_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_180_rs_net_1 ));
    CFG4 #( .INIT(16'hA9FF) )  
        \CoreGPIO_0/xhdl1.GEN_BITS[31].APB_32.INTR_reg_412_0_o2_0_0[31]  
        (.A(\CoreGPIO_0/CONFIG_reg[31][7] ), .B(
        \CoreGPIO_0/CONFIG_reg[31][6] ), .C(
        \CoreGPIO_0/CONFIG_reg[31][5] ), .D(
        \CoreGPIO_0/CONFIG_reg[31][3] ), .Y(
        \CoreGPIO_0/INTR_reg_412_0_o2_0[31] ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_187  (.A(VCC), 
        .B(VCC), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/MMUART0_SCK_F2H_SCP_net ), .IPB(), 
        .IPC());
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_14_set_RNILPRT  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_14_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_138_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_1_rs[2] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_1_[2]_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_53_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB8_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_7__1_sqmuxa ), .ALn(
        AFLSDF_INV_82_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(GND)
        , .Q(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_53_set_net_1 ));
    CFG3 #( .INIT(8'hF2) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_165  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_4_[4]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_504 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_165_i ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[30].REG_GEN.CONFIG_reg[30][1]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[1] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB15_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[30]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB5_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[30][1] ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_2_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB12_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_4__1_sqmuxa ), .ALn(
        AFLSDF_INV_83_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(GND)
        , .Q(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_2_set_net_1 ));
    CFG2 #( .INIT(4'h2) )  
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_a3_13[2]  (.A(
        \reg_apb_wrp_0/reg16x8_0/N_499 ), .B(
        \reg_apb_wrp_0/reg16x8_0/mem_8_[2]_net_1 ), .Y(
        \reg_apb_wrp_0/reg16x8_0/N_400 ));
    IOBI_IB_OB_EB \FIC_MSS_0/MDDR_DQ_15_PAD/U_IOBI  (.D(VCC), .E(VCC), 
        .YIN(\FIC_MSS_0/MDDR_DQ_15_PAD/YIN ), .DOUT(), .EOUT(), .Y());
    CFG4 #( .INIT(16'h0F35) )  
        \CoreGPIO_0/CONFIG_reg_o_2_31_am_1_RNO_1[6]  (.A(
        \CoreGPIO_0/CONFIG_reg[4][6] ), .B(
        \CoreGPIO_0/CONFIG_reg[20][6] ), .C(
        \CoreAPB3_0_APBmslave3_PADDR[6] ), .D(
        \CoreAPB3_0_APBmslave3_PADDR[5] ), .Y(
        \CoreGPIO_0/CONFIG_reg_o_2_6_1[6] ));
    CFG3 #( .INIT(8'hF2) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_152  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_3_[0]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_494 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_152_i ));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_14_[4]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[4] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB9_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_14__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_244_i ), .ADn(VCC), .SLn(
        VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_14_rs[4] ));
    CFG4 #( .INIT(16'h2000) )  
        \CoreGPIO_0/xhdl1.GEN_BITS[18].REG_GEN.CONFIG_reg[18]2_0_a4_0_a2  
        (.A(\CoreAPB3_0_APBmslave3_PADDR[3] ), .B(
        \CoreAPB3_0_APBmslave3_PADDR[2] ), .C(\CoreGPIO_0/N_598 ), .D(
        \CoreGPIO_0/N_606 ), .Y(\CoreGPIO_0/CONFIG_reg[18]2 ));
    CFG2 #( .INIT(4'h2) )  
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_a3_3[0]  (.A(
        \reg_apb_wrp_0/reg16x8_0/N_500 ), .B(
        \reg_apb_wrp_0/reg16x8_0/mem_13_[0]_net_1 ), .Y(
        \reg_apb_wrp_0/reg16x8_0/N_358 ));
    CFG4 #( .INIT(16'hAC0F) )  
        \CoreGPIO_0/CONFIG_reg_o_2_31_bm_RNO[6]  (.A(
        \CoreGPIO_0/CONFIG_reg[11][6] ), .B(
        \CoreGPIO_0/CONFIG_reg[27][6] ), .C(
        \CoreGPIO_0/CONFIG_reg_o_2_25_1_1[6] ), .D(
        \CoreAPB3_0_APBmslave3_PADDR[5] ), .Y(
        \CoreGPIO_0/CONFIG_reg_o_2_31_bm_RNO[6]_net_1 ));
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_119  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_14_[7]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_503 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_119_net_1 ));
    CFG2 #( .INIT(4'h4) )  \CoreGPIO_0/PRDATA_0_iv_0_a2_0[29]  (.A(
        \CoreGPIO_0.N_247 ), .B(\CoreGPIO_0/INTR_reg[29] ), .Y(
        \CoreGPIO_0.N_528 ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[3].APB_32.GPOUT_reg[3]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[3] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB10_rgbr_net_1 ), .EN(
        \CoreGPIO_0/GPOUT_reg_0_sqmuxa ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB0_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/GPOUT_reg[3] ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_29_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB14_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_6__1_sqmuxa ), .ALn(
        AFLSDF_INV_84_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(GND)
        , .Q(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_29_set_net_1 ));
    sdf_IOPAD_BI \FIC_MSS_0/MDDR_DQ_10_PAD/U_IOPAD  (.PAD(MDDR_DQ[10]), 
        .D(\FIC_MSS_0/DRAM_DQ_OUT_net_0[10] ), .E(
        \FIC_MSS_0/DRAM_DQ_OE_net_0[10] ), .Y(
        \FIC_MSS_0/MDDR_DQ_10_PAD_Y ));
    sdf_IOPAD_TRI \FIC_MSS_0/MDDR_DQS_TMATCH_0_OUT_PAD/U_IOPAD  (.PAD(
        MDDR_DQS_TMATCH_0_OUT), .D(
        \FIC_MSS_0/DRAM_FIFO_WE_OUT_net_0[0] ), .E(
        \FIC_MSS_0/MDDR_DQS_TMATCH_0_OUT_PAD/EOUT ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_105_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB9_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_13__1_sqmuxa ), .ALn(
        AFLSDF_INV_85_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(GND)
        , .Q(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_105_set_net_1 ));
    INV_BA AFLSDF_INV_68 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_100_net_1 ), .Y(
        AFLSDF_INV_68_net_1));
    CFG4 #( .INIT(16'h330A) )  
        \CoreGPIO_0/xhdl1.GEN_BITS[21].APB_32.INTR_reg_282_0[21]  (.A(
        \CoreGPIO_0/INTR_reg[21] ), .B(
        \CoreGPIO_0/INTR_reg_282_0_o2_1[21] ), .C(
        \CoreAPB3_0_APBmslave3_PWDATA[21] ), .D(\CoreGPIO_0/N_248 ), 
        .Y(\CoreGPIO_0/INTR_reg_282[21] ));
    IP_INTERFACE \FCCC_0/CCC_INST/IP_INTERFACE_7  (.A(VCC), .B(VCC), 
        .C(VCC), .IPA(\FCCC_0/CCC_INST/CLK3_net ), .IPB(), .IPC(
        \FCCC_0/CCC_INST/PWDATA_net[5] ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[6].gpin3[6]  (.D(
        \CoreGPIO_0/gpin2[6] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB12_rgbr_net_1 ), .EN(VCC), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB2_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0.xhdl1.GEN_BITS[6].gpin3[6] ));
    CFG4 #( .INIT(16'hA9FF) )  
        \CoreGPIO_0/xhdl1.GEN_BITS[30].APB_32.INTR_reg_399_0_o2_0_0[30]  
        (.A(\CoreGPIO_0/CONFIG_reg[30][7] ), .B(
        \CoreGPIO_0/CONFIG_reg[30][6] ), .C(
        \CoreGPIO_0/CONFIG_reg[30][5] ), .D(
        \CoreGPIO_0/CONFIG_reg[30][3] ), .Y(
        \CoreGPIO_0/INTR_reg_399_0_o2_0[30] ));
    CFG4 #( .INIT(16'h0F35) )  
        \CoreGPIO_0/CONFIG_reg_o_2_31_bm_1_RNO_1[7]  (.A(
        \CoreGPIO_0/CONFIG_reg[5][7] ), .B(
        \CoreGPIO_0/CONFIG_reg[21][7] ), .C(
        \CoreAPB3_0_APBmslave3_PADDR[6] ), .D(
        \CoreAPB3_0_APBmslave3_PADDR[5] ), .Y(
        \CoreGPIO_0/CONFIG_reg_o_2_21_1[7] ));
    sdf_IOPAD_TRI \FIC_MSS_0/MDDR_ADDR_1_PAD/U_IOPAD  (.PAD(
        MDDR_ADDR[1]), .D(\FIC_MSS_0/DRAM_ADDR_net_0[1] ), .E(
        \FIC_MSS_0/MDDR_ADDR_1_PAD/EOUT ));
    sdf_IOPAD_TRI \FIC_MSS_0/MDDR_ADDR_11_PAD/U_IOPAD  (.PAD(
        MDDR_ADDR[11]), .D(\FIC_MSS_0/DRAM_ADDR_net_0[11] ), .E(
        \FIC_MSS_0/MDDR_ADDR_11_PAD/EOUT ));
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_48  (
        .A(\reg_apb_wrp_0/reg16x8_0/mem_3_[3]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_494 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_48_net_1 ));
    CFG4 #( .INIT(16'hEFEE) )  
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_11[6]  (.A(
        \reg_apb_wrp_0/reg16x8_0/N_460 ), .B(
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_7[6]_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_0_[6]_net_1 ), .D(
        \reg_apb_wrp_0/reg16x8_0/N_496 ), .Y(
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_11[6]_net_1 ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[19].REG_GEN.CONFIG_reg[19][7]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[7] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB9_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[19]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_YR ), .ADn(VCC), .SLn(
        VCC), .SD(GND), .LAT(GND), .Q(\CoreGPIO_0/CONFIG_reg[19][7] ));
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_110  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_13_[6]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_500 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_110_net_1 ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[20].APB_32.INTR_reg[20]  (.D(
        \CoreGPIO_0/INTR_reg_269[20] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB13_rgbr_net_1 ), .EN(VCC), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB3_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/INTR_reg[20] ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[7].REG_GEN.CONFIG_reg[7][5]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[5] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB10_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[7]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB0_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[7][5] ));
    CFG4 #( .INIT(16'hF2F3) )  
        \CoreGPIO_0/xhdl1.GEN_BITS[31].APB_32.INTR_reg_412_0_o2_1_0[31]  
        (.A(\CoreGPIO_0/CONFIG_reg[31][6] ), .B(
        \CoreGPIO_0/edge_pos[31] ), .C(
        \CoreGPIO_0/INTR_reg_412_0_o2_0[31] ), .D(
        \CoreGPIO_0/CONFIG_reg[31][5] ), .Y(
        \CoreGPIO_0/INTR_reg_412_0_o2_1[31] ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[14].APB_32.INTR_reg[14]  (.D(
        \CoreGPIO_0/INTR_reg_191[14] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB13_rgbr_net_1 ), .EN(VCC), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB3_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/INTR_reg[14] ));
    CFG4 #( .INIT(16'h330A) )  
        \CoreGPIO_0/xhdl1.GEN_BITS[14].APB_32.INTR_reg_191_0[14]  (.A(
        \CoreGPIO_0/INTR_reg[14] ), .B(
        \CoreGPIO_0/INTR_reg_191_0_o2_1[14] ), .C(
        \CoreAPB3_0_APBmslave3_PWDATA[14] ), .D(\CoreGPIO_0/N_248 ), 
        .Y(\CoreGPIO_0/INTR_reg_191[14] ));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_173_rs_RNI3EQN  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_71_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_173_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_8_rs[7] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_8_[7]_net_1 ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_158  (.A(VCC), 
        .B(VCC), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/MGPIO10A_F2H_GPIN_net ), .IPB(), 
        .IPC());
    CFG3 #( .INIT(8'hF2) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_172  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_5_[0]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_490 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_172_i ));
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_115  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_14_[3]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_503 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_115_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_4_[4]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[4] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB11_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_4__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_165_i ), .ADn(VCC), .SLn(
        VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_4_rs[4] ));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_109_set_RNI0KRF  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_109_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_237_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_13_rs[5] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_13_[5]_net_1 ));
    CFG4 #( .INIT(16'h0F35) )  
        \CoreGPIO_0/CONFIG_reg_o_2_31_bm_1_RNO_1[2]  (.A(
        \CoreGPIO_0/CONFIG_reg[5][2] ), .B(
        \CoreGPIO_0/CONFIG_reg[21][2] ), .C(
        \CoreAPB3_0_APBmslave3_PADDR[6] ), .D(
        \CoreAPB3_0_APBmslave3_PADDR[5] ), .Y(
        \CoreGPIO_0/CONFIG_reg_o_2_21_1[2] ));
    CFG4 #( .INIT(16'hAC0F) )  
        \CoreGPIO_0/CONFIG_reg_o_2_31_bm_1_RNO_0[7]  (.A(
        \CoreGPIO_0/CONFIG_reg[9][7] ), .B(
        \CoreGPIO_0/CONFIG_reg[25][7] ), .C(
        \CoreGPIO_0/CONFIG_reg_o_2_18_1[7] ), .D(
        \CoreAPB3_0_APBmslave3_PADDR[5] ), .Y(
        \CoreGPIO_0/CONFIG_reg_o_2_31_bm_1_RNO_0[7]_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_60_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB5_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_15__1_sqmuxa ), .ALn(
        AFLSDF_INV_86_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(GND)
        , .Q(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_60_set_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_10_[6]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[6] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB13_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_10__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_203_i ), .ADn(VCC), .SLn(
        VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_10_rs[6] ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_207_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_88_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_207_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_207_rs_net_1 ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_170  (.A(VCC), 
        .B(VCC), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/MMUART1_RI_F2H_SCP_net ), .IPB(), 
        .IPC());
    RGB \FCCC_0/GL1_INST/U0_RGB1_RGB17  (.An(
        \FCCC_0/GL1_INST/U0_YNn_GSouth ), .ENn(GND), .YL(
        \FCCC_0/GL1_INST/U0_RGB1_RGB17_rgbl_net_1 ), .YR(
        \FCCC_0/GL1_INST/U0_RGB1_RGB17_rgbr_net_1 ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[17].REG_GEN.CONFIG_reg[17][2]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[2] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB16_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[17]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB6_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[17][2] ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_151_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_120_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_151_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_151_rs_net_1 ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_276  (.A(VCC), 
        .B(VCC), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[0] ), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[3] ), .IPC(
        \FIC_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[15] ));
    CFG4 #( .INIT(16'h0400) )  
        \reg_apb_wrp_0/reg16x8_0/WRITE_GEN.mem_6__2_i_a2[6]  (.A(
        \CoreAPB3_0_APBmslave3_PADDR[3] ), .B(
        \CoreAPB3_0_APBmslave3_PADDR[2] ), .C(
        \CoreAPB3_0_APBmslave3_PADDR[0] ), .D(
        \CoreAPB3_0_APBmslave3_PADDR[1] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/N_493 ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_33  (.A(GND), 
        .B(GND), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[9] ), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[16] ), .IPC());
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[8].REG_GEN.CONFIG_reg[8][2]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[2] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB15_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[8]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB5_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[8][2] ));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_1_[1]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[1] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB14_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_1__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_137_i ), .ADn(VCC), .SLn(
        VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_1_rs[1] ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_80  (.A(VCC), 
        .B(VCC), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[14] ), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[21] ), .IPC());
    CFG4 #( .INIT(16'h8000) )  
        \CoreGPIO_0/xhdl1.GEN_BITS[27].REG_GEN.CONFIG_reg[27]2_0_a4_0_a2  
        (.A(\CoreAPB3_0_APBmslave3_PADDR[3] ), .B(
        \CoreAPB3_0_APBmslave3_PADDR[2] ), .C(\CoreGPIO_0/N_598 ), .D(
        \CoreGPIO_0/N_610 ), .Y(\CoreGPIO_0/CONFIG_reg[27]2 ));
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_4  (
        .A(\reg_apb_wrp_0/reg16x8_0/mem_4_[2]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_504 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_4_net_1 ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_240  (.A(VCC), 
        .B(GND), .C(GND), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[52] ), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/F_WSTRB_net[0] ), .IPC(
        \FIC_MSS_0/MSS_ADLIB_INST/F_WVALID_net ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_152_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_122_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_152_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_152_rs_net_1 ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[14].APB_32.GPOUT_reg[14]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[14] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB13_rgbr_net_1 ), .EN(
        \CoreGPIO_0/GPOUT_reg_0_sqmuxa ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB3_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0.xhdl1.GEN_BITS[14].APB_32.GPOUT_reg[14] ));
    CFG4 #( .INIT(16'h7530) )  
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_7[6]  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_10_[6]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/mem_2_[6]_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/N_501 ), .D(
        \reg_apb_wrp_0/reg16x8_0/N_491 ), .Y(
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_7[6]_net_1 ));
    CFG4 #( .INIT(16'hF2F3) )  
        \CoreGPIO_0/xhdl1.GEN_BITS[27].APB_32.INTR_reg_360_0_o2_1_0[27]  
        (.A(\CoreGPIO_0/CONFIG_reg[27][6] ), .B(
        \CoreGPIO_0/edge_neg[27] ), .C(
        \CoreGPIO_0/INTR_reg_360_0_o2_0[27] ), .D(
        \CoreGPIO_0/CONFIG_reg[27][5] ), .Y(
        \CoreGPIO_0/INTR_reg_360_0_o2_1[27] ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[24].APB_32.edge_both[24]  (.D(
        \CoreGPIO_0/N_100_i_0 ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB9_rgbr_net_1 ), .EN(
        \CoreGPIO_0/N_155 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_YR ), .ADn(VCC), .SLn(
        VCC), .SD(GND), .LAT(GND), .Q(\CoreGPIO_0/edge_pos[24] ));
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_107  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_13_[3]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_500 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_107_net_1 ));
    CFG3 #( .INIT(8'hF2) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_205  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_10_[7]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_491 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_205_i ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_247  (.A(VCC), 
        .B(GND), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[59] ), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/F_WSTRB_net[7] ), .IPC());
    CFG4 #( .INIT(16'hAC0F) )  
        \CoreGPIO_0/CONFIG_reg_o_2_31_am_RNO_0[6]  (.A(
        \CoreGPIO_0/CONFIG_reg[14][6] ), .B(
        \CoreGPIO_0/CONFIG_reg[30][6] ), .C(
        \CoreGPIO_0/CONFIG_reg_o_2_13_1_1[6] ), .D(
        \CoreAPB3_0_APBmslave3_PADDR[5] ), .Y(
        \CoreGPIO_0/CONFIG_reg_o_2_31_am_RNO_0[6]_net_1 ));
    CFG4 #( .INIT(16'hAC0F) )  
        \CoreGPIO_0/CONFIG_reg_o_2_31_bm_1_RNO_0[6]  (.A(
        \CoreGPIO_0/CONFIG_reg[9][6] ), .B(
        \CoreGPIO_0/CONFIG_reg[25][6] ), .C(
        \CoreGPIO_0/CONFIG_reg_o_2_18_1[6] ), .D(
        \CoreAPB3_0_APBmslave3_PADDR[5] ), .Y(
        \CoreGPIO_0/CONFIG_reg_o_2_31_bm_1_RNO_0[6]_net_1 ));
    INV_BA AFLSDF_INV_20 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_83_net_1 ), .Y(
        AFLSDF_INV_20_net_1));
    CFG2 #( .INIT(4'h4) )  \CoreAPB3_0/iPSELS_1_0[5]  (.A(
        \FIC_MSS_0_FIC_0_APB_MASTER_PADDR[29] ), .B(
        \FIC_MSS_0_FIC_0_APB_MASTER_PADDR[30] ), .Y(
        \CoreAPB3_0/iPSELS_1[5] ));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/mem_14__RNISAMI[4]  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_116_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_244_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_14_rs[4] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_14_[4]_net_1 ));
    INV_BA AFLSDF_INV_80 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_31_net_1 ), .Y(
        AFLSDF_INV_80_net_1));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_6_[6]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[6] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB13_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_6__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_200_i ), .ADn(VCC), .SLn(
        VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_6_rs[6] ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_63_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB6_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_15__1_sqmuxa ), .ALn(
        AFLSDF_INV_87_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(GND)
        , .Q(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_63_set_net_1 ));
    CFG4 #( .INIT(16'hF2F3) )  
        \CoreGPIO_0/xhdl1.GEN_BITS[26].APB_32.INTR_reg_347_0_o2_1_0[26]  
        (.A(\CoreGPIO_0/CONFIG_reg[26][6] ), .B(
        \CoreGPIO_0/edge_pos[26] ), .C(
        \CoreGPIO_0/INTR_reg_347_0_o2_0[26] ), .D(
        \CoreGPIO_0/CONFIG_reg[26][5] ), .Y(
        \CoreGPIO_0/INTR_reg_347_0_o2_1[26] ));
    CFG4 #( .INIT(16'hEC00) )  \CoreAPB3_0/u_mux_p_to_b3/PRDATA[27]  (
        .A(\CoreGPIO_0.xhdl1.GEN_BITS[0].APB_32.GPOUT_reg9 ), .B(
        \CoreGPIO_0.N_532 ), .C(
        \CoreGPIO_0.xhdl1.GEN_BITS[27].APB_32.GPOUT_reg[27] ), .D(
        CoreAPB3_0_APBmslave5_PSELx), .Y(
        \FIC_MSS_0_FIC_0_APB_MASTER_PRDATA[27] ));
    SLE \reg_apb_wrp_0/reg16x8_0/data_out[0]  (.D(
        \reg_apb_wrp_0/reg16x8_0/temp_data[0]_net_1 ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB13_rgbr_net_1 ), .EN(VCC), .ALn(
        VCC), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreAPB3_0_APBmslave3_PRDATA[0] ));
    IOOUTFF_BYPASS \GPIO_OUT_obuf[0]/U0/U_IOOUTFF  (.A(
        \GPIO_OUT_obuf[0]/U0/DOUT1 ), .Y(\GPIO_OUT_obuf[0]/U0/DOUT ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_154  (.A(VCC), 
        .B(VCC), .C(VCC), .IPA(), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/SPI0_SS0_F2H_SCP_net ), .IPC());
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_167_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_68_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_167_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_167_rs_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_140_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_41_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_140_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_140_rs_net_1 ));
    CFG3 #( .INIT(8'hF2) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_199  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_10_[4]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_491 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_199_i ));
    CFG3 #( .INIT(8'h26) )  \reg_apb_wrp_0/fsm_ns_1_0_.m4  (.A(
        \reg_apb_wrp_0/fsm[1]_net_1 ), .B(\reg_apb_wrp_0/fsm[0]_net_1 )
        , .C(CoreAPB3_0_APBmslave3_PWRITE), .Y(
        \reg_apb_wrp_0/fsm_ns[1] ));
    IOINFF_BYPASS \FIC_MSS_0/MDDR_DQ_3_PAD/U_IOINFF  (.A(
        \FIC_MSS_0/MDDR_DQ_3_PAD_Y ), .Y(\FIC_MSS_0/MDDR_DQ_3_PAD/YIN )
        );
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[17].REG_GEN.CONFIG_reg[17][6]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[6] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB15_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[17]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB5_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[17][6] ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_237_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_109_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_237_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_237_rs_net_1 ));
    CFG2 #( .INIT(4'h8) )  
        \reg_apb_wrp_0/reg16x8_0/mem_0__1_sqmuxa_0_a2_0_a3  (.A(
        \reg_apb_wrp_0/reg16x8_0/N_496 ), .B(
        \reg_apb_wrp_0/wr_enable_net_1 ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_0__1_sqmuxa ));
    CFG4 #( .INIT(16'hF2F3) )  
        \CoreGPIO_0/xhdl1.GEN_BITS[12].APB_32.INTR_reg_165_0_o2_1_0[12]  
        (.A(\CoreGPIO_0/CONFIG_reg[12][6] ), .B(
        \CoreGPIO_0/edge_neg[12] ), .C(
        \CoreGPIO_0/INTR_reg_165_0_o2_0[12] ), .D(
        \CoreGPIO_0/CONFIG_reg[12][5] ), .Y(
        \CoreGPIO_0/INTR_reg_165_0_o2_1[12] ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_210  (.A(VCC), 
        .B(GND), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[28] ), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/F_AWLOCK_HMASTLOCK0_net[0] ), .IPC());
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_265  (.A(VCC), 
        .B(GND), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[25] ), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/F_ARBURST_HTRANS1_net[1] ), .IPC(
        \FIC_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWRITE_net ));
    sdf_IOPAD_TRI \FIC_MSS_0/MDDR_ODT_PAD/U_IOPAD  (.PAD(MDDR_ODT), .D(
        \FIC_MSS_0/MSS_ADLIB_INST_DRAM_ODT ), .E(
        \FIC_MSS_0/MDDR_ODT_PAD/EOUT ));
    sdf_IOPAD_TRI \FIC_MSS_0/MDDR_ADDR_7_PAD/U_IOPAD  (.PAD(
        MDDR_ADDR[7]), .D(\FIC_MSS_0/DRAM_ADDR_net_0[7] ), .E(
        \FIC_MSS_0/MDDR_ADDR_7_PAD/EOUT ));
    INV_BA AFLSDF_INV_93 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_27_net_1 ), .Y(
        AFLSDF_INV_93_net_1));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_39_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB11_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_6__1_sqmuxa ), .ALn(
        AFLSDF_INV_88_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(GND)
        , .Q(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_39_set_net_1 ));
    CFG3 #( .INIT(8'hF2) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_206  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_7_[1]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_498 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_206_i ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_131  (.A(VCC), 
        .B(GND), .C(VCC), .IPA(), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[13] ), .IPC());
    CFG3 #( .INIT(8'hB8) )  
        \CoreGPIO_0/xhdl1.GEN_BITS[1].APB_32.INTR_reg_22_0_m2_0[1]  (
        .A(\CoreGPIO_0/edge_neg[1] ), .B(\CoreGPIO_0/CONFIG_reg[1][5] )
        , .C(\CoreGPIO_0/edge_pos[1] ), .Y(\CoreGPIO_0/N_174 ));
    CFG2 #( .INIT(4'h7) )  \CoreGPIO_0/edge_both_2_sqmuxa_5_i  (.A(
        \CoreGPIO_0/N_248 ), .B(\CoreGPIO_0/CONFIG_reg[14][3] ), .Y(
        \CoreGPIO_0/edge_pos_2_sqmuxa_8_i_1 ));
    sdf_IOPADN_TRI \FIC_MSS_0/MDDR_CLK_PAD/U_IOPADN  (.PAD_P(
        MDDR_CLK_N), .OIN_P(\FIC_MSS_0/MSS_ADLIB_INST_DRAM_CLK ), 
        .EIN_P(VCC));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_217  (.A(VCC), 
        .B(VCC), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[1] ), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[13] ), .IPC(
        \FIC_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[25] ));
    CFG4 #( .INIT(16'h4000) )  
        \CoreGPIO_0/xhdl1.GEN_BITS[6].REG_GEN.CONFIG_reg[6]2_0_a4_0_a2  
        (.A(\CoreAPB3_0_APBmslave3_PADDR[2] ), .B(
        \CoreAPB3_0_APBmslave3_PADDR[3] ), .C(\CoreGPIO_0/N_603 ), .D(
        \CoreGPIO_0/N_604 ), .Y(\CoreGPIO_0/CONFIG_reg[6]2 ));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_73_set_RNI40PO  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_73_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_177_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_9_rs[1] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_9_[1]_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_243_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_115_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_243_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_243_rs_net_1 ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[10].APB_32.GPOUT_reg[10]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[10] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB16_rgbr_net_1 ), .EN(
        \CoreGPIO_0/GPOUT_reg_0_sqmuxa ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB6_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/GPOUT_reg[10] ));
    CFG3 #( .INIT(8'hF2) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_190  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_6_[1]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_493 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_190_i ));
    CFG4 #( .INIT(16'hAA08) )  
        \CoreGPIO_0/xhdl1.GEN_BITS[1].APB_32.edge_pos_23_iv_i_0[1]  (
        .A(\CoreGPIO_0/CONFIG_reg[1][3] ), .B(\CoreGPIO_0/edge_pos[1] )
        , .C(\CoreAPB3_0_APBmslave3_PWDATA[1] ), .D(\CoreGPIO_0/N_400 )
        , .Y(\CoreGPIO_0/N_107 ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_253  (.A(VCC), 
        .B(VCC), .C(GND), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[1] ), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[13] ), .IPC(
        \FIC_MSS_0/MSS_ADLIB_INST/F_ARSIZE_HSIZE1_net[1] ));
    INV_BA AFLSDF_INV_96 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_net_1 ), .Y(
        AFLSDF_INV_96_net_1));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_162  (.A(VCC), 
        .B(VCC), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/MGPIO12A_F2H_GPIN_net ), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/MGPIO15A_F2H_GPIN_net ), .IPC());
    CFG4 #( .INIT(16'h2000) )  
        \CoreGPIO_0/xhdl1.GEN_BITS[30].REG_GEN.CONFIG_reg[30]2_0_a4_0_a2  
        (.A(\CoreAPB3_0_APBmslave3_PADDR[3] ), .B(
        \CoreAPB3_0_APBmslave3_PADDR[2] ), .C(\CoreGPIO_0/N_598 ), .D(
        \CoreGPIO_0/N_605 ), .Y(\CoreGPIO_0/CONFIG_reg[30]2 ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_62  (.A(GND), 
        .B(VCC), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[23] ), .IPB(), .IPC()
        );
    IOBI_IB_OB_EB \FIC_MSS_0/MDDR_DQ_8_PAD/U_IOBI  (.D(VCC), .E(VCC), 
        .YIN(\FIC_MSS_0/MDDR_DQ_8_PAD/YIN ), .DOUT(), .EOUT(), .Y());
    CFG3 #( .INIT(8'hF2) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_195  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_10_[2]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_491 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_195_i ));
    CFG4 #( .INIT(16'hFF4F) )  \CoreGPIO_0/edge_both_2_sqmuxa_15_i_0  
        (.A(\CoreGPIO_0.N_247 ), .B(\CoreGPIO_0/INTR_reg21 ), .C(
        \CoreGPIO_0/CONFIG_reg[0][3] ), .D(\CoreGPIO_0/N_141_i ), .Y(
        \CoreGPIO_0/N_80 ));
    sdf_IOPAD_TRI \FIC_MSS_0/MDDR_CKE_PAD/U_IOPAD  (.PAD(MDDR_CKE), .D(
        \FIC_MSS_0/MSS_ADLIB_INST_DRAM_CKE ), .E(
        \FIC_MSS_0/MDDR_CKE_PAD/EOUT ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[1].REG_GEN.CONFIG_reg[1][2]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[2] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB16_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[1]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB6_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[1][2] ));
    IOOUTFF_BYPASS \GPIO_OUT_obuf[6]/U0/U_IOOUTFF  (.A(
        \GPIO_OUT_obuf[6]/U0/DOUT1 ), .Y(\GPIO_OUT_obuf[6]/U0/DOUT ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_274  (.A(GND), 
        .B(VCC), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/F_ARLEN_HBURST1_net[2] ), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/CLK_MDDR_APB_net ), .IPC());
    sdf_IOPAD_BI \FIC_MSS_0/MDDR_DQ_5_PAD/U_IOPAD  (.PAD(MDDR_DQ[5]), 
        .D(\FIC_MSS_0/DRAM_DQ_OUT_net_0[5] ), .E(
        \FIC_MSS_0/DRAM_DQ_OE_net_0[5] ), .Y(
        \FIC_MSS_0/MDDR_DQ_5_PAD_Y ));
    INV_BA AFLSDF_INV_125 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_22_net_1 ), .Y(
        AFLSDF_INV_125_net_1));
    CFG4 #( .INIT(16'hAA08) )  
        \CoreGPIO_0/xhdl1.GEN_BITS[0].APB_32.edge_pos_9_iv_i_0[0]  (.A(
        \CoreGPIO_0/CONFIG_reg[0][3] ), .B(\CoreGPIO_0/edge_pos[0] ), 
        .C(\CoreAPB3_0_APBmslave3_PWDATA[0] ), .D(\CoreGPIO_0/N_402 ), 
        .Y(\CoreGPIO_0/N_109 ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_223_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_64_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_223_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_223_rs_net_1 ));
    CFG4 #( .INIT(16'hAC0F) )  
        \CoreGPIO_0/CONFIG_reg_o_2_31_am_1_RNO_0[1]  (.A(
        \CoreGPIO_0/CONFIG_reg[8][1] ), .B(
        \CoreGPIO_0/CONFIG_reg[24][1] ), .C(
        \CoreGPIO_0/CONFIG_reg_o_2_3_1[1] ), .D(
        \CoreAPB3_0_APBmslave3_PADDR[5] ), .Y(
        \CoreGPIO_0/CONFIG_reg_o_2_31_am_1_RNO_0[1]_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_96_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB2_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_10__1_sqmuxa ), .ALn(
        AFLSDF_INV_89_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(GND)
        , .Q(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_96_set_net_1 ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[17].APB_32.GPOUT_reg[17]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[17] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB14_rgbr_net_1 ), .EN(
        \CoreGPIO_0/GPOUT_reg_0_sqmuxa ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB4_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0.xhdl1.GEN_BITS[17].APB_32.GPOUT_reg[17] ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_114_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB8_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_14__1_sqmuxa ), .ALn(
        AFLSDF_INV_90_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(GND)
        , .Q(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_114_set_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_4_[2]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[2] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB11_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_4__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_163_i ), .ADn(VCC), .SLn(
        VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_4_rs[2] ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_205_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_100_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_205_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_205_rs_net_1 ));
    CFG3 #( .INIT(8'hF2) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_136  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_1_[0]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_502 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_136_i ));
    CFG4 #( .INIT(16'hAC0F) )  
        \CoreGPIO_0/CONFIG_reg_o_2_31_bm_RNO_0[7]  (.A(
        \CoreGPIO_0/CONFIG_reg[15][7] ), .B(
        \CoreGPIO_0/CONFIG_reg[31][7] ), .C(
        \CoreGPIO_0/CONFIG_reg_o_2_28_1_1[7] ), .D(
        \CoreAPB3_0_APBmslave3_PADDR[5] ), .Y(
        \CoreGPIO_0/CONFIG_reg_o_2_31_bm_RNO_0[7]_net_1 ));
    CFG3 #( .INIT(8'hF2) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_159  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_3_[6]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_494 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_159_i ));
    IOINFF_BYPASS \FIC_MSS_0/MDDR_DQ_12_PAD/U_IOINFF  (.A(
        \FIC_MSS_0/MDDR_DQ_12_PAD_Y ), .Y(
        \FIC_MSS_0/MDDR_DQ_12_PAD/YIN ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_133_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_86_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_133_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_133_rs_net_1 ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_7  (.A(
        \FIC_MSS_0/FIC_MSS_0_FIC_0_APB_MASTER_PRDATA[5] ), .B(
        \FIC_MSS_0_FIC_0_APB_MASTER_PRDATA[12] ), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[5] ), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[12] ), .IPC());
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_78_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB16_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_9__1_sqmuxa ), .ALn(
        AFLSDF_INV_91_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(GND)
        , .Q(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_78_set_net_1 ));
    INV_BA AFLSDF_INV_32 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_55_net_1 ), .Y(
        AFLSDF_INV_32_net_1));
    INV_BA AFLSDF_INV_101 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_103_net_1 ), .Y(
        AFLSDF_INV_101_net_1));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[31].APB_32.edge_both[31]  (.D(
        \CoreGPIO_0/edge_neg_443[31] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB10_rgbr_net_1 ), .EN(
        \CoreGPIO_0/edge_pos_2_sqmuxa_19_i_1 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB0_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/edge_pos[31] ));
    CFG2 #( .INIT(4'h2) )  
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_a3_11[6]  (.A(
        \reg_apb_wrp_0/reg16x8_0/N_492 ), .B(
        \reg_apb_wrp_0/reg16x8_0/mem_9_[6]_net_1 ), .Y(
        \reg_apb_wrp_0/reg16x8_0/N_458 ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_202_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_123_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_202_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_202_rs_net_1 ));
    INV_BA AFLSDF_INV_2 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_34_net_1 ), .Y(
        AFLSDF_INV_2_net_1));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_13_[2]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[2] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB3_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_13__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_234_i ), .ADn(VCC), .SLn(
        VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_13_rs[2] ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[6].REG_GEN.CONFIG_reg[6][7]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[7] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB12_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[6]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB2_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[6][7] ));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_104_set_RNIHBD51  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_104_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_232_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_13_rs[0] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_13_[0]_net_1 ));
    INV_BA AFLSDF_INV_8 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_45_net_1 ), .Y(
        AFLSDF_INV_8_net_1));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[9].REG_GEN.CONFIG_reg[9][3]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[3] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB15_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[9]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB5_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[9][3] ));
    CFG3 #( .INIT(8'hF2) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_247  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_14_[7]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_503 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_247_i ));
    CFG4 #( .INIT(16'hEC00) )  \CoreAPB3_0/u_mux_p_to_b3/PRDATA[25]  (
        .A(\CoreGPIO_0.xhdl1.GEN_BITS[0].APB_32.GPOUT_reg9 ), .B(
        \CoreGPIO_0.N_536 ), .C(
        \CoreGPIO_0.xhdl1.GEN_BITS[25].APB_32.GPOUT_reg[25] ), .D(
        CoreAPB3_0_APBmslave5_PSELx), .Y(
        \FIC_MSS_0_FIC_0_APB_MASTER_PRDATA[25] ));
    CFG4 #( .INIT(16'hF2F3) )  
        \CoreGPIO_0/xhdl1.GEN_BITS[17].APB_32.INTR_reg_230_0_o2_1_0[17]  
        (.A(\CoreGPIO_0/CONFIG_reg[17][6] ), .B(
        \CoreGPIO_0/edge_neg[17] ), .C(
        \CoreGPIO_0/INTR_reg_230_0_o2_0[17] ), .D(
        \CoreGPIO_0/CONFIG_reg[17][5] ), .Y(
        \CoreGPIO_0/INTR_reg_230_0_o2_1[17] ));
    CFG4 #( .INIT(16'hEFEE) )  
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_8[2]  (.A(
        \reg_apb_wrp_0/reg16x8_0/N_390 ), .B(
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_1[2]_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_5_[2]_net_1 ), .D(
        \reg_apb_wrp_0/reg16x8_0/N_490 ), .Y(
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_8[2]_net_1 ));
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_56  (
        .A(\reg_apb_wrp_0/reg16x8_0/mem_15_[2]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_497 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_56_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_5_[1]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[1] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB12_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_5__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_174_i ), .ADn(VCC), .SLn(
        VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_5_rs[1] ));
    CFG3 #( .INIT(8'hF2) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_241  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_14_[1]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_503 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_241_i ));
    CFG2 #( .INIT(4'h8) )  
        \CoreGPIO_0/xhdl1.GEN_BITS[4].REG_GPOUT.un44_GPIO_OUT_i  (.A(
        \CoreGPIO_0.xhdl1.GEN_BITS[4].APB_32.GPOUT_reg[4] ), .B(
        \CoreGPIO_0/CONFIG_reg[4][0] ), .Y(\GPIO_OUT_net_2[4] ));
    CFG2 #( .INIT(4'h7) )  \CoreGPIO_0/edge_both_2_sqmuxa_17_i  (.A(
        \CoreGPIO_0/N_248 ), .B(\CoreGPIO_0/CONFIG_reg[11][3] ), .Y(
        \CoreGPIO_0/N_186 ));
    CFG2 #( .INIT(4'h4) )  \CoreGPIO_0/PRDATA_0_iv_0_a2_0[21]  (.A(
        \CoreGPIO_0.N_247 ), .B(\CoreGPIO_0/INTR_reg[21] ), .Y(
        \CoreGPIO_0.N_544 ));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_8_[5]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[5] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB18_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_8__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_169_i ), .ADn(VCC), .SLn(
        VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_8_rs[5] ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[18].REG_GEN.CONFIG_reg[18][7]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[7] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB17_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[18]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB7_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[18][7] ));
    sdf_IOPAD_TRI \FIC_MSS_0/MDDR_ADDR_10_PAD/U_IOPAD  (.PAD(
        MDDR_ADDR[10]), .D(\FIC_MSS_0/DRAM_ADDR_net_0[10] ), .E(
        \FIC_MSS_0/MDDR_ADDR_10_PAD/EOUT ));
    INV_BA AFLSDF_INV_60 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_46_net_1 ), .Y(
        AFLSDF_INV_60_net_1));
    INV_BA AFLSDF_INV_0 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_9_net_1 ), .Y(
        AFLSDF_INV_0_net_1));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[21].REG_GEN.CONFIG_reg[21][1]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[1] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB13_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[21]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB3_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[21][1] ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_180  (.A(VCC), 
        .B(VCC), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/MGPIO22B_F2H_GPIN_net ), .IPB(), 
        .IPC());
    CFG3 #( .INIT(8'hF2) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_150  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_2_[6]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_501 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_150_i ));
    sdf_IOPAD_TRI \FIC_MSS_0/MDDR_RESET_N_PAD/U_IOPAD  (.PAD(
        MDDR_RESET_N), .D(\FIC_MSS_0/MSS_ADLIB_INST_DRAM_RSTN ), .E(
        \FIC_MSS_0/MDDR_RESET_N_PAD/EOUT ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_286  (.A(VCC), 
        .B(VCC), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PADDR_net[9] ), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[13] ), .IPC());
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_48_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB17_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_3__1_sqmuxa ), .ALn(
        AFLSDF_INV_92_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(GND)
        , .Q(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_48_set_net_1 ));
    CFG2 #( .INIT(4'h2) )  
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_a3_3[1]  (.A(
        \reg_apb_wrp_0/reg16x8_0/N_500 ), .B(
        \reg_apb_wrp_0/reg16x8_0/mem_13_[1]_net_1 ), .Y(
        \reg_apb_wrp_0/reg16x8_0/N_374 ));
    CFG4 #( .INIT(16'h0F35) )  
        \CoreGPIO_0/CONFIG_reg_o_2_31_bm_1_RNO_1[1]  (.A(
        \CoreGPIO_0.xhdl1.GEN_BITS[5].REG_GEN.CONFIG_reg[5][1] ), .B(
        \CoreGPIO_0/CONFIG_reg[21][1] ), .C(
        \CoreAPB3_0_APBmslave3_PADDR[6] ), .D(
        \CoreAPB3_0_APBmslave3_PADDR[5] ), .Y(
        \CoreGPIO_0/CONFIG_reg_o_2_21_1[1] ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[5].REG_GEN.CONFIG_reg[5][7]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[7] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB13_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[5]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB3_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[5][7] ));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_0_[4]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[4] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB19_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_0__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_132_i ), .ADn(VCC), .SLn(
        VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_0_rs[4] ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[2].REG_GEN.CONFIG_reg[2][4]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[4] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB17_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[2]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB7_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[2][4] ));
    CFG4 #( .INIT(16'hAC0F) )  
        \CoreGPIO_0/CONFIG_reg_o_2_31_bm_1_RNO_0[5]  (.A(
        \CoreGPIO_0/CONFIG_reg[9][5] ), .B(
        \CoreGPIO_0/CONFIG_reg[25][5] ), .C(
        \CoreGPIO_0/CONFIG_reg_o_2_18_1[5] ), .D(
        \CoreAPB3_0_APBmslave3_PADDR[5] ), .Y(
        \CoreGPIO_0/CONFIG_reg_o_2_31_bm_1_RNO_0[5]_net_1 ));
    CFG2 #( .INIT(4'h8) )  
        \reg_apb_wrp_0/reg16x8_0/mem_1__1_sqmuxa_0_a2_0_a3  (.A(
        \reg_apb_wrp_0/reg16x8_0/N_502 ), .B(
        \reg_apb_wrp_0/wr_enable_net_1 ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_1__1_sqmuxa ));
    CFG4 #( .INIT(16'h0002) )  
        \CoreGPIO_0/xhdl1.GEN_BITS[0].APB_32.GPOUT_reg9_0_a2_2_a2  (.A(
        \CoreAPB3_0_APBmslave3_PADDR[5] ), .B(
        \CoreAPB3_0_APBmslave3_PADDR[4] ), .C(\CoreGPIO_0/N_243 ), .D(
        \CoreGPIO_0.RDATA_32.un12_PRDATA_o_0_o2_1 ), .Y(
        \CoreGPIO_0.xhdl1.GEN_BITS[0].APB_32.GPOUT_reg9 ));
    CFG3 #( .INIT(8'hF2) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_155  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_3_[3]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_494 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_155_i ));
    CFG3 #( .INIT(8'hF2) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_179  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_9_[2]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_492 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_179_i ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_246_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_118_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_246_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_246_rs_net_1 ));
    CFG4 #( .INIT(16'h0F35) )  
        \CoreGPIO_0/CONFIG_reg_o_2_31_bm_RNO_2[0]  (.A(
        \CoreGPIO_0/CONFIG_reg[7][0] ), .B(
        \CoreGPIO_0/CONFIG_reg[23][0] ), .C(
        \CoreAPB3_0_APBmslave3_PADDR[6] ), .D(
        \CoreAPB3_0_APBmslave3_PADDR[5] ), .Y(
        \CoreGPIO_0/CONFIG_reg_o_2_28_1_1[0] ));
    CFG4 #( .INIT(16'h0F35) )  
        \CoreGPIO_0/CONFIG_reg_o_2_31_bm_RNO_1[4]  (.A(
        \CoreGPIO_0/CONFIG_reg[3][4] ), .B(
        \CoreGPIO_0/CONFIG_reg[19][4] ), .C(
        \CoreAPB3_0_APBmslave3_PADDR[6] ), .D(
        \CoreAPB3_0_APBmslave3_PADDR[5] ), .Y(
        \CoreGPIO_0/CONFIG_reg_o_2_25_1_1[4] ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_235_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_107_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_235_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_235_rs_net_1 ));
    CFG4 #( .INIT(16'h0F35) )  
        \CoreGPIO_0/CONFIG_reg_o_2_31_bm_1_RNO_2[5]  (.A(
        \CoreGPIO_0/CONFIG_reg[1][5] ), .B(
        \CoreGPIO_0/CONFIG_reg[17][5] ), .C(
        \CoreAPB3_0_APBmslave3_PADDR[6] ), .D(
        \CoreAPB3_0_APBmslave3_PADDR[5] ), .Y(
        \CoreGPIO_0/CONFIG_reg_o_2_18_1[5] ));
    CFG4 #( .INIT(16'hA9FF) )  
        \CoreGPIO_0/xhdl1.GEN_BITS[16].APB_32.INTR_reg_217_0_o2_0_0[16]  
        (.A(\CoreGPIO_0/CONFIG_reg[16][7] ), .B(
        \CoreGPIO_0/CONFIG_reg[16][6] ), .C(
        \CoreGPIO_0/CONFIG_reg[16][5] ), .D(
        \CoreGPIO_0/CONFIG_reg[16][3] ), .Y(
        \CoreGPIO_0/INTR_reg_217_0_o2_0[16] ));
    CFG4 #( .INIT(16'h0004) )  
        \reg_apb_wrp_0/reg16x8_0/WRITE_GEN.mem_4__2_i_a2[4]  (.A(
        \CoreAPB3_0_APBmslave3_PADDR[3] ), .B(
        \CoreAPB3_0_APBmslave3_PADDR[2] ), .C(
        \CoreAPB3_0_APBmslave3_PADDR[0] ), .D(
        \CoreAPB3_0_APBmslave3_PADDR[1] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/N_504 ));
    CFG4 #( .INIT(16'hAA08) )  
        \CoreGPIO_0/xhdl1.GEN_BITS[5].APB_32.edge_neg_79_iv_i_0[5]  (
        .A(\CoreGPIO_0/CONFIG_reg[5][3] ), .B(\CoreGPIO_0/edge_neg[5] )
        , .C(\CoreAPB3_0_APBmslave3_PWDATA[5] ), .D(\CoreGPIO_0/N_405 )
        , .Y(\CoreGPIO_0/N_115 ));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_43_set_RNIP8NP  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_43_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_139_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_1_rs[3] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_1_[3]_net_1 ));
    CFG4 #( .INIT(16'hBBFB) )  \CoreGPIO_0/edge_neg_2_sqmuxa_7_i_0  (
        .A(\CoreGPIO_0/N_405 ), .B(\CoreGPIO_0/CONFIG_reg[5][3] ), .C(
        \CoreGPIO_0/INTR_reg21 ), .D(\CoreGPIO_0.N_247 ), .Y(
        \CoreGPIO_0/N_60 ));
    CFG4 #( .INIT(16'h5410) )  \CoreGPIO_0/PRDATA_iv_0_0_0_1[1]  (.A(
        \CoreAPB3_0_APBmslave3_PADDR[7] ), .B(
        \CoreAPB3_0_APBmslave3_PADDR[2] ), .C(
        \CoreGPIO_0/CONFIG_reg_o_2_31_am[1]_net_1 ), .D(
        \CoreGPIO_0/CONFIG_reg_o_2_31_bm[1]_net_1 ), .Y(
        \CoreGPIO_0.PRDATA_iv_0_0_0_0[1] ));
    RGB \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB4  (.An(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_YNn_GSouth ), .ENn(GND), .YL()
        , .YR(\MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB4_rgbr_net_1 ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[4].APB_32.GPOUT_reg[4]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[4] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB13_rgbr_net_1 ), .EN(
        \CoreGPIO_0/GPOUT_reg_0_sqmuxa ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB3_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0.xhdl1.GEN_BITS[4].APB_32.GPOUT_reg[4] ));
    CFG4 #( .INIT(16'hAA08) )  
        \CoreGPIO_0/xhdl1.GEN_BITS[2].APB_32.edge_pos_37_iv_i_0[2]  (
        .A(\CoreGPIO_0/CONFIG_reg[2][3] ), .B(\CoreGPIO_0/edge_pos[2] )
        , .C(\CoreAPB3_0_APBmslave3_PWDATA[2] ), .D(\CoreGPIO_0/N_396 )
        , .Y(\CoreGPIO_0/N_105 ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_232_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_104_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_232_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_232_rs_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_193_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_98_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_193_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_193_rs_net_1 ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_30  (.A(GND), 
        .B(GND), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[6] ), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[13] ), .IPC());
    SLE \reg_apb_wrp_0/reg16x8_0/mem_6_[3]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[3] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB7_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_6__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_194_i ), .ADn(VCC), .SLn(
        VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_6_rs[3] ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_168_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_9_net_1 ), .EN(VCC), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_168_i ), .ADn(VCC), .SLn(
        VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_168_rs_net_1 ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_93  (.A(VCC), 
        .B(VCC), .C(VCC), .IPA(\FIC_MSS_0/MSS_ADLIB_INST/RX_DVF_net ), 
        .IPB(), .IPC());
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[11].REG_GEN.CONFIG_reg[11][4]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[4] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB10_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[11]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB0_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[11][4] ));
    IP_INTERFACE \FCCC_0/CCC_INST/IP_INTERFACE_8  (.A(VCC), .B(GND), 
        .C(VCC), .IPA(\FCCC_0/CCC_INST/PWRITE_net ), .IPB(
        \FCCC_0/CCC_INST/NGMUX2_SEL_net ), .IPC(
        \FCCC_0/CCC_INST/PWDATA_net[6] ));
    CFG3 #( .INIT(8'hF2) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_182  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_5_[5]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_490 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_182_i ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_27_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB8_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_5__1_sqmuxa ), .ALn(
        AFLSDF_INV_93_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(GND)
        , .Q(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_27_set_net_1 ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[30].APB_32.INTR_reg[30]  (.D(
        \CoreGPIO_0/INTR_reg_399[30] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB13_rgbr_net_1 ), .EN(VCC), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB3_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/INTR_reg[30] ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_11_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB13_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_4__1_sqmuxa ), .ALn(
        AFLSDF_INV_94_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(GND)
        , .Q(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_11_set_net_1 ));
    IOTRI_OB_EB \FIC_MSS_0/MDDR_ADDR_3_PAD/U_IOOUT  (.D(VCC), .E(VCC), 
        .DOUT(), .EOUT(\FIC_MSS_0/MDDR_ADDR_3_PAD/EOUT ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[18].REG_GEN.CONFIG_reg[18][0]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[0] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB16_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[18]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB6_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[18][0] ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[4].REG_GEN.CONFIG_reg[4][5]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[5] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB12_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[4]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB2_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[4][5] ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[16].REG_GEN.CONFIG_reg[16][4]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[4] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB15_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[16]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB5_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[16][4] ));
    CFG3 #( .INIT(8'hF2) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_170  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_4_[7]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_504 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_170_i ));
    CFG4 #( .INIT(16'hEAFA) )  \FIC_MSS_0/MSS_ADLIB_INST_RNO_5  (.A(
        \FIC_MSS_0/CoreAPB3_0_APBmslave5_PRDATA_m_0_0[6] ), .B(
        \CoreGPIO_0.PRDATA_iv_0_0_0_0[6] ), .C(
        CoreAPB3_0_APBmslave5_PSELx), .D(
        \FIC_MSS_0/CoreAPB3_0_APBmslave5_PRDATA_m_0_1_1[6] ), .Y(
        \FIC_MSS_0/FIC_MSS_0_FIC_0_APB_MASTER_PRDATA[6] ));
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_51  (
        .A(\reg_apb_wrp_0/reg16x8_0/mem_7_[3]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_498 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_51_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_226_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_18_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_226_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_226_rs_net_1 ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[31].REG_GEN.CONFIG_reg[31][7]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[7] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB10_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[31]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB0_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[31][7] ));
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_80  (
        .A(\reg_apb_wrp_0/reg16x8_0/mem_0_[0]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_496 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_80_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_8_[7]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[7] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB10_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_8__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_173_i ), .ADn(VCC), .SLn(
        VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_8_rs[7] ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_244_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_116_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_244_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_244_rs_net_1 ));
    CFG3 #( .INIT(8'hF2) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_175  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_9_[0]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_492 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_175_i ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[7].REG_GEN.CONFIG_reg[7][0]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[0] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB11_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[7]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB1_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[7][0] ));
    CFG2 #( .INIT(4'h8) )  
        \reg_apb_wrp_0/reg16x8_0/mem_9__1_sqmuxa_0_a3  (.A(
        \reg_apb_wrp_0/reg16x8_0/N_492 ), .B(
        \reg_apb_wrp_0/wr_enable_net_1 ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_9__1_sqmuxa ));
    CFG4 #( .INIT(16'hAA08) )  
        \CoreGPIO_0/xhdl1.GEN_BITS[6].APB_32.edge_pos_93_iv_i_0_0[6]  
        (.A(\CoreGPIO_0/CONFIG_reg[6][3] ), .B(
        \CoreGPIO_0/edge_pos[6] ), .C(
        \CoreAPB3_0_APBmslave3_PWDATA[6] ), .D(\CoreGPIO_0/N_689 ), .Y(
        \CoreGPIO_0/N_99 ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_106_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB3_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_13__1_sqmuxa ), .ALn(
        AFLSDF_INV_95_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(GND)
        , .Q(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_106_set_net_1 ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_52  (.A(GND), 
        .B(GND), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[6] ), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[13] ), .IPC());
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_90  (
        .A(\reg_apb_wrp_0/reg16x8_0/mem_11_[2]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_505 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_90_net_1 ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_198  (.A(VCC), 
        .B(VCC), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[2] ), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[14] ), .IPC());
    CFG4 #( .INIT(16'h7530) )  
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_1[7]  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_15_[7]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/mem_7_[7]_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/N_498 ), .D(
        \reg_apb_wrp_0/reg16x8_0/N_497 ), .Y(
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_1[7]_net_1 ));
    CFG4 #( .INIT(16'hBBFB) )  \CoreGPIO_0/edge_neg_2_sqmuxa_10_i_0  (
        .A(\CoreGPIO_0/N_395 ), .B(\CoreGPIO_0/CONFIG_reg[2][3] ), .C(
        \CoreGPIO_0/INTR_reg21 ), .D(\CoreGPIO_0.N_247 ), .Y(
        \CoreGPIO_0/N_56 ));
    CFG4 #( .INIT(16'hB383) )  \CoreGPIO_0/CONFIG_reg_o_2_31_bm[7]  (
        .A(\CoreGPIO_0/CONFIG_reg_o_2_31_bm_RNO[7]_net_1 ), .B(
        \CoreGPIO_0/CONFIG_reg_o_2_31_bm_1[7] ), .C(
        \CoreAPB3_0_APBmslave3_PADDR[3] ), .D(
        \CoreGPIO_0/CONFIG_reg_o_2_31_bm_RNO_0[7]_net_1 ), .Y(
        \CoreGPIO_0/CONFIG_reg_o_2_31_bm[7]_net_1 ));
    CFG3 #( .INIT(8'hF2) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_227  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_12_[3]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_495 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_227_i ));
    sdf_IOPAD_TRI \FIC_MSS_0/MDDR_ADDR_4_PAD/U_IOPAD  (.PAD(
        MDDR_ADDR[4]), .D(\FIC_MSS_0/DRAM_ADDR_net_0[4] ), .E(
        \FIC_MSS_0/MDDR_ADDR_4_PAD/EOUT ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[26].REG_GEN.CONFIG_reg[26][3]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[3] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB17_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[26]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB7_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[26][3] ));
    CFG3 #( .INIT(8'hF2) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_239  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_13_[7]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_500 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_239_i ));
    CFG3 #( .INIT(8'hF2) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_221  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_8_[1]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_499 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_221_i ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[3].REG_GEN.CONFIG_reg[3][2]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[2] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB10_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[3]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB0_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[3][2] ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_101  (.A(VCC), 
        .B(VCC), .C(VCC), .IPA(\FIC_MSS_0/MSS_ADLIB_INST/RCGF_net[1] ), 
        .IPB(\FIC_MSS_0/MSS_ADLIB_INST/RCGF_net[8] ), .IPC());
    CFG2 #( .INIT(4'h2) )  
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_a3_11[2]  (.A(
        \reg_apb_wrp_0/reg16x8_0/N_492 ), .B(
        \reg_apb_wrp_0/reg16x8_0/mem_9_[2]_net_1 ), .Y(
        \reg_apb_wrp_0/reg16x8_0/N_398 ));
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_43  (
        .A(\reg_apb_wrp_0/reg16x8_0/mem_1_[3]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_502 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_43_net_1 ));
    CFG4 #( .INIT(16'h4657) )  
        \CoreGPIO_0/CONFIG_reg_o_2_31_am_1_1[2]  (.A(
        \CoreAPB3_0_APBmslave3_PADDR[4] ), .B(
        \CoreAPB3_0_APBmslave3_PADDR[3] ), .C(
        \CoreGPIO_0/CONFIG_reg_o_2_31_am_1_1_RNO[2]_net_1 ), .D(
        \CoreGPIO_0/CONFIG_reg_o_2_31_am_1_RNO_0[2]_net_1 ), .Y(
        \CoreGPIO_0/CONFIG_reg_o_2_31_am_1[2] ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_224_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_17_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_224_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_224_rs_net_1 ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_42  (.A(GND), 
        .B(GND), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[25] ), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_WRITE_net ), .IPC());
    sdf_IOPAD_BI \FIC_MSS_0/MDDR_DM_RDQS_0_PAD/U_IOPAD  (.PAD(
        MDDR_DM_RDQS[0]), .D(\FIC_MSS_0/DRAM_DM_RDQS_OUT_net_0[0] ), 
        .E(\FIC_MSS_0/DM_OE_net_0[0] ), .Y(
        \FIC_MSS_0/MDDR_DM_RDQS_0_PAD_Y ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_284  (.A(VCC), 
        .B(VCC), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PADDR_net[7] ), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[11] ), .IPC());
    CFG4 #( .INIT(16'hAC0F) )  
        \CoreGPIO_0/CONFIG_reg_o_2_31_bm_1_1_RNO[6]  (.A(
        \CoreGPIO_0/CONFIG_reg[13][6] ), .B(
        \CoreGPIO_0/CONFIG_reg[29][6] ), .C(
        \CoreGPIO_0/CONFIG_reg_o_2_21_1[6] ), .D(
        \CoreAPB3_0_APBmslave3_PADDR[5] ), .Y(
        \CoreGPIO_0/CONFIG_reg_o_2_31_bm_1_1_RNO[6]_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_208_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_49_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_208_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_208_rs_net_1 ));
    INV_BA AFLSDF_INV_6 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_119_net_1 ), .Y(
        AFLSDF_INV_6_net_1));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_250  (.A(VCC), 
        .B(GND), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[62] ), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/F_ARID_HSEL1_net[2] ), .IPC());
    CFG4 #( .INIT(16'h2000) )  
        \CoreGPIO_0/xhdl1.GEN_BITS[10].REG_GEN.CONFIG_reg[10]2_0_a4_0_a2  
        (.A(\CoreAPB3_0_APBmslave3_PADDR[3] ), .B(
        \CoreAPB3_0_APBmslave3_PADDR[2] ), .C(\CoreGPIO_0/N_604 ), .D(
        \CoreGPIO_0/N_610 ), .Y(\CoreGPIO_0/CONFIG_reg[10]2 ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[9].REG_GEN.CONFIG_reg[9][6]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[6] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB15_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[9]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB5_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[9][6] ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_210_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_51_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_210_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_210_rs_net_1 ));
    CFG4 #( .INIT(16'hAC0F) )  
        \CoreGPIO_0/CONFIG_reg_o_2_31_am_1_1_RNO[3]  (.A(
        \CoreGPIO_0/CONFIG_reg[12][3] ), .B(
        \CoreGPIO_0/CONFIG_reg[28][3] ), .C(
        \CoreGPIO_0/CONFIG_reg_o_2_6_1[3] ), .D(
        \CoreAPB3_0_APBmslave3_PADDR[5] ), .Y(
        \CoreGPIO_0/CONFIG_reg_o_2_31_am_1_1_RNO[3]_net_1 ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[10].REG_GEN.CONFIG_reg[10][6]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[6] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB17_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[10]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB7_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[10][6] ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[17].REG_GEN.CONFIG_reg[17][3]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[3] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB15_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[17]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB5_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[17][3] ));
    CFG4 #( .INIT(16'h0F35) )  
        \CoreGPIO_0/CONFIG_reg_o_2_31_am_RNO_2[3]  (.A(
        \CoreGPIO_0/CONFIG_reg[6][3] ), .B(
        \CoreGPIO_0/CONFIG_reg[22][3] ), .C(
        \CoreAPB3_0_APBmslave3_PADDR[6] ), .D(
        \CoreAPB3_0_APBmslave3_PADDR[5] ), .Y(
        \CoreGPIO_0/CONFIG_reg_o_2_13_1_1[3] ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[28].REG_GEN.CONFIG_reg[28][5]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[5] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB12_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[28]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB2_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[28][5] ));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/mem_14__RNI53II[7]  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_119_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_247_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_14_rs[7] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_14_[7]_net_1 ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_257  (.A(VCC), 
        .B(VCC), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[5] ), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[17] ), .IPC());
    CFG3 #( .INIT(8'h04) )  
        \CoreGPIO_0/xhdl1.GEN_BITS[4].APB_32.INTR_reg_61_0_0_RNO_0[4]  
        (.A(\CoreGPIO_0/CONFIG_reg[4][5] ), .B(
        \CoreGPIO_0/edge_both[4] ), .C(\CoreGPIO_0/CONFIG_reg[4][6] ), 
        .Y(\CoreGPIO_0/INTR_reg_61_0_0_53_tz_1 ));
    CFG4 #( .INIT(16'hBBFB) )  \CoreGPIO_0/edge_pos_2_sqmuxa_i_0  (.A(
        \CoreGPIO_0/N_402 ), .B(\CoreGPIO_0/CONFIG_reg[0][3] ), .C(
        \CoreGPIO_0/INTR_reg21 ), .D(\CoreGPIO_0.N_247 ), .Y(
        \CoreGPIO_0/N_74 ));
    INV_BA AFLSDF_INV_79 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_67_net_1 ), .Y(
        AFLSDF_INV_79_net_1));
    SLE \reg_apb_wrp_0/reg16x8_0/data_out[1]  (.D(
        \reg_apb_wrp_0/reg16x8_0/temp_data[1]_net_1 ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB15_rgbr_net_1 ), .EN(VCC), .ALn(
        VCC), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreAPB3_0_APBmslave3_PRDATA[1] ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB18_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_4__1_sqmuxa ), .ALn(
        AFLSDF_INV_96_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(GND)
        , .Q(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_set_net_1 ));
    IOINFF_BYPASS \FIC_MSS_0/MDDR_DM_RDQS_1_PAD/U_IOINFF  (.A(
        \FIC_MSS_0/MDDR_DM_RDQS_1_PAD_Y ), .Y(
        \FIC_MSS_0/MDDR_DM_RDQS_1_PAD/YIN ));
    INV_BA AFLSDF_INV_77 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_15_net_1 ), .Y(
        AFLSDF_INV_77_net_1));
    IOTRI_OB_EB \FIC_MSS_0/MDDR_RESET_N_PAD/U_IOOUT  (.D(VCC), .E(VCC), 
        .DOUT(), .EOUT(\FIC_MSS_0/MDDR_RESET_N_PAD/EOUT ));
    CFG4 #( .INIT(16'hAA08) )  
        \CoreGPIO_0/xhdl1.GEN_BITS[0].APB_32.edge_neg_9_iv_i_0[0]  (.A(
        \CoreGPIO_0/CONFIG_reg[0][3] ), .B(\CoreGPIO_0/edge_neg[0] ), 
        .C(\CoreAPB3_0_APBmslave3_PWDATA[0] ), .D(\CoreGPIO_0/N_401 ), 
        .Y(\CoreGPIO_0/N_123 ));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_0_[2]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[2] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB11_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_0__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_129_i ), .ADn(VCC), .SLn(
        VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_0_rs[2] ));
    CFG4 #( .INIT(16'hAA08) )  
        \CoreGPIO_0/xhdl1.GEN_BITS[6].APB_32.edge_both_RNO[6]  (.A(
        \CoreGPIO_0/CONFIG_reg[6][3] ), .B(\CoreGPIO_0/edge_both[6] ), 
        .C(\CoreAPB3_0_APBmslave3_PWDATA[6] ), .D(\CoreGPIO_0/N_252_i )
        , .Y(\CoreGPIO_0/N_22_i_0 ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_194  (.A(GND), 
        .B(VCC), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/F_AWID_HSEL0_net[2] ), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[10] ), .IPC());
    CFG4 #( .INIT(16'h0002) )  
        \reg_apb_wrp_0/reg16x8_0/WRITE_GEN.mem_8__2_i_a2[7]  (.A(
        \CoreAPB3_0_APBmslave3_PADDR[3] ), .B(
        \CoreAPB3_0_APBmslave3_PADDR[2] ), .C(
        \CoreAPB3_0_APBmslave3_PADDR[0] ), .D(
        \CoreAPB3_0_APBmslave3_PADDR[1] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/N_499 ));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/mem_6__RNIRPQL[2]  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_33_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_192_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_6_rs[2] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_6_[2]_net_1 ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[24].REG_GEN.CONFIG_reg[24][4]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[4] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB15_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[24]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB5_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[24][4] ));
    CFG3 #( .INIT(8'hF2) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_213  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_7_[5]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_498 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_213_i ));
    CFG3 #( .INIT(8'h20) )  
        \CoreGPIO_0/xhdl1.GEN_BITS[24].APB_32.edge_both_RNO[24]  (.A(
        \CoreGPIO_0/CONFIG_reg[24][3] ), .B(
        \CoreAPB3_0_APBmslave3_PWDATA[24] ), .C(
        \CoreGPIO_0/edge_pos[24] ), .Y(\CoreGPIO_0/N_100_i_0 ));
    CFG2 #( .INIT(4'h2) )  
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_a3_11[4]  (.A(
        \reg_apb_wrp_0/reg16x8_0/N_492 ), .B(
        \reg_apb_wrp_0/reg16x8_0/mem_9_[4]_net_1 ), .Y(
        \reg_apb_wrp_0/reg16x8_0/N_432 ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[20].REG_GEN.CONFIG_reg[20][2]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[2] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB14_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[20]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB4_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[20][2] ));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_252_rs_RNIDU0M  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_60_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_252_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_15_rs[7] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_15_[7]_net_1 ));
    CFG4 #( .INIT(16'hF2F3) )  
        \CoreGPIO_0/xhdl1.GEN_BITS[24].APB_32.INTR_reg_321_0_o2_1_0[24]  
        (.A(\CoreGPIO_0/CONFIG_reg[24][6] ), .B(
        \CoreGPIO_0/edge_pos[24] ), .C(
        \CoreGPIO_0/INTR_reg_321_0_o2_0[24] ), .D(
        \CoreGPIO_0/CONFIG_reg[24][5] ), .Y(
        \CoreGPIO_0/INTR_reg_321_0_o2_1[24] ));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_17_set_RNI59QO  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_17_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_224_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_12_rs[1] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_12_[1]_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_238_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_110_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_238_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_238_rs_net_1 ));
    IP_INTERFACE \FCCC_0/CCC_INST/IP_INTERFACE_1  (.A(VCC), .B(VCC), 
        .C(VCC), .IPA(\FCCC_0/CCC_INST/CLK1_net ), .IPB(
        \FCCC_0/CCC_INST/PENABLE_net ), .IPC());
    CFG4 #( .INIT(16'h0F35) )  
        \CoreGPIO_0/CONFIG_reg_o_2_31_am_RNO_1[5]  (.A(
        \CoreGPIO_0/CONFIG_reg[2][5] ), .B(
        \CoreGPIO_0/CONFIG_reg[18][5] ), .C(
        \CoreAPB3_0_APBmslave3_PADDR[6] ), .D(
        \CoreAPB3_0_APBmslave3_PADDR[5] ), .Y(
        \CoreGPIO_0/CONFIG_reg_o_2_10_1_1[5] ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_56_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB6_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_15__1_sqmuxa ), .ALn(
        AFLSDF_INV_97_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(GND)
        , .Q(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_56_set_net_1 ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_2  (.A(
        \FIC_MSS_0/FIC_MSS_0_FIC_0_APB_MASTER_PRDATA[0] ), .B(VCC), .C(
        VCC), .IPA(\FIC_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[0] ), 
        .IPB(), .IPC());
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_59  (
        .A(\reg_apb_wrp_0/reg16x8_0/mem_15_[1]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_497 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_59_net_1 ));
    IOOUTFF_BYPASS \GPIO_OUT_obuf[3]/U0/U_IOOUTFF  (.A(
        \GPIO_OUT_obuf[3]/U0/DOUT1 ), .Y(\GPIO_OUT_obuf[3]/U0/DOUT ));
    CFG4 #( .INIT(16'h7530) )  
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_7[3]  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_10_[3]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/mem_2_[3]_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/N_501 ), .D(
        \reg_apb_wrp_0/reg16x8_0/N_491 ), .Y(
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_7[3]_net_1 ));
    CFG2 #( .INIT(4'h2) )  
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_a3_11[7]  (.A(
        \reg_apb_wrp_0/reg16x8_0/N_492 ), .B(
        \reg_apb_wrp_0/reg16x8_0/mem_9_[7]_net_1 ), .Y(
        \reg_apb_wrp_0/reg16x8_0/N_478 ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[8].REG_GEN.CONFIG_reg[8][7]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[7] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB11_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[8]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB1_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[8][7] ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_37_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB8_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_6__1_sqmuxa ), .ALn(
        AFLSDF_INV_98_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(GND)
        , .Q(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_37_set_net_1 ));
    CFG4 #( .INIT(16'hEFEE) )  
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_9[6]  (.A(
        \reg_apb_wrp_0/reg16x8_0/N_458 ), .B(
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_3[6]_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_1_[6]_net_1 ), .D(
        \reg_apb_wrp_0/reg16x8_0/N_502 ), .Y(
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_9[6]_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_92_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB19_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_11__1_sqmuxa ), .ALn(
        AFLSDF_INV_99_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(GND)
        , .Q(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_92_set_net_1 ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[1].APB_32.INTR_reg[1]  (.D(
        \CoreGPIO_0/INTR_reg_22[1] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB15_rgbr_net_1 ), .EN(VCC), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB5_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0.xhdl1.GEN_BITS[1].APB_32.INTR_reg[1] ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[10].REG_GEN.CONFIG_reg[10][5]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[5] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB17_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[10]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB7_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[10][5] ));
    CFG4 #( .INIT(16'hAC0F) )  
        \CoreGPIO_0/CONFIG_reg_o_2_31_bm_RNO_0[3]  (.A(
        \CoreGPIO_0/CONFIG_reg[15][3] ), .B(
        \CoreGPIO_0/CONFIG_reg[31][3] ), .C(
        \CoreGPIO_0/CONFIG_reg_o_2_28_1_1[3] ), .D(
        \CoreAPB3_0_APBmslave3_PADDR[5] ), .Y(
        \CoreGPIO_0/CONFIG_reg_o_2_31_bm_RNO_0[3]_net_1 ));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/mem_10__RNIHJPE[7]  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_100_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_205_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_10_rs[7] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_10_[7]_net_1 ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[18].REG_GEN.CONFIG_reg[18][1]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[1] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB16_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[18]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB6_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[18][1] ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[30].REG_GEN.CONFIG_reg[30][0]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[0] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB14_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[30]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB4_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[30][0] ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_235  (.A(VCC), 
        .B(VCC), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[33] ), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[45] ), .IPC());
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_129  (.A(GND), 
        .B(GND), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[4] ), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[11] ), .IPC());
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_125  (.A(GND), 
        .B(GND), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[0] ), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[7] ), .IPC());
    sdf_IOPAD_TRI \FIC_MSS_0/MDDR_ADDR_15_PAD/U_IOPAD  (.PAD(
        MDDR_ADDR[15]), .D(\FIC_MSS_0/DRAM_ADDR_net_0[15] ), .E(
        \FIC_MSS_0/MDDR_ADDR_15_PAD/EOUT ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[2].APB_32.edge_neg[2]  (.D(
        \CoreGPIO_0/N_119 ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB17_rgbr_net_1 ), .EN(
        \CoreGPIO_0/N_56 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB7_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/edge_neg[2] ));
    CFG2 #( .INIT(4'h4) )  \CoreGPIO_0/edge_neg_2_sqmuxa_8_i_a2  (.A(
        \CoreGPIO_0/gpin2[4] ), .B(
        \CoreGPIO_0.xhdl1.GEN_BITS[4].gpin3[4] ), .Y(
        \CoreGPIO_0/N_397 ));
    CFG2 #( .INIT(4'h7) )  \CoreGPIO_0/edge_both_2_sqmuxa_8_i  (.A(
        \CoreGPIO_0/N_248 ), .B(\CoreGPIO_0/CONFIG_reg[20][3] ), .Y(
        \CoreGPIO_0/N_196 ));
    CFG4 #( .INIT(16'h0001) )  
        \reg_apb_wrp_0/reg16x8_0/temp_data_RNO[4]  (.A(
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_0[4]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_1[4]_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_13[4]_net_1 ), .D(
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_9[4]_net_1 ), .Y(
        \reg_apb_wrp_0/reg16x8_0/N_19_i_0 ));
    CFG4 #( .INIT(16'h7350) )  
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_0_5[5]  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_14_[5]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/mem_6_[5]_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/N_503 ), .D(
        \reg_apb_wrp_0/reg16x8_0/N_493 ), .Y(
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_0_5[5]_net_1 ));
    CFG2 #( .INIT(4'h4) )  \CoreGPIO_0/edge_neg_2_sqmuxa_25_i_a2  (.A(
        \CoreGPIO_0/gpin2[0] ), .B(
        \CoreGPIO_0.xhdl1.GEN_BITS[0].gpin3[0] ), .Y(
        \CoreGPIO_0/N_401 ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_20_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB5_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_12__1_sqmuxa ), .ALn(
        AFLSDF_INV_100_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_20_set_net_1 ));
    IOTRI_OB_EB \FIC_MSS_0/MDDR_ADDR_9_PAD/U_IOOUT  (.D(VCC), .E(VCC), 
        .DOUT(), .EOUT(\FIC_MSS_0/MDDR_ADDR_9_PAD/EOUT ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[1].gpin3[1]  (.D(
        \CoreGPIO_0/gpin2[1] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB16_rgbr_net_1 ), .EN(VCC), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB6_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0.xhdl1.GEN_BITS[1].gpin3[1] ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_250_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_56_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_250_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_250_rs_net_1 ));
    CFG3 #( .INIT(8'h20) )  
        \CoreGPIO_0/xhdl1.GEN_BITS[11].APB_32.edge_both_RNO[11]  (.A(
        \CoreGPIO_0/CONFIG_reg[11][3] ), .B(
        \CoreAPB3_0_APBmslave3_PWDATA[11] ), .C(
        \CoreGPIO_0/edge_neg[11] ), .Y(\CoreGPIO_0/edge_neg_163[11] ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_103_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB13_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_10__1_sqmuxa ), .ALn(
        AFLSDF_INV_101_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_103_set_net_1 ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[6].APB_32.edge_pos[6]  (.D(
        \CoreGPIO_0/N_99 ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB12_rgbr_net_1 ), .EN(
        \CoreGPIO_0/N_72 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB2_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/edge_pos[6] ));
    CFG3 #( .INIT(8'h04) )  
        \CoreGPIO_0/xhdl1.GEN_BITS[5].APB_32.INTR_reg_74_0_0_RNO_0[5]  
        (.A(\CoreGPIO_0/CONFIG_reg[5][5] ), .B(
        \CoreGPIO_0/edge_both[5] ), .C(\CoreGPIO_0/CONFIG_reg[5][6] ), 
        .Y(\CoreGPIO_0/INTR_reg_74_0_0_54_tz_1 ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_132  (.A(GND), 
        .B(VCC), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[14] ), .IPB(), 
        .IPC());
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_12  (.A(
        \FIC_MSS_0_FIC_0_APB_MASTER_PRDATA[17] ), .B(VCC), .C(VCC), 
        .IPA(\FIC_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[17] ), .IPB(), 
        .IPC());
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_84  (.A(VCC), 
        .B(VCC), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[25] ), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/RXDF_net[0] ), .IPC());
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[0].APB_32.edge_pos[0]  (.D(
        \CoreGPIO_0/N_109 ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB9_rgbr_net_1 ), .EN(
        \CoreGPIO_0/N_74 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_YR ), .ADn(VCC), .SLn(
        VCC), .SD(GND), .LAT(GND), .Q(\CoreGPIO_0/edge_pos[0] ));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/mem_7__RNIA31M[7]  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_1_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_217_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_7_rs[7] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_7_[7]_net_1 ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_90  (.A(VCC), 
        .B(VCC), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[31] ), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/RXDF_net[6] ), .IPC());
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[2].gpin3[2]  (.D(
        \CoreGPIO_0/gpin2[2] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB17_rgbr_net_1 ), .EN(VCC), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB7_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0.xhdl1.GEN_BITS[2].gpin3[2] ));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_7_[5]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[5] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB9_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_7__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_213_i ), .ADn(VCC), .SLn(
        VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_7_rs[5] ));
    CFG4 #( .INIT(16'h330A) )  
        \CoreGPIO_0/xhdl1.GEN_BITS[8].APB_32.INTR_reg_113_0[8]  (.A(
        \CoreGPIO_0/INTR_reg[8] ), .B(
        \CoreGPIO_0/INTR_reg_113_0_o2_1[8] ), .C(
        \CoreAPB3_0_APBmslave3_PWDATA[8] ), .D(\CoreGPIO_0/N_248 ), .Y(
        \CoreGPIO_0/INTR_reg_113[8] ));
    CFG3 #( .INIT(8'hF2) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_189  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_9_[7]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_492 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_189_i ));
    CFG3 #( .INIT(8'hF2) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_244  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_14_[4]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_503 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_244_i ));
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_55  (
        .A(\reg_apb_wrp_0/reg16x8_0/mem_3_[7]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_494 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_55_net_1 ));
    IOINFF_BYPASS \GPIO_IN_ibuf[2]/U0/U_IOINFF  (.A(
        \GPIO_IN_ibuf[2]/U0/YIN1 ), .Y(\GPIO_IN_ibuf[2]/U0/YIN ));
    SLE \reg_apb_wrp_0/reg16x8_0/data_out[2]  (.D(
        \reg_apb_wrp_0/reg16x8_0/temp_data[2]_net_1 ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB15_rgbr_net_1 ), .EN(VCC), .ALn(
        VCC), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreAPB3_0_APBmslave3_PRDATA[2] ));
    CFG4 #( .INIT(16'hEFEE) )  
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_8[7]  (.A(
        \reg_apb_wrp_0/reg16x8_0/N_470 ), .B(
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_1[7]_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_5_[7]_net_1 ), .D(
        \reg_apb_wrp_0/reg16x8_0/N_490 ), .Y(
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_8[7]_net_1 ));
    CFG2 #( .INIT(4'h7) )  \CoreGPIO_0/edge_both_2_sqmuxa_29_i  (.A(
        \CoreGPIO_0/N_248 ), .B(\CoreGPIO_0/CONFIG_reg[26][3] ), .Y(
        \CoreGPIO_0/N_159 ));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_210_rs_RNIKVRC  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_51_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_210_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_7_rs[3] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_7_[3]_net_1 ));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/mem_7__RNI947S[6]  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_3_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_215_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_7_rs[6] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_7_[6]_net_1 ));
    CFG2 #( .INIT(4'hE) )  \reg_apb_wrp_0/PREADY_RNO  (.A(
        CoreAPB3_0_APBmslave3_PWRITE), .B(\reg_apb_wrp_0/fsm[1]_net_1 )
        , .Y(\reg_apb_wrp_0/N_64_i_0 ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_23_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB6_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_12__1_sqmuxa ), .ALn(
        AFLSDF_INV_102_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_23_set_net_1 ));
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_74  (
        .A(\reg_apb_wrp_0/reg16x8_0/mem_9_[2]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_492 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_74_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_19_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB1_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_12__1_sqmuxa ), .ALn(
        AFLSDF_INV_103_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_19_set_net_1 ));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_183_rs_RNI77551  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_76_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_183_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_9_rs[4] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_9_[4]_net_1 ));
    INV_BA AFLSDF_INV_12 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_87_net_1 ), .Y(
        AFLSDF_INV_12_net_1));
    CFG4 #( .INIT(16'hBBFB) )  \CoreGPIO_0/edge_pos_2_sqmuxa_3_i_0  (
        .A(\CoreGPIO_0/N_406 ), .B(\CoreGPIO_0/CONFIG_reg[5][3] ), .C(
        \CoreGPIO_0/INTR_reg21 ), .D(\CoreGPIO_0.N_247 ), .Y(
        \CoreGPIO_0/N_70 ));
    IOINFF_BYPASS \FIC_MSS_0/MDDR_DQ_9_PAD/U_IOINFF  (.A(
        \FIC_MSS_0/MDDR_DQ_9_PAD_Y ), .Y(\FIC_MSS_0/MDDR_DQ_9_PAD/YIN )
        );
    CFG3 #( .INIT(8'hF2) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_144  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_2_[0]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_501 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_144_i ));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_2_[0]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[0] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB0_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_2__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_144_i ), .ADn(VCC), .SLn(
        VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_2_rs[0] ));
    CFG4 #( .INIT(16'h4657) )  
        \CoreGPIO_0/CONFIG_reg_o_2_31_bm_1_1[2]  (.A(
        \CoreAPB3_0_APBmslave3_PADDR[4] ), .B(
        \CoreAPB3_0_APBmslave3_PADDR[3] ), .C(
        \CoreGPIO_0/CONFIG_reg_o_2_31_bm_1_1_RNO[2]_net_1 ), .D(
        \CoreGPIO_0/CONFIG_reg_o_2_31_bm_1_RNO_0[2]_net_1 ), .Y(
        \CoreGPIO_0/CONFIG_reg_o_2_31_bm_1[2] ));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_206_rs_RNIB7OM  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_127_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_206_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_7_rs[1] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_7_[1]_net_1 ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[1].REG_GEN.CONFIG_reg[1][7]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[7] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB14_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[1]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB4_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[1][7] ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_137_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_12_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_137_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_137_rs_net_1 ));
    CFG3 #( .INIT(8'h20) )  
        \CoreGPIO_0/xhdl1.GEN_BITS[17].APB_32.edge_both_RNO[17]  (.A(
        \CoreGPIO_0/CONFIG_reg[17][3] ), .B(
        \CoreAPB3_0_APBmslave3_PWDATA[17] ), .C(
        \CoreGPIO_0/edge_neg[17] ), .Y(\CoreGPIO_0/edge_neg_247[17] ));
    CFG3 #( .INIT(8'h76) )  \reg_apb_wrp_0/PREADY_RNO_0  (.A(
        \reg_apb_wrp_0/fsm[1]_net_1 ), .B(\reg_apb_wrp_0/fsm[0]_net_1 )
        , .C(CoreAPB3_0_APBmslave3_PSELx), .Y(\reg_apb_wrp_0/N_44_i_0 )
        );
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[31].REG_GEN.CONFIG_reg[31][4]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[4] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB12_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[31]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB2_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[31][4] ));
    CFG2 #( .INIT(4'h4) )  \CoreGPIO_0/PRDATA_0_iv_0_a2_0[19]  (.A(
        \CoreGPIO_0.N_247 ), .B(\CoreGPIO_0/INTR_reg[19] ), .Y(
        \CoreGPIO_0.N_548 ));
    IOIN_IB \GPIO_IN_ibuf[5]/U0/U_IOIN  (.YIN(\GPIO_IN_ibuf[5]/U0/YIN )
        , .E(GND), .Y(\GPIO_IN_c[5] ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_107_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB4_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_13__1_sqmuxa ), .ALn(
        AFLSDF_INV_104_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_107_set_net_1 ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_81  (.A(VCC), 
        .B(VCC), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[15] ), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[22] ), .IPC());
    CFG3 #( .INIT(8'hF2) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_180  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_5_[4]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_490 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_180_i ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_241_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_113_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_241_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_241_rs_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_66_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB8_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_8__1_sqmuxa ), .ALn(
        AFLSDF_INV_105_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_66_set_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_94_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB17_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_11__1_sqmuxa ), .ALn(
        AFLSDF_INV_106_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_94_set_net_1 ));
    sdf_IOPAD_TRI \FIC_MSS_0/MDDR_RAS_N_PAD/U_IOPAD  (.PAD(MDDR_RAS_N), 
        .D(\FIC_MSS_0/MSS_ADLIB_INST_DRAM_RASN ), .E(
        \FIC_MSS_0/MDDR_RAS_N_PAD/EOUT ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[10].APB_32.INTR_reg[10]  (.D(
        \CoreGPIO_0/INTR_reg_139[10] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB17_rgbr_net_1 ), .EN(VCC), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB7_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0.xhdl1.GEN_BITS[10].APB_32.INTR_reg[10] ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[14].REG_GEN.CONFIG_reg[14][1]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[1] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB15_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[14]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB5_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[14][1] ));
    INV_BA AFLSDF_INV_128 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_24_net_1 ), .Y(
        AFLSDF_INV_128_net_1));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[6].REG_GEN.CONFIG_reg[6][4]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[4] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB14_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[6]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB4_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[6][4] ));
    CFG3 #( .INIT(8'hF2) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_185  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_9_[5]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_492 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_185_i ));
    CFG2 #( .INIT(4'h2) )  \CoreGPIO_0/edge_pos_2_sqmuxa_6_i_a2  (.A(
        \CoreGPIO_0/gpin2[2] ), .B(
        \CoreGPIO_0.xhdl1.GEN_BITS[2].gpin3[2] ), .Y(
        \CoreGPIO_0/N_396 ));
    CFG2 #( .INIT(4'h8) )  
        \CoreGPIO_0/xhdl1.GEN_BITS[2].REG_GPOUT.un24_GPIO_OUT_i  (.A(
        \CoreGPIO_0/GPOUT_reg[2] ), .B(\CoreGPIO_0/CONFIG_reg[2][0] ), 
        .Y(\GPIO_OUT_net_2[2] ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[18].APB_32.edge_both[18]  (.D(
        \CoreGPIO_0/edge_neg_261[18] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB17_rgbr_net_1 ), .EN(
        \CoreGPIO_0/N_192 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB7_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/edge_neg[18] ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[12].REG_GEN.CONFIG_reg[12][0]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[0] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB12_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[12]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB2_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[12][0] ));
    CFG4 #( .INIT(16'hA9FF) )  
        \CoreGPIO_0/xhdl1.GEN_BITS[11].APB_32.INTR_reg_152_0_o2_0_0[11]  
        (.A(\CoreGPIO_0/CONFIG_reg[11][7] ), .B(
        \CoreGPIO_0/CONFIG_reg[11][6] ), .C(
        \CoreGPIO_0/CONFIG_reg[11][5] ), .D(
        \CoreGPIO_0/CONFIG_reg[11][3] ), .Y(
        \CoreGPIO_0/INTR_reg_152_0_o2_0[11] ));
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_57  (
        .A(\reg_apb_wrp_0/reg16x8_0/mem_15_[0]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_497 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_57_net_1 ));
    IOBI_IB_OB_EB \FIC_MSS_0/MDDR_DM_RDQS_1_PAD/U_IOBI  (.D(VCC), .E(
        VCC), .YIN(\FIC_MSS_0/MDDR_DM_RDQS_1_PAD/YIN ), .DOUT(), .EOUT(
        ), .Y());
    CFG2 #( .INIT(4'h4) )  \CoreGPIO_0/edge_neg_2_sqmuxa_i_0_0_a2  (.A(
        \CoreGPIO_0/gpin2[6] ), .B(
        \CoreGPIO_0.xhdl1.GEN_BITS[6].gpin3[6] ), .Y(
        \CoreGPIO_0/N_688 ));
    sdf_IOPAD_TRI \GPIO_OUT_obuf[5]/U0/U_IOPAD  (.PAD(GPIO_OUT[5]), .D(
        \GPIO_OUT_obuf[5]/U0/DOUT ), .E(\GPIO_OUT_obuf[5]/U0/EOUT ));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_7_[7]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[7] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB3_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_7__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_217_i ), .ADn(VCC), .SLn(
        VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_7_rs[7] ));
    CFG4 #( .INIT(16'h330A) )  
        \CoreGPIO_0/xhdl1.GEN_BITS[12].APB_32.INTR_reg_165_0[12]  (.A(
        \CoreGPIO_0/INTR_reg[12] ), .B(
        \CoreGPIO_0/INTR_reg_165_0_o2_1[12] ), .C(
        \CoreAPB3_0_APBmslave3_PWDATA[12] ), .D(\CoreGPIO_0/N_248 ), 
        .Y(\CoreGPIO_0/INTR_reg_165[12] ));
    CFG4 #( .INIT(16'hCC0A) )  
        \CoreGPIO_0/xhdl1.GEN_BITS[3].APB_32.INTR_reg_48_0[3]  (.A(
        \CoreGPIO_0.xhdl1.GEN_BITS[3].APB_32.INTR_reg[3] ), .B(
        \CoreGPIO_0/un34_intr ), .C(\CoreAPB3_0_APBmslave3_PWDATA[3] ), 
        .D(\CoreGPIO_0/N_248 ), .Y(\CoreGPIO_0/INTR_reg_48[3] ));
    IOINFF_BYPASS \GPIO_IN_ibuf[3]/U0/U_IOINFF  (.A(
        \GPIO_IN_ibuf[3]/U0/YIN1 ), .Y(\GPIO_IN_ibuf[3]/U0/YIN ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_221_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_5_net_1 ), .EN(VCC), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_221_i ), .ADn(VCC), .SLn(
        VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_221_rs_net_1 ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[5].REG_GEN.CONFIG_reg[5][4]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[4] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB14_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[5]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB4_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[5][4] ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[4].REG_GEN.CONFIG_reg[4][0]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[0] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB12_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[4]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB2_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[4][0] ));
    sdf_IOPAD_IN \GPIO_IN_ibuf[1]/U0/U_IOPAD  (.PAD(GPIO_IN[1]), .Y(
        \GPIO_IN_ibuf[1]/U0/YIN1 ));
    CFG2 #( .INIT(4'h2) )  
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_a3_11[0]  (.A(
        \reg_apb_wrp_0/reg16x8_0/N_492 ), .B(
        \reg_apb_wrp_0/reg16x8_0/mem_9_[0]_net_1 ), .Y(
        \reg_apb_wrp_0/reg16x8_0/N_366 ));
    CFG3 #( .INIT(8'h20) )  
        \CoreGPIO_0/xhdl1.GEN_BITS[19].APB_32.edge_both_RNO[19]  (.A(
        \CoreGPIO_0/CONFIG_reg[19][3] ), .B(
        \CoreAPB3_0_APBmslave3_PWDATA[19] ), .C(
        \CoreGPIO_0/edge_neg[19] ), .Y(\CoreGPIO_0/edge_neg_275[19] ));
    INV_BA AFLSDF_INV_35 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_65_net_1 ), .Y(
        AFLSDF_INV_35_net_1));
    CFG3 #( .INIT(8'h10) )  \CoreGPIO_0/RDATA_32.un12_PRDATA_o_0_a2  (
        .A(\CoreGPIO_0.RDATA_32.un12_PRDATA_o_0_o2_1 ), .B(
        \CoreGPIO_0/N_243 ), .C(\CoreGPIO_0/N_603 ), .Y(
        \CoreGPIO_0.RDATA_32.un12_PRDATA_o ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[30].REG_GEN.CONFIG_reg[30][3]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[3] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB12_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[30]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB2_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[30][3] ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_66  (.A(GND), 
        .B(VCC), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[27] ), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[0] ), .IPC());
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[28].REG_GEN.CONFIG_reg[28][3]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[3] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB14_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[28]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB4_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[28][3] ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_30_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB12_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_2__1_sqmuxa ), .ALn(
        AFLSDF_INV_107_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_30_set_net_1 ));
    IOIN_IB \FIC_MSS_0/MDDR_DQS_1_PAD/U_IOP  (.YIN(
        \FIC_MSS_0/MDDR_DQS_1_PAD/YIN ), .E(GND), .Y());
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_204_rs_RNI6O5C  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_125_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_204_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_7_rs[0] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_7_[0]_net_1 ));
    CFG3 #( .INIT(8'hF2) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_253  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_15_[4]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_497 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_253_i ));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/mem_2__RNIOC1E[1]  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_28_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_145_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_2_rs[1] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_2_[1]_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_197_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_96_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_197_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_197_rs_net_1 ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[2].REG_GEN.CONFIG_reg[2][5]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[5] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB17_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[2]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB7_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[2][5] ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[23].REG_GEN.CONFIG_reg[23][0]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[0] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB11_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[23]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB1_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[23][0] ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[7].REG_GEN.CONFIG_reg[7][3]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[3] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB10_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[7]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB0_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[7][3] ));
    CFG3 #( .INIT(8'hF2) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_224  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_12_[1]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_495 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_224_i ));
    CFG4 #( .INIT(16'h7530) )  
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_7[2]  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_10_[2]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/mem_2_[2]_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/N_501 ), .D(
        \reg_apb_wrp_0/reg16x8_0/N_491 ), .Y(
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_7[2]_net_1 ));
    CFG3 #( .INIT(8'hF2) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_218  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_11_[6]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_505 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_218_i ));
    CFG3 #( .INIT(8'hF2) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_132  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_0_[4]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_496 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_132_i ));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/mem_6__RNI3UQI[6]  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_121_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_200_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_6_rs[6] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_6_[6]_net_1 ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[5].gpin3[5]  (.D(
        \CoreGPIO_0/gpin2[5] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB10_rgbr_net_1 ), .EN(VCC), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB0_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0.xhdl1.GEN_BITS[5].gpin3[5] ));
    IOINFF_BYPASS \FIC_MSS_0/MDDR_DQ_14_PAD/U_IOINFF  (.A(
        \FIC_MSS_0/MDDR_DQ_14_PAD_Y ), .Y(
        \FIC_MSS_0/MDDR_DQ_14_PAD/YIN ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_213_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_54_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_213_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_213_rs_net_1 ));
    CFG4 #( .INIT(16'h0400) )  
        \CoreGPIO_0/xhdl1.GEN_BITS[12].REG_GEN.CONFIG_reg[12]2_0_a4_0_a2  
        (.A(\CoreAPB3_0_APBmslave3_PADDR[7] ), .B(\CoreGPIO_0/N_605 ), 
        .C(\CoreGPIO_0/N_243 ), .D(\CoreGPIO_0/INTR_reg21 ), .Y(
        \CoreGPIO_0/CONFIG_reg[12]2 ));
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_72  (
        .A(\reg_apb_wrp_0/reg16x8_0/mem_9_[0]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_492 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_72_net_1 ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[26].APB_32.GPOUT_reg[26]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[26] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB16_rgbr_net_1 ), .EN(
        \CoreGPIO_0/GPOUT_reg_0_sqmuxa ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB6_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/GPOUT_reg[26] ));
    CFG4 #( .INIT(16'hC5CA) )  
        \CoreGPIO_0/xhdl1.GEN_BITS[5].APB_32.INTR_reg_74_0_0_m2[5]  (
        .A(\CoreGPIO_0.xhdl1.GEN_BITS[5].gpin3[5] ), .B(
        \CoreGPIO_0/N_171 ), .C(\CoreGPIO_0/CONFIG_reg[5][6] ), .D(
        \CoreGPIO_0/CONFIG_reg[5][5] ), .Y(
        \CoreGPIO_0/INTR_reg_74_0_0_m2[5] ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_279  (.A(VCC), 
        .B(VCC), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PADDR_net[2] ), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[6] ), .IPC());
    CFG4 #( .INIT(16'hCC0A) )  
        \CoreGPIO_0/xhdl1.GEN_BITS[2].APB_32.INTR_reg_35_0_0[2]  (.A(
        \CoreGPIO_0/INTR_reg[2] ), .B(\CoreGPIO_0/N_1577_tz ), .C(
        \CoreAPB3_0_APBmslave3_PWDATA[2] ), .D(\CoreGPIO_0/N_248 ), .Y(
        \CoreGPIO_0/INTR_reg_35[2] ));
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_124  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_3_[1]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_494 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_124_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_3_[4]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[4] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB10_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_3__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_156_i ), .ADn(VCC), .SLn(
        VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_3_rs[4] ));
    CFG4 #( .INIT(16'hECA0) )  \FIC_MSS_0/MSS_ADLIB_INST_RNO_9  (.A(
        \CoreAPB3_0_APBmslave3_PRDATA[2] ), .B(
        CoreAPB3_0_APBmslave5_PSELx), .C(CoreAPB3_0_APBmslave3_PSELx), 
        .D(\CoreGPIO_0.PRDATA_iv_0_0_1[2] ), .Y(
        \FIC_MSS_0/CoreAPB3_0_APBmslave5_PRDATA_m_0_0[2] ));
    IOIN_IB \FIC_MSS_0/MDDR_DQS_0_PAD/U_IOP  (.YIN(
        \FIC_MSS_0/MDDR_DQS_0_PAD/YIN ), .E(GND), .Y());
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[27].REG_GEN.CONFIG_reg[27][6]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[6] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB9_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[27]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_YR ), .ADn(VCC), .SLn(
        VCC), .SD(GND), .LAT(GND), .Q(\CoreGPIO_0/CONFIG_reg[27][6] ));
    CFG2 #( .INIT(4'h4) )  \CoreGPIO_0/edge_neg_2_sqmuxa_9_i_a2  (.A(
        \CoreGPIO_0/gpin2[3] ), .B(
        \CoreGPIO_0.xhdl1.GEN_BITS[3].gpin3[3] ), .Y(
        \CoreGPIO_0/N_686 ));
    INV_BA AFLSDF_INV_74 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_74_net_1 ), .Y(
        AFLSDF_INV_74_net_1));
    CFG4 #( .INIT(16'hB383) )  \CoreGPIO_0/CONFIG_reg_o_2_31_bm[5]  (
        .A(\CoreGPIO_0/CONFIG_reg_o_2_31_bm_RNO[5]_net_1 ), .B(
        \CoreGPIO_0/CONFIG_reg_o_2_31_bm_1[5] ), .C(
        \CoreAPB3_0_APBmslave3_PADDR[3] ), .D(
        \CoreGPIO_0/CONFIG_reg_o_2_31_bm_RNO_0[5]_net_1 ), .Y(
        \CoreGPIO_0/CONFIG_reg_o_2_31_bm[5]_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_33_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB12_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_6__1_sqmuxa ), .ALn(
        AFLSDF_INV_108_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_33_set_net_1 ));
    IOINFF_BYPASS \FIC_MSS_0/MDDR_DQ_1_PAD/U_IOINFF  (.A(
        \FIC_MSS_0/MDDR_DQ_1_PAD_Y ), .Y(\FIC_MSS_0/MDDR_DQ_1_PAD/YIN )
        );
    sdf_IOPAD_TRI \FIC_MSS_0/MDDR_ADDR_3_PAD/U_IOPAD  (.PAD(
        MDDR_ADDR[3]), .D(\FIC_MSS_0/DRAM_ADDR_net_0[3] ), .E(
        \FIC_MSS_0/MDDR_ADDR_3_PAD/EOUT ));
    CFG4 #( .INIT(16'hA820) )  
        \CoreGPIO_0/xhdl1.GEN_BITS[3].REG_INT.un34_intr_u_ns  (.A(
        \CoreGPIO_0/CONFIG_reg[3][3] ), .B(
        \CoreGPIO_0/CONFIG_reg[3][7] ), .C(\CoreGPIO_0/un34_intr_u_bm )
        , .D(\CoreGPIO_0/un34_intr_u_ns_1 ), .Y(\CoreGPIO_0/un34_intr )
        );
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_205  (.A(VCC), 
        .B(GND), .C(GND), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/F_AWADDR_HADDR0_net[23] ), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/F_AWLEN_HBURST0_net[1] ), .IPC(
        \FIC_MSS_0/MSS_ADLIB_INST/F_WLAST_net ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_52_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB10_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_3__1_sqmuxa ), .ALn(
        AFLSDF_INV_109_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_52_set_net_1 ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[22].APB_32.edge_both[22]  (.D(
        \CoreGPIO_0/edge_neg_317[22] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB13_rgbr_net_1 ), .EN(
        \CoreGPIO_0/N_200 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB3_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/edge_neg[22] ));
    CFG4 #( .INIT(16'h0F35) )  
        \CoreGPIO_0/CONFIG_reg_o_2_31_am_1_RNO_1[5]  (.A(
        \CoreGPIO_0/CONFIG_reg[4][5] ), .B(
        \CoreGPIO_0/CONFIG_reg[20][5] ), .C(
        \CoreAPB3_0_APBmslave3_PADDR[6] ), .D(
        \CoreAPB3_0_APBmslave3_PADDR[5] ), .Y(
        \CoreGPIO_0/CONFIG_reg_o_2_6_1[5] ));
    IOTRI_OB_EB \FIC_MSS_0/MDDR_ADDR_10_PAD/U_IOOUT  (.D(VCC), .E(VCC), 
        .DOUT(), .EOUT(\FIC_MSS_0/MDDR_ADDR_10_PAD/EOUT ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_166_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_67_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_166_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_166_rs_net_1 ));
    CFG4 #( .INIT(16'hF2F3) )  
        \CoreGPIO_0/xhdl1.GEN_BITS[30].APB_32.INTR_reg_399_0_o2_1_0[30]  
        (.A(\CoreGPIO_0/CONFIG_reg[30][6] ), .B(
        \CoreGPIO_0/edge_pos[30] ), .C(
        \CoreGPIO_0/INTR_reg_399_0_o2_0[30] ), .D(
        \CoreGPIO_0/CONFIG_reg[30][5] ), .Y(
        \CoreGPIO_0/INTR_reg_399_0_o2_1[30] ));
    IOTRI_OB_EB \FIC_MSS_0/MDDR_WE_N_PAD/U_IOOUT  (.D(VCC), .E(VCC), 
        .DOUT(), .EOUT(\FIC_MSS_0/MDDR_WE_N_PAD/EOUT ));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_1_[5]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[5] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB15_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_1__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_141_i ), .ADn(VCC), .SLn(
        VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_1_rs[5] ));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_11_[0]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[0] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB16_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_11__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_207_i ), .ADn(VCC), .SLn(
        VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_11_rs[0] ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[14].REG_GEN.CONFIG_reg[14][0]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[0] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB14_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[14]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB4_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[14][0] ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[1].gpin1[1]  (.D(\GPIO_IN_c[1] ), 
        .CLK(\FCCC_0/GL1_INST/U0_RGB1_RGB16_rgbr_net_1 ), .EN(VCC), 
        .ALn(\MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB6_rgbr_net_1 ), 
        .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/gpin1[1] ));
    CFG4 #( .INIT(16'h0100) )  
        \reg_apb_wrp_0/reg16x8_0/WRITE_GEN.mem_2__2_i_a2[6]  (.A(
        \CoreAPB3_0_APBmslave3_PADDR[3] ), .B(
        \CoreAPB3_0_APBmslave3_PADDR[2] ), .C(
        \CoreAPB3_0_APBmslave3_PADDR[0] ), .D(
        \CoreAPB3_0_APBmslave3_PADDR[1] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/N_501 ));
    CFG4 #( .INIT(16'hEFEE) )  
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_9[1]  (.A(
        \reg_apb_wrp_0/reg16x8_0/N_382 ), .B(
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_3[1]_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_1_[1]_net_1 ), .D(
        \reg_apb_wrp_0/reg16x8_0/N_502 ), .Y(
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_9[1]_net_1 ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[12].REG_GEN.CONFIG_reg[12][1]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[1] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB12_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[12]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB2_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[12][1] ));
    CFG3 #( .INIT(8'h20) )  
        \CoreGPIO_0/xhdl1.GEN_BITS[12].APB_32.edge_both_RNO[12]  (.A(
        \CoreGPIO_0/CONFIG_reg[12][3] ), .B(
        \CoreAPB3_0_APBmslave3_PWDATA[12] ), .C(
        \CoreGPIO_0/edge_neg[12] ), .Y(\CoreGPIO_0/edge_neg_177[12] ));
    CFG4 #( .INIT(16'h0F35) )  
        \CoreGPIO_0/CONFIG_reg_o_2_31_am_RNO_2[5]  (.A(
        \CoreGPIO_0/CONFIG_reg[6][5] ), .B(
        \CoreGPIO_0/CONFIG_reg[22][5] ), .C(
        \CoreAPB3_0_APBmslave3_PADDR[6] ), .D(
        \CoreAPB3_0_APBmslave3_PADDR[5] ), .Y(
        \CoreGPIO_0/CONFIG_reg_o_2_13_1_1[5] ));
    CFG4 #( .INIT(16'h330A) )  
        \CoreGPIO_0/xhdl1.GEN_BITS[17].APB_32.INTR_reg_230_0[17]  (.A(
        \CoreGPIO_0/INTR_reg[17] ), .B(
        \CoreGPIO_0/INTR_reg_230_0_o2_1[17] ), .C(
        \CoreAPB3_0_APBmslave3_PWDATA[17] ), .D(\CoreGPIO_0/N_248 ), 
        .Y(\CoreGPIO_0/INTR_reg_230[17] ));
    CFG4 #( .INIT(16'hAC0F) )  
        \CoreGPIO_0/CONFIG_reg_o_2_31_am_RNO[1]  (.A(
        \CoreGPIO_0/CONFIG_reg[10][1] ), .B(
        \CoreGPIO_0/CONFIG_reg[26][1] ), .C(
        \CoreGPIO_0/CONFIG_reg_o_2_10_1_1[1] ), .D(
        \CoreAPB3_0_APBmslave3_PADDR[5] ), .Y(
        \CoreGPIO_0/CONFIG_reg_o_2_31_am_RNO[1]_net_1 ));
    CFG4 #( .INIT(16'h7530) )  
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_7[0]  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_10_[0]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/mem_2_[0]_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/N_501 ), .D(
        \reg_apb_wrp_0/reg16x8_0/N_491 ), .Y(
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_7[0]_net_1 ));
    INV_BA AFLSDF_INV_99 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_92_net_1 ), .Y(
        AFLSDF_INV_99_net_1));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_102  (.A(VCC), 
        .B(VCC), .C(VCC), .IPA(\FIC_MSS_0/MSS_ADLIB_INST/RCGF_net[2] ), 
        .IPB(\FIC_MSS_0/MSS_ADLIB_INST/RCGF_net[9] ), .IPC());
    RGB \FCCC_0/GL1_INST/U0_RGB1_RGB19  (.An(
        \FCCC_0/GL1_INST/U0_YNn_GSouth ), .ENn(GND), .YL(
        \FCCC_0/GL1_INST/U0_RGB1_RGB19_rgbl_net_1 ), .YR());
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_150_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_38_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_150_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_150_rs_net_1 ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_34  (.A(VCC), 
        .B(GND), .C(VCC), .IPA(), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[17] ), .IPC());
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[3].REG_GEN.CONFIG_reg[3][7]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[7] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB9_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[3]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_YR ), .ADn(VCC), .SLn(
        VCC), .SD(GND), .LAT(GND), .Q(\CoreGPIO_0/CONFIG_reg[3][7] ));
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_64  (
        .A(\reg_apb_wrp_0/reg16x8_0/mem_8_[2]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_499 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_64_net_1 ));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_250_rs_RNIB6LI  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_56_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_250_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_15_rs[2] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_15_[2]_net_1 ));
    INV_BA AFLSDF_INV_42 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_82_net_1 ), .Y(
        AFLSDF_INV_42_net_1));
    INV_BA AFLSDF_INV_115 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_6_net_1 ), .Y(
        AFLSDF_INV_115_net_1));
    INV_BA AFLSDF_INV_97 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_56_net_1 ), .Y(
        AFLSDF_INV_97_net_1));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_138_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_14_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_138_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_138_rs_net_1 ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[10].REG_GEN.CONFIG_reg[10][3]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[3] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB17_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[10]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB7_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[10][3] ));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_6_[1]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[1] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB6_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_6__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_190_i ), .ADn(VCC), .SLn(
        VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_6_rs[1] ));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_20_set_RNI616Q  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_20_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_228_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_12_rs[4] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_12_[4]_net_1 ));
    CFG4 #( .INIT(16'hAC0F) )  
        \CoreGPIO_0/CONFIG_reg_o_2_31_bm_1_1_RNO[1]  (.A(
        \CoreGPIO_0/CONFIG_reg[13][1] ), .B(
        \CoreGPIO_0/CONFIG_reg[29][1] ), .C(
        \CoreGPIO_0/CONFIG_reg_o_2_21_1[1] ), .D(
        \CoreAPB3_0_APBmslave3_PADDR[5] ), .Y(
        \CoreGPIO_0/CONFIG_reg_o_2_31_bm_1_1_RNO[1]_net_1 ));
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_24  (
        .A(\reg_apb_wrp_0/reg16x8_0/mem_1_[7]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_502 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_24_net_1 ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[20].REG_GEN.CONFIG_reg[20][5]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[5] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB12_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[20]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB2_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[20][5] ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[28].REG_GEN.CONFIG_reg[28][6]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[6] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB12_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[28]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB2_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[28][6] ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[13].REG_GEN.CONFIG_reg[13][1]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[1] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB13_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[13]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB3_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[13][1] ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_178  (.A(VCC), 
        .B(VCC), .C(VCC), .IPA(), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/MMUART0_DSR_F2H_SCP_net ), .IPC());
    CFG3 #( .INIT(8'h40) )  \CoreGPIO_0/PRDATA_0_iv_0_a2[18]  (.A(
        \CoreGPIO_0.N_246 ), .B(\CoreGPIO_0/GPOUT_reg[18] ), .C(
        \CoreAPB3_0_APBmslave3_PADDR[5] ), .Y(\CoreGPIO_0.N_549 ));
    CFG3 #( .INIT(8'h54) )  \reg_apb_wrp_0/fsm_RNIENS51[1]  (.A(
        \reg_apb_wrp_0/fsm[1]_net_1 ), .B(\reg_apb_wrp_0/fsm[0]_net_1 )
        , .C(CoreAPB3_0_APBmslave3_PSELx), .Y(\reg_apb_wrp_0/N_45_i_0 )
        );
    sdf_IOPAD_TRI \FIC_MSS_0/MDDR_BA_0_PAD/U_IOPAD  (.PAD(MDDR_BA[0]), 
        .D(\FIC_MSS_0/DRAM_BA_net_0[0] ), .E(
        \FIC_MSS_0/MDDR_BA_0_PAD/EOUT ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[1].gpin2[1]  (.D(
        \CoreGPIO_0/gpin1[1] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB16_rgbr_net_1 ), .EN(VCC), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB6_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(\CoreGPIO_0/gpin2[1] )
        );
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[11].APB_32.edge_both[11]  (.D(
        \CoreGPIO_0/edge_neg_163[11] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB9_rgbr_net_1 ), .EN(
        \CoreGPIO_0/N_186 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_YR ), .ADn(VCC), .SLn(
        VCC), .SD(GND), .LAT(GND), .Q(\CoreGPIO_0/edge_neg[11] ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_253_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_58_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_253_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_253_rs_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_216_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_93_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_216_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_216_rs_net_1 ));
    INV_BA AFLSDF_INV_31 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_86_net_1 ), .Y(
        AFLSDF_INV_31_net_1));
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_106  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_13_[2]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_500 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_106_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_1_[7]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[7] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB16_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_1__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_143_i ), .ADn(VCC), .SLn(
        VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_1_rs[7] ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_31  (.A(GND), 
        .B(GND), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[7] ), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[14] ), .IPC());
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[2].APB_32.edge_pos[2]  (.D(
        \CoreGPIO_0/N_105 ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB17_rgbr_net_1 ), .EN(
        \CoreGPIO_0/N_64 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB7_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/edge_pos[2] ));
    CFG2 #( .INIT(4'h7) )  \CoreGPIO_0/edge_both_2_sqmuxa_4_i  (.A(
        \CoreGPIO_0/N_248 ), .B(\CoreGPIO_0/CONFIG_reg[15][3] ), .Y(
        \CoreGPIO_0/edge_pos_2_sqmuxa_7_i_1 ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[21].APB_32.edge_both[21]  (.D(
        \CoreGPIO_0/edge_neg_303[21] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB13_rgbr_net_1 ), .EN(
        \CoreGPIO_0/N_198 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB3_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/edge_neg[21] ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[7].REG_GEN.CONFIG_reg[7][6]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[6] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB10_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[7]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB0_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[7][6] ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_56  (.A(GND), 
        .B(GND), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[10] ), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[17] ), .IPC());
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/mem_10__RNIDDPI[5]  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_102_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_201_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_10_rs[5] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_10_[5]_net_1 ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[11].REG_GEN.CONFIG_reg[11][2]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[2] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB10_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[11]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB0_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[11][2] ));
    CFG4 #( .INIT(16'h5410) )  \CoreGPIO_0/PRDATA_iv_0_0_0_1[2]  (.A(
        \CoreAPB3_0_APBmslave3_PADDR[7] ), .B(
        \CoreAPB3_0_APBmslave3_PADDR[2] ), .C(
        \CoreGPIO_0/CONFIG_reg_o_2_31_am[2]_net_1 ), .D(
        \CoreGPIO_0/CONFIG_reg_o_2_31_bm[2]_net_1 ), .Y(
        \CoreGPIO_0.PRDATA_iv_0_0_0_0[2] ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_164_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_6_net_1 ), .EN(VCC), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_164_i ), .ADn(VCC), .SLn(
        VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_164_rs_net_1 ));
    CFG4 #( .INIT(16'hCC0A) )  
        \CoreGPIO_0/xhdl1.GEN_BITS[1].APB_32.INTR_reg_22_0_0[1]  (.A(
        \CoreGPIO_0.xhdl1.GEN_BITS[1].APB_32.INTR_reg[1] ), .B(
        \CoreGPIO_0/N_1576_tz ), .C(\CoreAPB3_0_APBmslave3_PWDATA[1] ), 
        .D(\CoreGPIO_0/N_248 ), .Y(\CoreGPIO_0/INTR_reg_22[1] ));
    sdf_IOPAD_TRI \FIC_MSS_0/MDDR_ADDR_8_PAD/U_IOPAD  (.PAD(
        MDDR_ADDR[8]), .D(\FIC_MSS_0/DRAM_ADDR_net_0[8] ), .E(
        \FIC_MSS_0/MDDR_ADDR_8_PAD/EOUT ));
    CFG4 #( .INIT(16'hA9FF) )  
        \CoreGPIO_0/xhdl1.GEN_BITS[14].APB_32.INTR_reg_191_0_o2_0_0[14]  
        (.A(\CoreGPIO_0/CONFIG_reg[14][7] ), .B(
        \CoreGPIO_0/CONFIG_reg[14][6] ), .C(
        \CoreGPIO_0/CONFIG_reg[14][5] ), .D(
        \CoreGPIO_0/CONFIG_reg[14][3] ), .Y(
        \CoreGPIO_0/INTR_reg_191_0_o2_0[14] ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_179_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_74_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_179_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_179_rs_net_1 ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[8].REG_GEN.CONFIG_reg[8][4]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[4] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB15_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[8]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB5_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[8][4] ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_141  (.A(VCC), 
        .B(VCC), .C(VCC), .IPA(\FIC_MSS_0/MSS_ADLIB_INST/F2HCALIB_net )
        , .IPB(\FIC_MSS_0/MSS_ADLIB_INST/SPI0_CLK_IN_net ), .IPC());
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[10].APB_32.edge_both[10]  (.D(
        \CoreGPIO_0/edge_neg_149[10] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB17_rgbr_net_1 ), .EN(
        \CoreGPIO_0/N_184 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB7_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/edge_pos[10] ));
    CFG2 #( .INIT(4'h4) )  \CoreGPIO_0/PRDATA_0_iv_0_a2_0[11]  (.A(
        \CoreGPIO_0.N_247 ), .B(\CoreGPIO_0/INTR_reg[11] ), .Y(
        \CoreGPIO_0.N_564 ));
    CFG4 #( .INIT(16'hAC0F) )  
        \CoreGPIO_0/CONFIG_reg_o_2_31_am_1_RNO_0[0]  (.A(
        \CoreGPIO_0/CONFIG_reg[8][0] ), .B(
        \CoreGPIO_0/CONFIG_reg[24][0] ), .C(
        \CoreGPIO_0/CONFIG_reg_o_2_3_1[0] ), .D(
        \CoreAPB3_0_APBmslave3_PADDR[5] ), .Y(
        \CoreGPIO_0/CONFIG_reg_o_2_31_am_1_RNO_0[0]_net_1 ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_85  (.A(VCC), 
        .B(VCC), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[26] ), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/RXDF_net[1] ), .IPC());
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[28].REG_GEN.CONFIG_reg[28][4]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[4] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB14_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[28]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB4_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[28][4] ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[25].REG_GEN.CONFIG_reg[25][3]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[3] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB15_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[25]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB5_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[25][3] ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_46  (.A(VCC), 
        .B(GND), .C(VCC), .IPA(), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[0] ), .IPC());
    SLE \reg_apb_wrp_0/reg16x8_0/mem_13_[3]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[3] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB4_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_13__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_235_i ), .ADn(VCC), .SLn(
        VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_13_rs[3] ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_54_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB8_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_7__1_sqmuxa ), .ALn(
        AFLSDF_INV_110_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_54_set_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_3_[2]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[2] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB17_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_3__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_154_i ), .ADn(VCC), .SLn(
        VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_3_rs[2] ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_174  (.A(VCC), 
        .B(VCC), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/MGPIO25B_F2H_GPIN_net ), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/MMUART0_DTR_F2H_SCP_net ), .IPC());
    CFG4 #( .INIT(16'hAC0F) )  
        \CoreGPIO_0/CONFIG_reg_o_2_31_am_RNO_0[2]  (.A(
        \CoreGPIO_0/CONFIG_reg[14][2] ), .B(
        \CoreGPIO_0/CONFIG_reg[30][2] ), .C(
        \CoreGPIO_0/CONFIG_reg_o_2_13_1_1[2] ), .D(
        \CoreAPB3_0_APBmslave3_PADDR[5] ), .Y(
        \CoreGPIO_0/CONFIG_reg_o_2_31_am_RNO_0[2]_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_198_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_39_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_198_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_198_rs_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_214_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_92_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_214_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_214_rs_net_1 ));
    IOTRI_OB_EB \FIC_MSS_0/MDDR_ADDR_8_PAD/U_IOOUT  (.D(VCC), .E(VCC), 
        .DOUT(), .EOUT(\FIC_MSS_0/MDDR_ADDR_8_PAD/EOUT ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_62_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB7_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_15__1_sqmuxa ), .ALn(
        AFLSDF_INV_111_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_62_set_net_1 ));
    CFG4 #( .INIT(16'hAA08) )  
        \CoreGPIO_0/xhdl1.GEN_BITS[3].APB_32.edge_both_51_iv_i[3]  (.A(
        \CoreGPIO_0/CONFIG_reg[3][3] ), .B(\CoreGPIO_0/edge_both[3] ), 
        .C(\CoreAPB3_0_APBmslave3_PWDATA[3] ), .D(\CoreGPIO_0/N_253_i )
        , .Y(\CoreGPIO_0/edge_both_51_iv_i_0[3] ));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_4_[6]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[6] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB17_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_4__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_168_i ), .ADn(VCC), .SLn(
        VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_4_rs[6] ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[31].APB_32.GPOUT_reg[31]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[31] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB9_rgbr_net_1 ), .EN(
        \CoreGPIO_0/GPOUT_reg_0_sqmuxa ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_YR ), .ADn(VCC), .SLn(
        VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0.xhdl1.GEN_BITS[31].APB_32.GPOUT_reg[31] ));
    CFG4 #( .INIT(16'hEC00) )  \CoreAPB3_0/u_mux_p_to_b3/PRDATA[29]  (
        .A(\CoreGPIO_0.xhdl1.GEN_BITS[0].APB_32.GPOUT_reg9 ), .B(
        \CoreGPIO_0.N_528 ), .C(
        \CoreGPIO_0.xhdl1.GEN_BITS[29].APB_32.GPOUT_reg[29] ), .D(
        CoreAPB3_0_APBmslave5_PSELx), .Y(
        \FIC_MSS_0_FIC_0_APB_MASTER_PRDATA[29] ));
    SLE \reg_apb_wrp_0/reg16x8_0/temp_data[3]  (.D(
        \reg_apb_wrp_0/reg16x8_0/N_11_i_0 ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB11_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/rd_enable_net_1 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB1_rgbl_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/temp_data[3]_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_9_[4]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[4] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB13_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_9__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_183_i ), .ADn(VCC), .SLn(
        VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_9_rs[4] ));
    CFG4 #( .INIT(16'hB383) )  \CoreGPIO_0/CONFIG_reg_o_2_31_am[0]  (
        .A(\CoreGPIO_0/CONFIG_reg_o_2_31_am_RNO[0]_net_1 ), .B(
        \CoreGPIO_0/CONFIG_reg_o_2_31_am_1[0] ), .C(
        \CoreAPB3_0_APBmslave3_PADDR[3] ), .D(
        \CoreGPIO_0/CONFIG_reg_o_2_31_am_RNO_0[0]_net_1 ), .Y(
        \CoreGPIO_0/CONFIG_reg_o_2_31_am[0]_net_1 ));
    CFG2 #( .INIT(4'h7) )  \CoreGPIO_0/edge_both_2_sqmuxa_28_i  (.A(
        \CoreGPIO_0/N_248 ), .B(\CoreGPIO_0/CONFIG_reg[27][3] ), .Y(
        \CoreGPIO_0/N_161 ));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_18_set_RNI9K6V  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_18_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_226_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_12_rs[2] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_12_[2]_net_1 ));
    CFG4 #( .INIT(16'hC5CA) )  
        \CoreGPIO_0/xhdl1.GEN_BITS[1].APB_32.INTR_reg_22_0_m2[1]  (.A(
        \CoreGPIO_0.xhdl1.GEN_BITS[1].gpin3[1] ), .B(
        \CoreGPIO_0/N_174 ), .C(\CoreGPIO_0/CONFIG_reg[1][6] ), .D(
        \CoreGPIO_0/CONFIG_reg[1][5] ), .Y(\CoreGPIO_0/N_177 ));
    sdf_IOPAD_IN \GPIO_IN_ibuf[5]/U0/U_IOPAD  (.PAD(GPIO_IN[5]), .Y(
        \GPIO_IN_ibuf[5]/U0/YIN1 ));
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_58  (
        .A(\reg_apb_wrp_0/reg16x8_0/mem_15_[4]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_497 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_58_net_1 ));
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_62  (
        .A(\reg_apb_wrp_0/reg16x8_0/mem_15_[5]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_497 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_62_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_17_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB2_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_12__1_sqmuxa ), .ALn(
        AFLSDF_INV_112_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_17_set_net_1 ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_111  (.A(VCC), 
        .B(VCC), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/FAB_XDATAIN_net[3] ), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/FAB_VSTATUS_net[0] ), .IPC());
    CFG2 #( .INIT(4'h4) )  \CoreGPIO_0/PRDATA_0_iv_0_a2_0[27]  (.A(
        \CoreGPIO_0.N_247 ), .B(\CoreGPIO_0/INTR_reg[27] ), .Y(
        \CoreGPIO_0.N_532 ));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_5_[5]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[5] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB5_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_5__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_182_i ), .ADn(VCC), .SLn(
        VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_5_rs[5] ));
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_22  (
        .A(\reg_apb_wrp_0/reg16x8_0/mem_12_[6]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_495 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_22_net_1 ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_273  (.A(GND), 
        .B(VCC), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/F_ARLEN_HBURST1_net[1] ), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PSEL_net ), .IPC());
    IOTRI_OB_EB \FIC_MSS_0/MDDR_CS_N_PAD/U_IOOUT  (.D(VCC), .E(VCC), 
        .DOUT(), .EOUT(\FIC_MSS_0/MDDR_CS_N_PAD/EOUT ));
    CFG4 #( .INIT(16'h4000) )  
        \CoreGPIO_0/xhdl1.GEN_BITS[1].REG_GEN.CONFIG_reg[1]2_0_a4_0_a2  
        (.A(\CoreAPB3_0_APBmslave3_PADDR[3] ), .B(
        \CoreAPB3_0_APBmslave3_PADDR[2] ), .C(\CoreGPIO_0/N_604 ), .D(
        \CoreGPIO_0/N_606 ), .Y(\CoreGPIO_0/CONFIG_reg[1]2 ));
    CFG3 #( .INIT(8'hF2) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_139  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_1_[3]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_502 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_139_i ));
    CFG3 #( .INIT(8'h08) )  
        \CoreGPIO_0/xhdl1.GEN_BITS[16].REG_GEN.CONFIG_reg[16]2_0_a4_0_a2_1  
        (.A(\CoreAPB3_0_APBmslave3_PADDR[6] ), .B(
        \CoreGPIO_0/INTR_reg21 ), .C(\CoreAPB3_0_APBmslave3_PADDR[7] ), 
        .Y(\CoreGPIO_0/N_598 ));
    CFG2 #( .INIT(4'h8) )  
        \reg_apb_wrp_0/reg16x8_0/mem_7__1_sqmuxa_0_a3  (.A(
        \reg_apb_wrp_0/reg16x8_0/N_498 ), .B(
        \reg_apb_wrp_0/wr_enable_net_1 ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_7__1_sqmuxa ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_85_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB19_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_0__1_sqmuxa ), .ALn(
        AFLSDF_INV_113_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_85_set_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_10_[2]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[2] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB14_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_10__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_195_i ), .ADn(VCC), .SLn(
        VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_10_rs[2] ));
    CCC #( .INIT(210'h0000007FB8000044D64000307C6318C6318C61EC0404040400301)
        , .VCOFREQUENCY(800.0) )  \FCCC_0/CCC_INST/INST_CCC_IP  (.Y0(), 
        .Y1(), .Y2(), .Y3(), .PRDATA({nc271, nc272, nc273, nc274, 
        nc275, nc276, nc277, nc278}), .LOCK(FCCC_0_LOCK), .BUSY(), 
        .CLK0(\FCCC_0/CCC_INST/CLK0_net ), .CLK1(
        \FCCC_0/CCC_INST/CLK1_net ), .CLK2(\FCCC_0/CCC_INST/CLK2_net ), 
        .CLK3(\FCCC_0/CCC_INST/CLK3_net ), .NGMUX0_SEL(
        \FCCC_0/CCC_INST/NGMUX0_SEL_net ), .NGMUX1_SEL(
        \FCCC_0/CCC_INST/NGMUX1_SEL_net ), .NGMUX2_SEL(
        \FCCC_0/CCC_INST/NGMUX2_SEL_net ), .NGMUX3_SEL(
        \FCCC_0/CCC_INST/NGMUX3_SEL_net ), .NGMUX0_HOLD_N(
        \FCCC_0/CCC_INST/NGMUX0_HOLD_N_net ), .NGMUX1_HOLD_N(
        \FCCC_0/CCC_INST/NGMUX1_HOLD_N_net ), .NGMUX2_HOLD_N(
        \FCCC_0/CCC_INST/NGMUX2_HOLD_N_net ), .NGMUX3_HOLD_N(
        \FCCC_0/CCC_INST/NGMUX3_HOLD_N_net ), .NGMUX0_ARST_N(
        \FCCC_0/CCC_INST/NGMUX0_ARST_N_net ), .NGMUX1_ARST_N(
        \FCCC_0/CCC_INST/NGMUX1_ARST_N_net ), .NGMUX2_ARST_N(
        \FCCC_0/CCC_INST/NGMUX2_ARST_N_net ), .NGMUX3_ARST_N(
        \FCCC_0/CCC_INST/NGMUX3_ARST_N_net ), .PLL_BYPASS_N(
        \FCCC_0/CCC_INST/PLL_BYPASS_N_net ), .PLL_ARST_N(
        \FCCC_0/CCC_INST/PLL_ARST_N_net ), .PLL_POWERDOWN_N(
        \FCCC_0/CCC_INST/PLL_POWERDOWN_N_net ), .GPD0_ARST_N(
        \FCCC_0/CCC_INST/GPD0_ARST_N_net ), .GPD1_ARST_N(
        \FCCC_0/CCC_INST/GPD1_ARST_N_net ), .GPD2_ARST_N(
        \FCCC_0/CCC_INST/GPD2_ARST_N_net ), .GPD3_ARST_N(
        \FCCC_0/CCC_INST/GPD3_ARST_N_net ), .PRESET_N(
        \FCCC_0/CCC_INST/PRESET_N_net ), .PCLK(
        \FCCC_0/CCC_INST/PCLK_net ), .PSEL(\FCCC_0/CCC_INST/PSEL_net ), 
        .PENABLE(\FCCC_0/CCC_INST/PENABLE_net ), .PWRITE(
        \FCCC_0/CCC_INST/PWRITE_net ), .PADDR({
        \FCCC_0/CCC_INST/PADDR_net[7] , \FCCC_0/CCC_INST/PADDR_net[6] , 
        \FCCC_0/CCC_INST/PADDR_net[5] , \FCCC_0/CCC_INST/PADDR_net[4] , 
        \FCCC_0/CCC_INST/PADDR_net[3] , \FCCC_0/CCC_INST/PADDR_net[2] })
        , .PWDATA({\FCCC_0/CCC_INST/PWDATA_net[7] , 
        \FCCC_0/CCC_INST/PWDATA_net[6] , 
        \FCCC_0/CCC_INST/PWDATA_net[5] , 
        \FCCC_0/CCC_INST/PWDATA_net[4] , 
        \FCCC_0/CCC_INST/PWDATA_net[3] , 
        \FCCC_0/CCC_INST/PWDATA_net[2] , 
        \FCCC_0/CCC_INST/PWDATA_net[1] , 
        \FCCC_0/CCC_INST/PWDATA_net[0] }), .CLK0_PAD(GND), .CLK1_PAD(
        GND), .CLK2_PAD(GND), .CLK3_PAD(GND), .GL0(), .GL1(), .GL2(), 
        .GL3(\FCCC_0/GL1_net ), .RCOSC_25_50MHZ(
        OSC_0_RCOSC_25_50MHZ_CCC_OUT_RCOSC_25_50MHZ_CCC), .RCOSC_1MHZ(
        GND), .XTLOSC(GND));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[5].gpin2[5]  (.D(
        \CoreGPIO_0/gpin1[5] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB10_rgbr_net_1 ), .EN(VCC), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB0_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(\CoreGPIO_0/gpin2[5] )
        );
    IOTRI_OB_EB \FIC_MSS_0/MDDR_ADDR_13_PAD/U_IOOUT  (.D(VCC), .E(VCC), 
        .DOUT(), .EOUT(\FIC_MSS_0/MDDR_ADDR_13_PAD/EOUT ));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/mem_10__RNIH13P[1]  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_98_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_193_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_10_rs[1] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_10_[1]_net_1 ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[16].REG_GEN.CONFIG_reg[16][1]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[1] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB15_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[16]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB5_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[16][1] ));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_78_set_RNIFTT11  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_78_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_187_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_9_rs[6] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_9_[6]_net_1 ));
    IOTRI_OB_EB \FIC_MSS_0/MDDR_ADDR_12_PAD/U_IOOUT  (.D(VCC), .E(VCC), 
        .DOUT(), .EOUT(\FIC_MSS_0/MDDR_ADDR_12_PAD/EOUT ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_104_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB11_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_13__1_sqmuxa ), .ALn(
        AFLSDF_INV_114_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_104_set_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_12_[0]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[0] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB1_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_12__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_222_i ), .ADn(VCC), .SLn(
        VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_12_rs[0] ));
    IP_INTERFACE \FCCC_0/CCC_INST/IP_INTERFACE_11  (.A(VCC), .B(VCC), 
        .C(VCC), .IPA(\FCCC_0/CCC_INST/PLL_POWERDOWN_N_net ), .IPB(
        \FCCC_0/CCC_INST/NGMUX3_HOLD_N_net ), .IPC());
    CFG4 #( .INIT(16'h1000) )  
        \CoreGPIO_0/xhdl1.GEN_BITS[24].REG_GEN.CONFIG_reg[24]2_0_a4_0_a2  
        (.A(\CoreAPB3_0_APBmslave3_PADDR[3] ), .B(
        \CoreAPB3_0_APBmslave3_PADDR[2] ), .C(\CoreGPIO_0/N_598 ), .D(
        \CoreGPIO_0/N_610 ), .Y(\CoreGPIO_0/CONFIG_reg[24]2 ));
    INV_BA AFLSDF_INV_78 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_117_net_1 ), .Y(
        AFLSDF_INV_78_net_1));
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_5  (
        .A(\reg_apb_wrp_0/reg16x8_0/mem_8_[1]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_499 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_5_net_1 ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_126  (.A(GND), 
        .B(GND), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[1] ), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[8] ), .IPC());
    CFG3 #( .INIT(8'hF2) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_130  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_0_[3]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_496 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_130_i ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[19].REG_GEN.CONFIG_reg[19][6]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[6] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB9_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[19]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_YR ), .ADn(VCC), .SLn(
        VCC), .SD(GND), .LAT(GND), .Q(\CoreGPIO_0/CONFIG_reg[19][6] ));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/mem_11__RNICVCQ[7]  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_95_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_220_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_11_rs[7] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_11_[7]_net_1 ));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/mem_3__RNIU02R[3]  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_48_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_155_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_3_rs[3] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_3_[3]_net_1 ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[1].REG_GEN.CONFIG_reg[1][4]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[4] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB14_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[1]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB4_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[1][4] ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_169  (.A(VCC), 
        .B(VCC), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/MMUART1_DSR_F2H_SCP_net ), .IPB(), 
        .IPC());
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_165  (.A(VCC), 
        .B(VCC), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/SPI1_SS0_F2H_SCP_net ), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/SPI1_SS3_F2H_SCP_net ), .IPC());
    CFG3 #( .INIT(8'hF2) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_209  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_11_[1]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_505 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_209_i ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_72  (.A(VCC), 
        .B(VCC), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[6] ), .IPB(), 
        .IPC());
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[4].REG_GEN.CONFIG_reg[4][3]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[3] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB12_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[4]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB2_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[4][3] ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_6_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB9_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_4__1_sqmuxa ), .ALn(
        AFLSDF_INV_115_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_6_set_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_13_[5]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[5] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB5_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_13__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_237_i ), .ADn(VCC), .SLn(
        VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_13_rs[5] ));
    IOBI_IB_OB_EB \FIC_MSS_0/MDDR_DQ_13_PAD/U_IOBI  (.D(VCC), .E(VCC), 
        .YIN(\FIC_MSS_0/MDDR_DQ_13_PAD/YIN ), .DOUT(), .EOUT(), .Y());
    CFG3 #( .INIT(8'hF2) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_135  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_0_[7]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_496 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_135_i ));
    CFG4 #( .INIT(16'h7350) )  
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_5[0]  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_14_[0]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/mem_6_[0]_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/N_503 ), .D(
        \reg_apb_wrp_0/reg16x8_0/N_493 ), .Y(
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_5[0]_net_1 ));
    sdf_IOPAD_TRI \FIC_MSS_0/MDDR_ADDR_13_PAD/U_IOPAD  (.PAD(
        MDDR_ADDR[13]), .D(\FIC_MSS_0/DRAM_ADDR_net_0[13] ), .E(
        \FIC_MSS_0/MDDR_ADDR_13_PAD/EOUT ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[19].APB_32.edge_both[19]  (.D(
        \CoreGPIO_0/edge_neg_275[19] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB9_rgbr_net_1 ), .EN(
        \CoreGPIO_0/N_194 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_YR ), .ADn(VCC), .SLn(
        VCC), .SD(GND), .LAT(GND), .Q(\CoreGPIO_0/edge_neg[19] ));
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_40  (
        .A(\reg_apb_wrp_0/reg16x8_0/mem_5_[2]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_490 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_40_net_1 ));
    INV_BA AFLSDF_INV_52 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_127_net_1 ), .Y(
        AFLSDF_INV_52_net_1));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_188  (.A(VCC), 
        .B(VCC), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/MGPIO30B_F2H_GPIN_net ), .IPB(), 
        .IPC());
    CFG4 #( .INIT(16'hEC00) )  \CoreAPB3_0/u_mux_p_to_b3/PRDATA[11]  (
        .A(\CoreGPIO_0.xhdl1.GEN_BITS[0].APB_32.GPOUT_reg9 ), .B(
        \CoreGPIO_0.N_564 ), .C(
        \CoreGPIO_0.xhdl1.GEN_BITS[11].APB_32.GPOUT_reg[11] ), .D(
        CoreAPB3_0_APBmslave5_PSELx), .Y(
        \FIC_MSS_0_FIC_0_APB_MASTER_PRDATA[11] ));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_5_[7]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[7] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB9_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_5__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_186_i ), .ADn(VCC), .SLn(
        VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_5_rs[7] ));
    RGB \FCCC_0/GL1_INST/U0_RGB1_RGB4  (.An(\FCCC_0/GL1_INST/U0_YNn ), 
        .ENn(GND), .YL(\FCCC_0/GL1_INST/U0_RGB1_RGB4_rgbl_net_1 ), .YR(
        \FCCC_0/GL1_INST/U0_RGB1_RGB4_rgbr_net_1 ));
    CFG2 #( .INIT(4'h2) )  
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_a3_5[2]  (.A(
        \reg_apb_wrp_0/reg16x8_0/N_495 ), .B(
        \reg_apb_wrp_0/reg16x8_0/mem_12_[2]_net_1 ), .Y(
        \reg_apb_wrp_0/reg16x8_0/N_392 ));
    CFG2 #( .INIT(4'h4) )  \CoreGPIO_0/PRDATA_0_iv_0_a2_0[22]  (.A(
        \CoreGPIO_0.N_247 ), .B(\CoreGPIO_0/INTR_reg[22] ), .Y(
        \CoreGPIO_0.N_542 ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_254_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_62_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_254_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_254_rs_net_1 ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[2].REG_GEN.CONFIG_reg[2][0]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[0] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB16_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[2]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB6_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[2][0] ));
    INV_BA AFLSDF_INV_15 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_38_net_1 ), .Y(
        AFLSDF_INV_15_net_1));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_13_[4]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[4] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB5_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_13__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_236_i ), .ADn(VCC), .SLn(
        VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_13_rs[4] ));
    SLE \reg_apb_wrp_0/PREADY  (.D(\reg_apb_wrp_0/N_64_i_0 ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB12_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/N_44_i_0 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB2_rgbr_net_1 ), .ADn(
        GND), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        CoreAPB3_0_APBmslave3_PREADY));
    IOBI_IB_OB_EB \FIC_MSS_0/MDDR_DQ_0_PAD/U_IOBI  (.D(VCC), .E(VCC), 
        .YIN(\FIC_MSS_0/MDDR_DQ_0_PAD/YIN ), .DOUT(), .EOUT(), .Y());
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[10].REG_GEN.CONFIG_reg[10][2]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[2] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB16_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[10]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB6_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[10][2] ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_189_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_79_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_189_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_189_rs_net_1 ));
    CFG3 #( .INIT(8'hF2) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_148  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_2_[4]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_501 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_148_i ));
    IP_INTERFACE \FCCC_0/CCC_INST/IP_INTERFACE_14  (.A(VCC), .B(VCC), 
        .C(VCC), .IPA(\FCCC_0/CCC_INST/NGMUX2_ARST_N_net ), .IPB(
        \FCCC_0/CCC_INST/GPD0_ARST_N_net ), .IPC(
        \FCCC_0/CCC_INST/PADDR_net[4] ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_221  (.A(VCC), 
        .B(VCC), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[5] ), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[17] ), .IPC());
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_64_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB14_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_8__1_sqmuxa ), .ALn(
        AFLSDF_INV_116_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_64_set_net_1 ));
    CFG4 #( .INIT(16'hA9FF) )  
        \CoreGPIO_0/xhdl1.GEN_BITS[25].APB_32.INTR_reg_334_0_o2_0_0[25]  
        (.A(\CoreGPIO_0/CONFIG_reg[25][7] ), .B(
        \CoreGPIO_0/CONFIG_reg[25][6] ), .C(
        \CoreGPIO_0/CONFIG_reg[25][5] ), .D(
        \CoreGPIO_0/CONFIG_reg[25][3] ), .Y(
        \CoreGPIO_0/INTR_reg_334_0_o2_0[25] ));
    CFG4 #( .INIT(16'hF2F3) )  
        \CoreGPIO_0/xhdl1.GEN_BITS[14].APB_32.INTR_reg_191_0_o2_1_0[14]  
        (.A(\CoreGPIO_0/CONFIG_reg[14][6] ), .B(
        \CoreGPIO_0/edge_neg[14] ), .C(
        \CoreGPIO_0/INTR_reg_191_0_o2_0[14] ), .D(
        \CoreGPIO_0/CONFIG_reg[14][5] ), .Y(
        \CoreGPIO_0/INTR_reg_191_0_o2_1[14] ));
    INV_BA AFLSDF_INV_103 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_19_net_1 ), .Y(
        AFLSDF_INV_103_net_1));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_63  (.A(GND), 
        .B(GND), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[24] ), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[31] ), .IPC());
    CFG2 #( .INIT(4'h8) )  
        \CoreGPIO_0/xhdl1.GEN_BITS[0].REG_GPOUT.un5_GPIO_OUT_i  (.A(
        \CoreGPIO_0/GPOUT_reg[0] ), .B(\CoreGPIO_0/CONFIG_reg[0][0] ), 
        .Y(\GPIO_OUT_net_2[0] ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_16  (.A(
        \FIC_MSS_0_FIC_0_APB_MASTER_PRDATA[21] ), .B(
        \FIC_MSS_0_FIC_0_APB_MASTER_PRDATA[28] ), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[21] ), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[28] ), .IPC());
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/mem_6__RNI3P1N[0]  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_29_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_188_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_6_rs[0] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_6_[0]_net_1 ));
    CFG4 #( .INIT(16'h7350) )  
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_6[1]  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_8_[1]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/mem_0_[1]_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/N_499 ), .D(
        \reg_apb_wrp_0/reg16x8_0/N_496 ), .Y(
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_6[1]_net_1 ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_123  (.A(VCC), 
        .B(GND), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/FAB_HOSTDISCON_net ), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[5] ), .IPC());
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[6].REG_GEN.CONFIG_reg[6][5]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[5] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB12_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[6]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB2_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[6][5] ));
    CFG2 #( .INIT(4'h6) )  \CoreGPIO_0/edge_both_2_sqmuxa_23_i_x2  (.A(
        \CoreGPIO_0/gpin2[5] ), .B(
        \CoreGPIO_0.xhdl1.GEN_BITS[5].gpin3[5] ), .Y(
        \CoreGPIO_0/N_139_i ));
    CFG4 #( .INIT(16'hAC0F) )  
        \CoreGPIO_0/CONFIG_reg_o_2_31_bm_RNO[1]  (.A(
        \CoreGPIO_0/CONFIG_reg[11][1] ), .B(
        \CoreGPIO_0/CONFIG_reg[27][1] ), .C(
        \CoreGPIO_0/CONFIG_reg_o_2_25_1_1[1] ), .D(
        \CoreAPB3_0_APBmslave3_PADDR[5] ), .Y(
        \CoreGPIO_0/CONFIG_reg_o_2_31_bm_RNO[1]_net_1 ));
    CFG4 #( .INIT(16'h0F35) )  
        \CoreGPIO_0/CONFIG_reg_o_2_31_bm_RNO_2[2]  (.A(
        \CoreGPIO_0/CONFIG_reg[7][2] ), .B(
        \CoreGPIO_0/CONFIG_reg[23][2] ), .C(
        \CoreAPB3_0_APBmslave3_PADDR[6] ), .D(
        \CoreAPB3_0_APBmslave3_PADDR[5] ), .Y(
        \CoreGPIO_0/CONFIG_reg_o_2_28_1_1[2] ));
    CFG4 #( .INIT(16'hA9FF) )  
        \CoreGPIO_0/xhdl1.GEN_BITS[18].APB_32.INTR_reg_243_0_o2_0_0[18]  
        (.A(\CoreGPIO_0/CONFIG_reg[18][7] ), .B(
        \CoreGPIO_0/CONFIG_reg[18][6] ), .C(
        \CoreGPIO_0/CONFIG_reg[18][5] ), .D(
        \CoreGPIO_0/CONFIG_reg[18][3] ), .Y(
        \CoreGPIO_0/INTR_reg_243_0_o2_0[18] ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[0].REG_GEN.CONFIG_reg[0][1]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[1] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB15_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[0]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB5_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0.xhdl1.GEN_BITS[0].REG_GEN.CONFIG_reg[0][1] ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[27].REG_GEN.CONFIG_reg[27][3]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[3] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB9_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[27]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_YR ), .ADn(VCC), .SLn(
        VCC), .SD(GND), .LAT(GND), .Q(\CoreGPIO_0/CONFIG_reg[27][3] ));
    sdf_IOPAD_TRI \FIC_MSS_0/MMUART_0_TXD_PAD/U_IOPAD  (.PAD(
        MMUART_0_TXD), .D(
        \FIC_MSS_0/MSS_ADLIB_INST_MMUART0_TXD_USBC_DIR_MGPIO27B_OUT ), 
        .E(\FIC_MSS_0/MSS_ADLIB_INST_MMUART0_TXD_USBC_DIR_MGPIO27B_OE )
        );
    IOBI_IB_OB_EB \FIC_MSS_0/MDDR_DQ_11_PAD/U_IOBI  (.D(VCC), .E(VCC), 
        .YIN(\FIC_MSS_0/MDDR_DQ_11_PAD/YIN ), .DOUT(), .EOUT(), .Y());
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_92_set_RNI9O0E  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_92_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_214_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_11_rs[4] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_11_[4]_net_1 ));
    CFG2 #( .INIT(4'h8) )  
        \CoreGPIO_0/xhdl1.GEN_BITS[14].REG_GEN.CONFIG_reg[14]2_0_a4_0_a2_0  
        (.A(\CoreAPB3_0_APBmslave3_PADDR[5] ), .B(
        \CoreAPB3_0_APBmslave3_PADDR[4] ), .Y(\CoreGPIO_0/N_605 ));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_9_[2]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[2] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB15_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_9__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_179_i ), .ADn(VCC), .SLn(
        VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_9_rs[2] ));
    CFG3 #( .INIT(8'hB8) )  
        \CoreGPIO_0/xhdl1.GEN_BITS[5].APB_32.INTR_reg_74_0_m2_0_i_m2[5]  
        (.A(\CoreGPIO_0/edge_neg[5] ), .B(
        \CoreGPIO_0/CONFIG_reg[5][5] ), .C(\CoreGPIO_0/edge_pos[5] ), 
        .Y(\CoreGPIO_0/N_171 ));
    CFG4 #( .INIT(16'hAC0F) )  
        \CoreGPIO_0/CONFIG_reg_o_2_31_am_1_1_RNO[5]  (.A(
        \CoreGPIO_0/CONFIG_reg[12][5] ), .B(
        \CoreGPIO_0/CONFIG_reg[28][5] ), .C(
        \CoreGPIO_0/CONFIG_reg_o_2_6_1[5] ), .D(
        \CoreAPB3_0_APBmslave3_PADDR[5] ), .Y(
        \CoreGPIO_0/CONFIG_reg_o_2_31_am_1_1_RNO[5]_net_1 ));
    sdf_IOPAD_IN \GPIO_IN_ibuf[3]/U0/U_IOPAD  (.PAD(GPIO_IN[3]), .Y(
        \GPIO_IN_ibuf[3]/U0/YIN1 ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[5].REG_GEN.CONFIG_reg[5][5]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[5] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB13_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[5]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB3_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[5][5] ));
    CFG4 #( .INIT(16'h0F35) )  
        \CoreGPIO_0/CONFIG_reg_o_2_31_bm_1_RNO_2[0]  (.A(
        \CoreGPIO_0/CONFIG_reg[1][0] ), .B(
        \CoreGPIO_0/CONFIG_reg[17][0] ), .C(
        \CoreAPB3_0_APBmslave3_PADDR[6] ), .D(
        \CoreAPB3_0_APBmslave3_PADDR[5] ), .Y(
        \CoreGPIO_0/CONFIG_reg_o_2_18_1[0] ));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_137_rs_RNIHDC41  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_12_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_137_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_1_rs[1] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_1_[1]_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_98_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB2_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_10__1_sqmuxa ), .ALn(
        AFLSDF_INV_117_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_98_set_net_1 ));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/mem_14__RNI2R8D[6]  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_118_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_246_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_14_rs[6] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_14_[6]_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/data_out[5]  (.D(
        \reg_apb_wrp_0/reg16x8_0/temp_data[5]_net_1 ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB10_rgbr_net_1 ), .EN(VCC), .ALn(
        VCC), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreAPB3_0_APBmslave3_PRDATA[5] ));
    CFG2 #( .INIT(4'h7) )  \CoreGPIO_0/edge_both_2_sqmuxa_6_i  (.A(
        \CoreGPIO_0/N_248 ), .B(\CoreGPIO_0/CONFIG_reg[22][3] ), .Y(
        \CoreGPIO_0/N_200 ));
    CFG4 #( .INIT(16'h0080) )  
        \reg_apb_wrp_0/reg16x8_0/WRITE_GEN.mem_13__2_i_0_0_a2[5]  (.A(
        \CoreAPB3_0_APBmslave3_PADDR[3] ), .B(
        \CoreAPB3_0_APBmslave3_PADDR[2] ), .C(
        \CoreAPB3_0_APBmslave3_PADDR[0] ), .D(
        \CoreAPB3_0_APBmslave3_PADDR[1] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/N_500 ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_184  (.A(VCC), 
        .B(VCC), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/MGPIO28B_F2H_GPIN_net ), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/MGPIO31B_F2H_GPIN_net ), .IPC());
    CFG4 #( .INIT(16'hF2F3) )  
        \CoreGPIO_0/xhdl1.GEN_BITS[13].APB_32.INTR_reg_178_0_o2_1_0[13]  
        (.A(\CoreGPIO_0/CONFIG_reg[13][6] ), .B(
        \CoreGPIO_0/edge_neg[13] ), .C(
        \CoreGPIO_0/INTR_reg_178_0_o2_0[13] ), .D(
        \CoreGPIO_0/CONFIG_reg[13][5] ), .Y(
        \CoreGPIO_0/INTR_reg_178_0_o2_1[13] ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_26_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB1_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_2__1_sqmuxa ), .ALn(
        AFLSDF_INV_118_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_26_set_net_1 ));
    INV_BA AFLSDF_INV_94 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_11_net_1 ), .Y(
        AFLSDF_INV_94_net_1));
    CFG3 #( .INIT(8'hF2) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_240  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_14_[0]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_503 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_240_i ));
    IP_INTERFACE \FCCC_0/CCC_INST/IP_INTERFACE_15  (.A(VCC), .B(VCC), 
        .C(VCC), .IPA(\FCCC_0/CCC_INST/NGMUX3_ARST_N_net ), .IPB(
        \FCCC_0/CCC_INST/GPD1_ARST_N_net ), .IPC(
        \FCCC_0/CCC_INST/PADDR_net[5] ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[25].REG_GEN.CONFIG_reg[25][2]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[2] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB16_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[25]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB6_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[25][2] ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_161_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_net_1 ), .EN(VCC), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_161_i ), .ADn(VCC), .SLn(
        VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_161_rs_net_1 ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_91  (.A(VCC), 
        .B(VCC), .C(VCC), .IPA(\FIC_MSS_0/MSS_ADLIB_INST/TX_CLKPF_net )
        , .IPB(\FIC_MSS_0/MSS_ADLIB_INST/RXDF_net[7] ), .IPC());
    CFG3 #( .INIT(8'h04) )  
        \CoreGPIO_0/xhdl1.GEN_BITS[1].APB_32.INTR_reg_22_0_0_RNO_0[1]  
        (.A(\CoreGPIO_0/CONFIG_reg[1][5] ), .B(
        \CoreGPIO_0/edge_both[1] ), .C(\CoreGPIO_0/CONFIG_reg[1][6] ), 
        .Y(\CoreGPIO_0/INTR_reg_22_0_0_51_tz_1 ));
    CFG4 #( .INIT(16'hDC00) )  \CoreAPB3_0/u_mux_p_to_b3/PRDATA[18]  (
        .A(\CoreGPIO_0.N_247 ), .B(\CoreGPIO_0.N_549 ), .C(
        \CoreGPIO_0.xhdl1.GEN_BITS[18].APB_32.INTR_reg[18] ), .D(
        CoreAPB3_0_APBmslave5_PSELx), .Y(
        \FIC_MSS_0_FIC_0_APB_MASTER_PRDATA[18] ));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_4_[3]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[3] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB9_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_4__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_164_i ), .ADn(VCC), .SLn(
        VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_4_rs[3] ));
    CFG3 #( .INIT(8'hF2) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_242  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_14_[2]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_503 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_242_i ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[4].APB_32.edge_both[4]  (.D(
        \CoreGPIO_0/N_91 ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB13_rgbr_net_1 ), .EN(
        \CoreGPIO_0/N_84 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB3_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/edge_both[4] ));
    CFG4 #( .INIT(16'h330A) )  
        \CoreGPIO_0/xhdl1.GEN_BITS[11].APB_32.INTR_reg_152_0[11]  (.A(
        \CoreGPIO_0/INTR_reg[11] ), .B(
        \CoreGPIO_0/INTR_reg_152_0_o2_1[11] ), .C(
        \CoreAPB3_0_APBmslave3_PWDATA[11] ), .D(\CoreGPIO_0/N_248 ), 
        .Y(\CoreGPIO_0/INTR_reg_152[11] ));
    sdf_IOPADN_BI \FIC_MSS_0/MDDR_DQS_1_PAD/U_IOPADN  (.PAD_P(
        MDDR_DQS_N[1]), .OIN_P(\FIC_MSS_0/DRAM_DQS_OUT_net_0[1] ), 
        .EIN_P(\FIC_MSS_0/DRAM_DQS_OE_net_0[1] ), .N2POUT_P(
        \FIC_MSS_0/MDDR_DQS_1_PAD/U2_N2P ));
    CFG4 #( .INIT(16'hB383) )  \CoreGPIO_0/CONFIG_reg_o_2_31_am[4]  (
        .A(\CoreGPIO_0/CONFIG_reg_o_2_31_am_RNO[4]_net_1 ), .B(
        \CoreGPIO_0/CONFIG_reg_o_2_31_am_1[4] ), .C(
        \CoreAPB3_0_APBmslave3_PADDR[3] ), .D(
        \CoreGPIO_0/CONFIG_reg_o_2_31_am_RNO_0[4]_net_1 ), .Y(
        \CoreGPIO_0/CONFIG_reg_o_2_31_am[4]_net_1 ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_35  (.A(VCC), 
        .B(GND), .C(VCC), .IPA(), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[18] ), .IPC());
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[20].REG_GEN.CONFIG_reg[20][6]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[6] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB12_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[20]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB2_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[20][6] ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_162_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_2_net_1 ), .EN(VCC), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_162_i ), .ADn(VCC), .SLn(
        VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_162_rs_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/data_out[3]  (.D(
        \reg_apb_wrp_0/reg16x8_0/temp_data[3]_net_1 ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB12_rgbr_net_1 ), .EN(VCC), .ALn(
        VCC), .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreAPB3_0_APBmslave3_PRDATA[3] ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_10_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB14_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_1__1_sqmuxa ), .ALn(
        AFLSDF_INV_119_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_10_set_net_1 ));
    sdf_IOPAD_TRI \FIC_MSS_0/MDDR_WE_N_PAD/U_IOPAD  (.PAD(MDDR_WE_N), 
        .D(\FIC_MSS_0/MSS_ADLIB_INST_DRAM_WEN ), .E(
        \FIC_MSS_0/MDDR_WE_N_PAD/EOUT ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[6].APB_32.INTR_reg[6]  (.D(
        \CoreGPIO_0/INTR_reg_87[6] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB12_rgbr_net_1 ), .EN(VCC), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB2_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0.xhdl1.GEN_BITS[6].APB_32.INTR_reg[6] ));
    CFG4 #( .INIT(16'hEC00) )  \CoreAPB3_0/u_mux_p_to_b3/PRDATA[14]  (
        .A(\CoreGPIO_0.xhdl1.GEN_BITS[0].APB_32.GPOUT_reg9 ), .B(
        \CoreGPIO_0.N_558 ), .C(
        \CoreGPIO_0.xhdl1.GEN_BITS[14].APB_32.GPOUT_reg[14] ), .D(
        CoreAPB3_0_APBmslave5_PSELx), .Y(
        \FIC_MSS_0_FIC_0_APB_MASTER_PRDATA[14] ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_175_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_72_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_175_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_175_rs_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_0_[6]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[6] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB17_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_0__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_134_i ), .ADn(VCC), .SLn(
        VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_0_rs[6] ));
    sdf_IOPAD_IN \MSS_RESET_N_F2M_ibuf/U0/U_IOPAD  (.PAD(
        MSS_RESET_N_F2M), .Y(\MSS_RESET_N_F2M_ibuf/U0/YIN1 ));
    CFG3 #( .INIT(8'hF2) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_143  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_1_[7]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_502 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_143_i ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[0].APB_32.GPOUT_reg[0]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[0] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB11_rgbr_net_1 ), .EN(
        \CoreGPIO_0/GPOUT_reg_0_sqmuxa ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB1_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/GPOUT_reg[0] ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_249_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_59_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_249_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_249_rs_net_1 ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_283  (.A(VCC), 
        .B(VCC), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PADDR_net[6] ), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[10] ), .IPC());
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_24_set_RNINOSM  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_24_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_143_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_1_rs[7] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_1_[7]_net_1 ));
    IOTRI_OB_EB \GPIO_OUT_obuf[4]/U0/U_IOTRI  (.D(\GPIO_OUT_net_2[4] ), 
        .E(VCC), .DOUT(\GPIO_OUT_obuf[4]/U0/DOUT1 ), .EOUT(
        \GPIO_OUT_obuf[4]/U0/EOUT1 ));
    CFG3 #( .INIT(8'h40) )  \CoreGPIO_0/PRDATA_iv_0_a2_0[3]  (.A(
        \CoreGPIO_0.N_246 ), .B(\CoreGPIO_0/GPOUT_reg[3] ), .C(
        \CoreAPB3_0_APBmslave3_PADDR[5] ), .Y(\CoreGPIO_0.N_496 ));
    CFG3 #( .INIT(8'h20) )  
        \CoreGPIO_0/xhdl1.GEN_BITS[31].APB_32.edge_both_RNO[31]  (.A(
        \CoreGPIO_0/CONFIG_reg[31][3] ), .B(
        \CoreAPB3_0_APBmslave3_PWDATA[31] ), .C(
        \CoreGPIO_0/edge_pos[31] ), .Y(\CoreGPIO_0/edge_neg_443[31] ));
    CFG4 #( .INIT(16'h0F35) )  
        \CoreGPIO_0/CONFIG_reg_o_2_31_am_1_RNO_2[3]  (.A(
        \CoreGPIO_0/CONFIG_reg[0][3] ), .B(
        \CoreGPIO_0/CONFIG_reg[16][3] ), .C(
        \CoreAPB3_0_APBmslave3_PADDR[6] ), .D(
        \CoreAPB3_0_APBmslave3_PADDR[5] ), .Y(
        \CoreGPIO_0/CONFIG_reg_o_2_3_1[3] ));
    CFG2 #( .INIT(4'h8) )  
        \reg_apb_wrp_0/reg16x8_0/mem_3__1_sqmuxa_0_a3  (.A(
        \reg_apb_wrp_0/reg16x8_0/N_494 ), .B(
        \reg_apb_wrp_0/wr_enable_net_1 ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_3__1_sqmuxa ));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_77_set_RNIBIHR  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_77_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_185_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_9_rs[5] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_9_[5]_net_1 ));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_89_set_RNIGNAI  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_89_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_209_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_11_rs[1] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_11_[1]_net_1 ));
    CFG4 #( .INIT(16'h8F88) )  \FIC_MSS_0/MSS_ADLIB_INST_RNO_12  (.A(
        \CoreAPB3_0_APBmslave3_PRDATA[6] ), .B(
        CoreAPB3_0_APBmslave3_PSELx), .C(\CoreGPIO_0.N_247 ), .D(
        \FIC_MSS_0/CoreAPB3_0_APBmslave5_PRDATA_m_c_c_0[6] ), .Y(
        \FIC_MSS_0/CoreAPB3_0_APBmslave5_PRDATA_m_0_0[6] ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[4].REG_GEN.CONFIG_reg[4][6]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[6] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB12_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[4]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB2_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[4][6] ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_228  (.A(VCC), 
        .B(VCC), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[26] ), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[38] ), .IPC(
        \FIC_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[50] ));
    CFG4 #( .INIT(16'h0F35) )  
        \CoreGPIO_0/CONFIG_reg_o_2_31_am_RNO_2[1]  (.A(
        \CoreGPIO_0.xhdl1.GEN_BITS[6].REG_GEN.CONFIG_reg[6][1] ), .B(
        \CoreGPIO_0/CONFIG_reg[22][1] ), .C(
        \CoreAPB3_0_APBmslave3_PADDR[6] ), .D(
        \CoreAPB3_0_APBmslave3_PADDR[5] ), .Y(
        \CoreGPIO_0/CONFIG_reg_o_2_13_1_1[1] ));
    CFG4 #( .INIT(16'h0F35) )  
        \CoreGPIO_0/CONFIG_reg_o_2_31_am_RNO_1[3]  (.A(
        \CoreGPIO_0/CONFIG_reg[2][3] ), .B(
        \CoreGPIO_0/CONFIG_reg[18][3] ), .C(
        \CoreAPB3_0_APBmslave3_PADDR[6] ), .D(
        \CoreAPB3_0_APBmslave3_PADDR[5] ), .Y(
        \CoreGPIO_0/CONFIG_reg_o_2_10_1_1[3] ));
    CFG3 #( .INIT(8'hF2) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_128  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_0_[1]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_496 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_128_i ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_211_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_90_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_211_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_211_rs_net_1 ));
    CFG4 #( .INIT(16'h7530) )  
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_7[4]  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_10_[4]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/mem_2_[4]_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/N_501 ), .D(
        \reg_apb_wrp_0/reg16x8_0/N_491 ), .Y(
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_7[4]_net_1 ));
    CFG4 #( .INIT(16'h7530) )  
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_1[0]  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_15_[0]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/mem_7_[0]_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/N_498 ), .D(
        \reg_apb_wrp_0/reg16x8_0/N_497 ), .Y(
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_1[0]_net_1 ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[25].REG_GEN.CONFIG_reg[25][0]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[0] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB16_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[25]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB6_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[25][0] ));
    CFG3 #( .INIT(8'hF2) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_141  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_1_[5]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_502 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_141_i ));
    CFG4 #( .INIT(16'hF2F3) )  
        \CoreGPIO_0/xhdl1.GEN_BITS[21].APB_32.INTR_reg_282_0_o2_1_0[21]  
        (.A(\CoreGPIO_0/CONFIG_reg[21][6] ), .B(
        \CoreGPIO_0/edge_neg[21] ), .C(
        \CoreGPIO_0/INTR_reg_282_0_o2_0[21] ), .D(
        \CoreGPIO_0/CONFIG_reg[21][5] ), .Y(
        \CoreGPIO_0/INTR_reg_282_0_o2_1[21] ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[16].REG_GEN.CONFIG_reg[16][6]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[6] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB11_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[16]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB1_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[16][6] ));
    sdf_IOPAD_TRI \FIC_MSS_0/MDDR_ADDR_0_PAD/U_IOPAD  (.PAD(
        MDDR_ADDR[0]), .D(\FIC_MSS_0/DRAM_ADDR_net_0[0] ), .E(
        \FIC_MSS_0/MDDR_ADDR_0_PAD/EOUT ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_270  (.A(VCC), 
        .B(GND), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[30] ), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/F_RREADY_net ), .IPC());
    IOTRI_OB_EB \FIC_MSS_0/MDDR_ADDR_7_PAD/U_IOOUT  (.D(VCC), .E(VCC), 
        .DOUT(), .EOUT(\FIC_MSS_0/MDDR_ADDR_7_PAD/EOUT ));
    RGB \FCCC_0/GL1_INST/U0_RGB1_RGB13  (.An(
        \FCCC_0/GL1_INST/U0_YNn_GSouth ), .ENn(GND), .YL(
        \FCCC_0/GL1_INST/U0_RGB1_RGB13_rgbl_net_1 ), .YR(
        \FCCC_0/GL1_INST/U0_RGB1_RGB13_rgbr_net_1 ));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_172_rs_RNIK1KK  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_13_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_172_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_5_rs[0] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_5_[0]_net_1 ));
    CFG3 #( .INIT(8'h04) )  
        \CoreGPIO_0/xhdl1.GEN_BITS[2].APB_32.INTR_reg_35_0_0_RNO_0[2]  
        (.A(\CoreGPIO_0/CONFIG_reg[2][5] ), .B(
        \CoreGPIO_0/edge_both[2] ), .C(\CoreGPIO_0/CONFIG_reg[2][6] ), 
        .Y(\CoreGPIO_0/INTR_reg_35_0_0_52_tz_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_13_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB11_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_5__1_sqmuxa ), .ALn(
        AFLSDF_INV_120_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_13_set_net_1 ));
    IOIN_IB \GPIO_IN_ibuf[1]/U0/U_IOIN  (.YIN(\GPIO_IN_ibuf[1]/U0/YIN )
        , .E(GND), .Y(\GPIO_IN_c[1] ));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_11_[1]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[1] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB16_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_11__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_209_i ), .ADn(VCC), .SLn(
        VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_11_rs[1] ));
    CFG2 #( .INIT(4'h2) )  \reg_apb_wrp_0/wr_enable_RNO  (.A(
        CoreAPB3_0_APBmslave3_PWRITE), .B(\reg_apb_wrp_0/fsm[0]_net_1 )
        , .Y(\reg_apb_wrp_0/N_70 ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_229_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_21_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_229_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_229_rs_net_1 ));
    CFG3 #( .INIT(8'h01) )  \reg_apb_wrp_0/reg16x8_0/temp_data_RNO[3]  
        (.A(\reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_8[3]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_13[3]_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_9[3]_net_1 ), .Y(
        \reg_apb_wrp_0/reg16x8_0/N_11_i_0 ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[3].REG_GEN.CONFIG_reg[3][4]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[4] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB10_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[3]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB0_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[3][4] ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_277  (.A(VCC), 
        .B(VCC), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[1] ), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[4] ), .IPC());
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[19].REG_GEN.CONFIG_reg[19][2]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[2] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB10_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[19]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB0_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[19][2] ));
    INV_BA AFLSDF_INV_106 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_94_net_1 ), .Y(
        AFLSDF_INV_106_net_1));
    CFG4 #( .INIT(16'hDC00) )  \CoreAPB3_0/u_mux_p_to_b3/PRDATA[10]  (
        .A(\CoreGPIO_0.N_247 ), .B(\CoreGPIO_0.N_565 ), .C(
        \CoreGPIO_0.xhdl1.GEN_BITS[10].APB_32.INTR_reg[10] ), .D(
        CoreAPB3_0_APBmslave5_PSELx), .Y(
        \FIC_MSS_0_FIC_0_APB_MASTER_PRDATA[10] ));
    CFG2 #( .INIT(4'h8) )  \FIC_MSS_0/MSS_ADLIB_INST_RNO_22  (.A(
        CoreAPB3_0_APBmslave5_PSELx), .B(
        \CoreGPIO_0.xhdl1.GEN_BITS[1].APB_32.INTR_reg[1] ), .Y(
        \FIC_MSS_0/CoreAPB3_0_APBmslave5_PRDATA_m_c_c_0[1] ));
    INV_BA AFLSDF_INV_11 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_4_net_1 ), .Y(
        AFLSDF_INV_11_net_1));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_149_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_36_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_149_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_149_rs_net_1 ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[19].REG_GEN.CONFIG_reg[19][0]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[0] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB9_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[19]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_YR ), .ADn(VCC), .SLn(
        VCC), .SD(GND), .LAT(GND), .Q(\CoreGPIO_0/CONFIG_reg[19][0] ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_151  (.A(VCC), 
        .B(VCC), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/CAN_TXBUS_F2H_SCP_net ), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/MGPIO6A_F2H_GPIN_net ), .IPC());
    CFG2 #( .INIT(4'h8) )  \CoreGPIO_0/GPOUT_reg_0_sqmuxa_0_a4_0_a2  (
        .A(\CoreGPIO_0/INTR_reg21 ), .B(
        \CoreGPIO_0.xhdl1.GEN_BITS[0].APB_32.GPOUT_reg9 ), .Y(
        \CoreGPIO_0/GPOUT_reg_0_sqmuxa ));
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_34  (
        .A(\reg_apb_wrp_0/reg16x8_0/mem_2_[4]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_501 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_34_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_5_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB4_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_8__1_sqmuxa ), .ALn(
        AFLSDF_INV_121_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_5_set_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_11_[7]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[7] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB17_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_11__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_220_i ), .ADn(VCC), .SLn(
        VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_11_rs[7] ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_89  (.A(VCC), 
        .B(VCC), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[30] ), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/RXDF_net[5] ), .IPC());
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[3].gpin1[3]  (.D(\GPIO_IN_c[3] ), 
        .CLK(\FCCC_0/GL1_INST/U0_RGB1_RGB9_rgbr_net_1 ), .EN(VCC), 
        .ALn(\MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_YR ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(GND), .Q(\CoreGPIO_0/gpin1[3] ));
    IOIN_IB \GPIO_IN_ibuf[3]/U0/U_IOIN  (.YIN(\GPIO_IN_ibuf[3]/U0/YIN )
        , .E(GND), .Y(\GPIO_IN_c[3] ));
    CFG4 #( .INIT(16'hECA0) )  \FIC_MSS_0/MSS_ADLIB_INST_RNO_13  (.A(
        \CoreAPB3_0_APBmslave3_PRDATA[3] ), .B(
        \CoreGPIO_0.RDATA_32.un12_PRDATA_o ), .C(
        CoreAPB3_0_APBmslave3_PSELx), .D(
        \FIC_MSS_0/CoreAPB3_0_APBmslave5_PRDATA_m_c_c_1[3] ), .Y(
        \FIC_MSS_0/CoreAPB3_0_APBmslave5_PRDATA_m_0_0[3] ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[15].REG_GEN.CONFIG_reg[15][5]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[5] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB10_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[15]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB0_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[15][5] ));
    CFG2 #( .INIT(4'h2) )  
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_a3_11[1]  (.A(
        \reg_apb_wrp_0/reg16x8_0/N_492 ), .B(
        \reg_apb_wrp_0/reg16x8_0/mem_9_[1]_net_1 ), .Y(
        \reg_apb_wrp_0/reg16x8_0/N_382 ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[0].APB_32.INTR_reg[0]  (.D(
        \CoreGPIO_0/INTR_reg_9[0] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB10_rgbr_net_1 ), .EN(VCC), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB0_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/INTR_reg[0] ));
    CFG3 #( .INIT(8'hF2) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_220  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_11_[7]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_505 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_220_i ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[27].REG_GEN.CONFIG_reg[27][5]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[5] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB9_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[27]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_YR ), .ADn(VCC), .SLn(
        VCC), .SD(GND), .LAT(GND), .Q(\CoreGPIO_0/CONFIG_reg[27][5] ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_53  (.A(GND), 
        .B(GND), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[7] ), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[14] ), .IPC());
    CFG3 #( .INIT(8'h20) )  
        \CoreGPIO_0/xhdl1.GEN_BITS[9].APB_32.edge_both_RNO[9]  (.A(
        \CoreGPIO_0/CONFIG_reg[9][3] ), .B(
        \CoreAPB3_0_APBmslave3_PWDATA[9] ), .C(
        \CoreGPIO_0/edge_neg[9] ), .Y(\CoreGPIO_0/edge_neg_135[9] ));
    RGB \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB5  (.An(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_YNn_GSouth ), .ENn(GND), .YL()
        , .YR(\MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB5_rgbr_net_1 ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_245  (.A(VCC), 
        .B(GND), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[57] ), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/F_WSTRB_net[5] ), .IPC());
    INV_BA AFLSDF_INV_45 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_43_net_1 ), .Y(
        AFLSDF_INV_45_net_1));
    CFG4 #( .INIT(16'hAC0F) )  
        \CoreGPIO_0/CONFIG_reg_o_2_31_bm_1_1_RNO[2]  (.A(
        \CoreGPIO_0/CONFIG_reg[13][2] ), .B(
        \CoreGPIO_0/CONFIG_reg[29][2] ), .C(
        \CoreGPIO_0/CONFIG_reg_o_2_21_1[2] ), .D(
        \CoreAPB3_0_APBmslave3_PADDR[5] ), .Y(
        \CoreGPIO_0/CONFIG_reg_o_2_31_bm_1_1_RNO[2]_net_1 ));
    INV_BA AFLSDF_INV_118 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_26_net_1 ), .Y(
        AFLSDF_INV_118_net_1));
    CFG3 #( .INIT(8'hF2) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_222  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_12_[0]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_495 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_222_i ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_136_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_10_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_136_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_136_rs_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_129_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_82_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_129_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_129_rs_net_1 ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[14].REG_GEN.CONFIG_reg[14][5]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[5] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB13_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[14]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB3_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[14][5] ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[28].REG_GEN.CONFIG_reg[28][0]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[0] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB14_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[28]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB4_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[28][0] ));
    CFG4 #( .INIT(16'hBBFB) )  \CoreGPIO_0/edge_pos_2_sqmuxa_6_i_0  (
        .A(\CoreGPIO_0/N_396 ), .B(\CoreGPIO_0/CONFIG_reg[2][3] ), .C(
        \CoreGPIO_0/INTR_reg21 ), .D(\CoreGPIO_0.N_247 ), .Y(
        \CoreGPIO_0/N_64 ));
    IOINFF_BYPASS \MSS_RESET_N_F2M_ibuf/U0/U_IOINFF  (.A(
        \MSS_RESET_N_F2M_ibuf/U0/YIN1 ), .Y(
        \MSS_RESET_N_F2M_ibuf/U0/YIN ));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_174_rs_RNIPG6V  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_15_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_174_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_5_rs[1] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_5_[1]_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_36_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB13_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_2__1_sqmuxa ), .ALn(
        AFLSDF_INV_122_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_36_set_net_1 ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_22  (.A(VCC), 
        .B(GND), .C(VCC), .IPA(), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_SIZE_net[1] ), .IPC());
    CFG4 #( .INIT(16'h4000) )  \FIC_MSS_0/MSS_ADLIB_INST_RNO_23  (.A(
        \CoreGPIO_0.N_246 ), .B(CoreAPB3_0_APBmslave5_PSELx), .C(
        \CoreGPIO_0.xhdl1.GEN_BITS[4].APB_32.GPOUT_reg[4] ), .D(
        \CoreAPB3_0_APBmslave3_PADDR[5] ), .Y(
        \FIC_MSS_0/CoreAPB3_0_APBmslave5_PRDATA_m_c_c[4] ));
    INV_BA AFLSDF_INV_70 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_42_net_1 ), .Y(
        AFLSDF_INV_70_net_1));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[23].APB_32.INTR_reg[23]  (.D(
        \CoreGPIO_0/INTR_reg_308[23] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB13_rgbr_net_1 ), .EN(VCC), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB3_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/INTR_reg[23] ));
    CFG3 #( .INIT(8'h20) )  
        \CoreGPIO_0/xhdl1.GEN_BITS[15].APB_32.edge_pos_RNO[15]  (.A(
        \CoreGPIO_0/CONFIG_reg[15][3] ), .B(
        \CoreAPB3_0_APBmslave3_PWDATA[15] ), .C(
        \CoreGPIO_0/edge_neg[15] ), .Y(\CoreGPIO_0/edge_pos_219[15] ));
    CFG4 #( .INIT(16'hA9FF) )  
        \CoreGPIO_0/xhdl1.GEN_BITS[15].APB_32.INTR_reg_204_0_o2_0_0[15]  
        (.A(\CoreGPIO_0/CONFIG_reg[15][7] ), .B(
        \CoreGPIO_0/CONFIG_reg[15][6] ), .C(
        \CoreGPIO_0/CONFIG_reg[15][5] ), .D(
        \CoreGPIO_0/CONFIG_reg[15][3] ), .Y(
        \CoreGPIO_0/INTR_reg_204_0_o2_0[15] ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_43  (.A(GND), 
        .B(GND), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[26] ), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_SEL_net ), .IPC());
    IOINFF_BYPASS \FIC_MSS_0/MDDR_DQ_15_PAD/U_IOINFF  (.A(
        \FIC_MSS_0/MDDR_DQ_15_PAD_Y ), .Y(
        \FIC_MSS_0/MDDR_DQ_15_PAD/YIN ));
    sdf_IOPAD_BI \FIC_MSS_0/MDDR_DQ_6_PAD/U_IOPAD  (.PAD(MDDR_DQ[6]), 
        .D(\FIC_MSS_0/DRAM_DQ_OUT_net_0[6] ), .E(
        \FIC_MSS_0/DRAM_DQ_OE_net_0[6] ), .Y(
        \FIC_MSS_0/MDDR_DQ_6_PAD_Y ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[12].REG_GEN.CONFIG_reg[12][4]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[4] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB14_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[12]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB4_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[12][4] ));
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_123  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_6_[7]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_493 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_123_net_1 ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[1].APB_32.edge_pos[1]  (.D(
        \CoreGPIO_0/N_107 ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB16_rgbr_net_1 ), .EN(
        \CoreGPIO_0/N_66 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB6_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/edge_pos[1] ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[16].REG_GEN.CONFIG_reg[16][2]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[2] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB15_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[16]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB5_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[16][2] ));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_8_[0]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[0] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB7_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_8__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_219_i ), .ADn(VCC), .SLn(
        VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_8_rs[0] ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[12].REG_GEN.CONFIG_reg[12][5]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[5] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB12_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[12]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB2_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[12][5] ));
    CFG4 #( .INIT(16'hA9FF) )  
        \CoreGPIO_0/xhdl1.GEN_BITS[7].APB_32.INTR_reg_100_0_o2_0_0[7]  
        (.A(\CoreGPIO_0/CONFIG_reg[7][7] ), .B(
        \CoreGPIO_0/CONFIG_reg[7][6] ), .C(
        \CoreGPIO_0/CONFIG_reg[7][5] ), .D(
        \CoreGPIO_0/CONFIG_reg[7][3] ), .Y(
        \CoreGPIO_0/INTR_reg_100_0_o2_0[7] ));
    CFG4 #( .INIT(16'h330A) )  
        \CoreGPIO_0/xhdl1.GEN_BITS[15].APB_32.INTR_reg_204_0[15]  (.A(
        \CoreGPIO_0/INTR_reg[15] ), .B(
        \CoreGPIO_0/INTR_reg_204_0_o2_1[15] ), .C(
        \CoreAPB3_0_APBmslave3_PWDATA[15] ), .D(\CoreGPIO_0/N_248 ), 
        .Y(\CoreGPIO_0/INTR_reg_204[15] ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[4].gpin1[4]  (.D(\GPIO_IN_c[4] ), 
        .CLK(\FCCC_0/GL1_INST/U0_RGB1_RGB12_rgbr_net_1 ), .EN(VCC), 
        .ALn(\MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB2_rgbr_net_1 ), 
        .ADn(VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/gpin1[4] ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_222  (.A(VCC), 
        .B(VCC), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[6] ), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/F_WDATA_HWDATA01_net[18] ), .IPC());
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_142  (.A(VCC), 
        .B(VCC), .C(VCC), .IPA(), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/SPI1_CLK_IN_net ), .IPC());
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_60  (.A(GND), 
        .B(VCC), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[21] ), .IPB(), .IPC()
        );
    CFG2 #( .INIT(4'h7) )  \CoreGPIO_0/edge_both_2_sqmuxa_27_i  (.A(
        \CoreGPIO_0/N_248 ), .B(\CoreGPIO_0/CONFIG_reg[28][3] ), .Y(
        \CoreGPIO_0/N_163 ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_215  (.A(GND), 
        .B(GND), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/F_AWSIZE_HSIZE0_net[1] ), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/F_WID_HREADY01_net[3] ), .IPC());
    IOOUTFF_BYPASS \GPIO_OUT_obuf[4]/U0/U_IOOUTFF  (.A(
        \GPIO_OUT_obuf[4]/U0/DOUT1 ), .Y(\GPIO_OUT_obuf[4]/U0/DOUT ));
    CFG2 #( .INIT(4'h4) )  \CoreGPIO_0/PRDATA_0_iv_0_a2_0[25]  (.A(
        \CoreGPIO_0.N_247 ), .B(\CoreGPIO_0/INTR_reg[25] ), .Y(
        \CoreGPIO_0.N_536 ));
    CFG4 #( .INIT(16'h0F35) )  
        \CoreGPIO_0/CONFIG_reg_o_2_31_am_1_RNO_1[7]  (.A(
        \CoreGPIO_0/CONFIG_reg[4][7] ), .B(
        \CoreGPIO_0/CONFIG_reg[20][7] ), .C(
        \CoreAPB3_0_APBmslave3_PADDR[6] ), .D(
        \CoreAPB3_0_APBmslave3_PADDR[5] ), .Y(
        \CoreGPIO_0/CONFIG_reg_o_2_6_1[7] ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[8].REG_GEN.CONFIG_reg[8][5]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[5] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB9_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[8]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_YR ), .ADn(VCC), .SLn(
        VCC), .SD(GND), .LAT(GND), .Q(\CoreGPIO_0/CONFIG_reg[8][5] ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[17].REG_GEN.CONFIG_reg[17][4]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[4] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB14_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[17]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB4_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[17][4] ));
    INV_BA AFLSDF_INV_104 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_107_net_1 ), .Y(
        AFLSDF_INV_104_net_1));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_251_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_61_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_251_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_251_rs_net_1 ));
    CFG4 #( .INIT(16'hA9FF) )  
        \CoreGPIO_0/xhdl1.GEN_BITS[23].APB_32.INTR_reg_308_0_o2_0_0[23]  
        (.A(\CoreGPIO_0/CONFIG_reg[23][7] ), .B(
        \CoreGPIO_0/CONFIG_reg[23][6] ), .C(
        \CoreGPIO_0/CONFIG_reg[23][5] ), .D(
        \CoreGPIO_0/CONFIG_reg[23][3] ), .Y(
        \CoreGPIO_0/INTR_reg_308_0_o2_0[23] ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[25].APB_32.INTR_reg[25]  (.D(
        \CoreGPIO_0/INTR_reg_334[25] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB14_rgbr_net_1 ), .EN(VCC), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB4_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/INTR_reg[25] ));
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_121  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_6_[6]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_493 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_121_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_185_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_77_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_185_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_185_rs_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_118_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB13_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_14__1_sqmuxa ), .ALn(
        AFLSDF_INV_123_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_118_set_net_1 ));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_25_set_RNI0VMT  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_25_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_184_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_5_rs[6] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_5_[6]_net_1 ));
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_53  (
        .A(\reg_apb_wrp_0/reg16x8_0/mem_7_[4]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_498 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_53_net_1 ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[13].REG_GEN.CONFIG_reg[13][5]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[5] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB13_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[13]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB3_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[13][5] ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_127  (.A(GND), 
        .B(GND), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[2] ), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/F2H_INTERRUPT_net[9] ), .IPC());
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[11].APB_32.GPOUT_reg[11]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[11] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB13_rgbr_net_1 ), .EN(
        \CoreGPIO_0/GPOUT_reg_0_sqmuxa ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB3_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0.xhdl1.GEN_BITS[11].APB_32.GPOUT_reg[11] ));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_11_[6]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[6] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB16_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_11__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_218_i ), .ADn(VCC), .SLn(
        VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_11_rs[6] ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[22].REG_GEN.CONFIG_reg[22][7]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[7] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB12_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[22]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB2_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[22][7] ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[10].REG_GEN.CONFIG_reg[10][7]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[7] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB17_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[10]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB7_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[10][7] ));
    IOINFF_BYPASS \FIC_MSS_0/MDDR_DQ_2_PAD/U_IOINFF  (.A(
        \FIC_MSS_0/MDDR_DQ_2_PAD_Y ), .Y(\FIC_MSS_0/MDDR_DQ_2_PAD/YIN )
        );
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_102  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_10_[5]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_491 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_102_net_1 ));
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_32  (
        .A(\reg_apb_wrp_0/reg16x8_0/mem_2_[3]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_501 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_32_net_1 ));
    IOBI_IB_OB_EB \FIC_MSS_0/MDDR_DQ_2_PAD/U_IOBI  (.D(VCC), .E(VCC), 
        .YIN(\FIC_MSS_0/MDDR_DQ_2_PAD/YIN ), .DOUT(), .EOUT(), .Y());
    IOINFF_BYPASS \FIC_MSS_0/MDDR_DQS_TMATCH_0_IN_PAD/U_IOINFF  (.A(
        \FIC_MSS_0/MDDR_DQS_TMATCH_0_IN_PAD_Y ), .Y(
        \FIC_MSS_0/MDDR_DQS_TMATCH_0_IN_PAD/YIN ));
    RGB \FCCC_0/GL1_INST/U0_RGB1  (.An(\FCCC_0/GL1_INST/U0_YNn ), .ENn(
        GND), .YL(), .YR(\FCCC_0/GL1_INST/U0_RGB1_YR ));
    CFG4 #( .INIT(16'h330A) )  
        \CoreGPIO_0/xhdl1.GEN_BITS[16].APB_32.INTR_reg_217_0[16]  (.A(
        \CoreGPIO_0/INTR_reg[16] ), .B(
        \CoreGPIO_0/INTR_reg_217_0_o2_1[16] ), .C(
        \CoreAPB3_0_APBmslave3_PWDATA[16] ), .D(\CoreGPIO_0/N_248 ), 
        .Y(\CoreGPIO_0/INTR_reg_217[16] ));
    sdf_IOPAD_BI \FIC_MSS_0/MDDR_DQ_3_PAD/U_IOPAD  (.PAD(MDDR_DQ[3]), 
        .D(\FIC_MSS_0/DRAM_DQ_OUT_net_0[3] ), .E(
        \FIC_MSS_0/DRAM_DQ_OE_net_0[3] ), .Y(
        \FIC_MSS_0/MDDR_DQ_3_PAD_Y ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_196_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_37_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_196_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_196_rs_net_1 ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[31].REG_GEN.CONFIG_reg[31][2]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[2] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB11_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[31]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB1_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[31][2] ));
    CFG4 #( .INIT(16'h0F35) )  
        \CoreGPIO_0/CONFIG_reg_o_2_31_am_1_RNO_1[2]  (.A(
        \CoreGPIO_0/CONFIG_reg[4][2] ), .B(
        \CoreGPIO_0/CONFIG_reg[20][2] ), .C(
        \CoreAPB3_0_APBmslave3_PADDR[6] ), .D(
        \CoreAPB3_0_APBmslave3_PADDR[5] ), .Y(
        \CoreGPIO_0/CONFIG_reg_o_2_6_1[2] ));
    CFG4 #( .INIT(16'hAC0F) )  
        \CoreGPIO_0/CONFIG_reg_o_2_31_am_1_RNO_0[7]  (.A(
        \CoreGPIO_0/CONFIG_reg[8][7] ), .B(
        \CoreGPIO_0/CONFIG_reg[24][7] ), .C(
        \CoreGPIO_0/CONFIG_reg_o_2_3_1[7] ), .D(
        \CoreAPB3_0_APBmslave3_PADDR[5] ), .Y(
        \CoreGPIO_0/CONFIG_reg_o_2_31_am_1_RNO_0[7]_net_1 ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_112  (.A(VCC), 
        .B(VCC), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/FAB_XDATAIN_net[4] ), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/FAB_VSTATUS_net[1] ), .IPC());
    CFG4 #( .INIT(16'hAC0F) )  
        \CoreGPIO_0/CONFIG_reg_o_2_31_am_RNO_0[1]  (.A(
        \CoreGPIO_0/CONFIG_reg[14][1] ), .B(
        \CoreGPIO_0/CONFIG_reg[30][1] ), .C(
        \CoreGPIO_0/CONFIG_reg_o_2_13_1_1[1] ), .D(
        \CoreAPB3_0_APBmslave3_PADDR[5] ), .Y(
        \CoreGPIO_0/CONFIG_reg_o_2_31_am_RNO_0[1]_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_0_[3]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[3] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB9_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_0__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_130_i ), .ADn(VCC), .SLn(
        VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_0_rs[3] ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[5].APB_32.GPOUT_reg[5]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[5] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB11_rgbr_net_1 ), .EN(
        \CoreGPIO_0/GPOUT_reg_0_sqmuxa ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB1_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0.xhdl1.GEN_BITS[5].APB_32.GPOUT_reg[5] ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[31].REG_GEN.CONFIG_reg[31][0]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[0] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB11_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[31]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB1_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[31][0] ));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_186_rs_RNI5E981  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_27_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_186_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_5_rs[7] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_5_[7]_net_1 ));
    CFG4 #( .INIT(16'hEC00) )  \CoreAPB3_0/u_mux_p_to_b3/PRDATA[12]  (
        .A(\CoreGPIO_0.xhdl1.GEN_BITS[0].APB_32.GPOUT_reg9 ), .B(
        \CoreGPIO_0.N_562 ), .C(
        \CoreGPIO_0.xhdl1.GEN_BITS[12].APB_32.GPOUT_reg[12] ), .D(
        CoreAPB3_0_APBmslave5_PSELx), .Y(
        \FIC_MSS_0_FIC_0_APB_MASTER_PRDATA[12] ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_134_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_87_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_134_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_134_rs_net_1 ));
    CFG4 #( .INIT(16'hAC0F) )  
        \CoreGPIO_0/CONFIG_reg_o_2_31_am_1_1_RNO[7]  (.A(
        \CoreGPIO_0/CONFIG_reg[12][7] ), .B(
        \CoreGPIO_0/CONFIG_reg[28][7] ), .C(
        \CoreGPIO_0/CONFIG_reg_o_2_6_1[7] ), .D(
        \CoreAPB3_0_APBmslave3_PADDR[5] ), .Y(
        \CoreGPIO_0/CONFIG_reg_o_2_31_am_1_1_RNO[7]_net_1 ));
    CFG2 #( .INIT(4'h8) )  \CoreGPIO_0/PRDATA_0_iv_0_0_a2_0_0[7]  (.A(
        \CoreAPB3_0_APBmslave3_PADDR[5] ), .B(
        \CoreGPIO_0/GPOUT_reg[7] ), .Y(
        \CoreGPIO_0/PRDATA_0_iv_0_0_a2_0_0[7]_net_1 ));
    INV_BA AFLSDF_INV_98 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_37_net_1 ), .Y(
        AFLSDF_INV_98_net_1));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_58_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB6_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_15__1_sqmuxa ), .ALn(
        AFLSDF_INV_124_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_58_set_net_1 ));
    CFG4 #( .INIT(16'h4000) )  
        \CoreGPIO_0/xhdl1.GEN_BITS[21].REG_GEN.CONFIG_reg[21]2_0_a4_0_a2  
        (.A(\CoreAPB3_0_APBmslave3_PADDR[3] ), .B(
        \CoreAPB3_0_APBmslave3_PADDR[2] ), .C(\CoreGPIO_0/N_598 ), .D(
        \CoreGPIO_0/N_603 ), .Y(\CoreGPIO_0/CONFIG_reg[21]2 ));
    CFG2 #( .INIT(4'h6) )  \CoreGPIO_0/edge_both_2_sqmuxa_14_i_x2  (.A(
        \CoreGPIO_0/gpin2[1] ), .B(
        \CoreGPIO_0.xhdl1.GEN_BITS[1].gpin3[1] ), .Y(
        \CoreGPIO_0/N_142_i ));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_243_rs_RNIP2DD  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_115_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_243_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_14_rs[3] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_14_[3]_net_1 ));
    CFG4 #( .INIT(16'hAC0F) )  
        \CoreGPIO_0/CONFIG_reg_o_2_31_bm_1_RNO_0[3]  (.A(
        \CoreGPIO_0/CONFIG_reg[9][3] ), .B(
        \CoreGPIO_0/CONFIG_reg[25][3] ), .C(
        \CoreGPIO_0/CONFIG_reg_o_2_18_1[3] ), .D(
        \CoreAPB3_0_APBmslave3_PADDR[5] ), .Y(
        \CoreGPIO_0/CONFIG_reg_o_2_31_bm_1_RNO_0[3]_net_1 ));
    INV_BA AFLSDF_INV_100 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_20_net_1 ), .Y(
        AFLSDF_INV_100_net_1));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[26].REG_GEN.CONFIG_reg[26][6]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[6] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB17_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[26]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB7_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[26][6] ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[2].REG_GEN.CONFIG_reg[2][3]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[3] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB17_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[2]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB7_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[2][3] ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_139  (.A(VCC), 
        .B(VCC), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/SMBSUS_NI1_net ), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/F2_DMAREADY_net[1] ), .IPC());
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_135  (.A(VCC), 
        .B(MSS_RESET_N_F2M_ibuf), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/SMBALERT_NI0_net ), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/USER_MSS_RESET_N_net ), .IPC());
    CFG2 #( .INIT(4'h2) )  
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_a3_3[2]  (.A(
        \reg_apb_wrp_0/reg16x8_0/N_500 ), .B(
        \reg_apb_wrp_0/reg16x8_0/mem_13_[2]_net_1 ), .Y(
        \reg_apb_wrp_0/reg16x8_0/N_390 ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_22_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB1_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_12__1_sqmuxa ), .ALn(
        AFLSDF_INV_125_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_22_set_net_1 ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_280  (.A(VCC), 
        .B(VCC), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PADDR_net[3] ), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[7] ), .IPC());
    INV_BA AFLSDF_INV_102 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_23_net_1 ), .Y(
        AFLSDF_INV_102_net_1));
    CFG3 #( .INIT(8'hF2) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_217  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_7_[7]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_498 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_217_i ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[24].REG_GEN.CONFIG_reg[24][5]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[5] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB11_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[24]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB1_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[24][5] ));
    CFG4 #( .INIT(16'hAC0F) )  
        \CoreGPIO_0/CONFIG_reg_o_2_31_am_1_RNO_0[6]  (.A(
        \CoreGPIO_0/CONFIG_reg[8][6] ), .B(
        \CoreGPIO_0/CONFIG_reg[24][6] ), .C(
        \CoreGPIO_0/CONFIG_reg_o_2_3_1[6] ), .D(
        \CoreAPB3_0_APBmslave3_PADDR[5] ), .Y(
        \CoreGPIO_0/CONFIG_reg_o_2_31_am_1_RNO_0[6]_net_1 ));
    RGB \FCCC_0/GL1_INST/U0_RGB1_RGB2  (.An(\FCCC_0/GL1_INST/U0_YNn ), 
        .ENn(GND), .YL(\FCCC_0/GL1_INST/U0_RGB1_RGB2_rgbl_net_1 ), .YR(
        \FCCC_0/GL1_INST/U0_RGB1_RGB2_rgbr_net_1 ));
    CFG3 #( .INIT(8'hF2) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_211  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_11_[2]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_505 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_211_i ));
    CFG4 #( .INIT(16'h7350) )  
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_0_0[5]  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_13_[5]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/mem_5_[5]_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/N_500 ), .D(
        \reg_apb_wrp_0/reg16x8_0/N_490 ), .Y(
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_0_0[5]_net_1 ));
    CFG2 #( .INIT(4'h4) )  \CoreGPIO_0/edge_neg_2_sqmuxa_11_i_a2  (.A(
        \CoreGPIO_0/gpin2[1] ), .B(
        \CoreGPIO_0.xhdl1.GEN_BITS[1].gpin3[1] ), .Y(
        \CoreGPIO_0/N_399 ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[6].REG_GEN.CONFIG_reg[6][0]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[0] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB14_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[6]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB4_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[6][0] ));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_132_rs_RNIOCGF  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_85_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_132_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_0_rs[4] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_0_[4]_net_1 ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[20].REG_GEN.CONFIG_reg[20][7]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[7] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB12_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[20]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB2_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[20][7] ));
    IOENFF_BYPASS \GPIO_OUT_obuf[1]/U0/U_IOENFF  (.A(
        \GPIO_OUT_obuf[1]/U0/EOUT1 ), .Y(\GPIO_OUT_obuf[1]/U0/EOUT ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_287  (.A(VCC), 
        .B(VCC), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PADDR_net[10] ), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/MDDR_FABRIC_PWDATA_net[14] ), .IPC());
    INV_BA AFLSDF_INV_7 (.A(\FCCC_0/GL1_net ), .Y(AFLSDF_INV_7_net_1));
    IOINFF_BYPASS \GPIO_IN_ibuf[4]/U0/U_IOINFF  (.A(
        \GPIO_IN_ibuf[4]/U0/YIN1 ), .Y(\GPIO_IN_ibuf[4]/U0/YIN ));
    CFG4 #( .INIT(16'hEFEE) )  
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_9[3]  (.A(
        \reg_apb_wrp_0/reg16x8_0/N_414 ), .B(
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_3[3]_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_1_[3]_net_1 ), .D(
        \reg_apb_wrp_0/reg16x8_0/N_502 ), .Y(
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_9[3]_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_12_[1]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[1] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB4_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_12__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_224_i ), .ADn(VCC), .SLn(
        VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_12_rs[1] ));
    IOINFF_BYPASS \FIC_MSS_0/MDDR_DQ_6_PAD/U_IOINFF  (.A(
        \FIC_MSS_0/MDDR_DQ_6_PAD_Y ), .Y(\FIC_MSS_0/MDDR_DQ_6_PAD/YIN )
        );
    INV_BA AFLSDF_INV_41 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_112_net_1 ), .Y(
        AFLSDF_INV_41_net_1));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[25].REG_GEN.CONFIG_reg[25][1]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[1] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB16_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[25]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB6_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[25][1] ));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_106_set_RNINRVV  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_106_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_234_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_13_rs[2] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_13_[2]_net_1 ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[23].APB_32.GPOUT_reg[23]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[23] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB13_rgbr_net_1 ), .EN(
        \CoreGPIO_0/GPOUT_reg_0_sqmuxa ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB3_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0.xhdl1.GEN_BITS[23].APB_32.GPOUT_reg[23] ));
    CFG4 #( .INIT(16'h0001) )  
        \reg_apb_wrp_0/reg16x8_0/temp_data_RNO[0]  (.A(
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_11[0]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_10[0]_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_9[0]_net_1 ), .D(
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_8[0]_net_1 ), .Y(
        \reg_apb_wrp_0/reg16x8_0/N_5_i_0 ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[5].REG_GEN.CONFIG_reg[5][0]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[0] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB14_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[5]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB4_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[5][0] ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_13  (.A(
        \FIC_MSS_0_FIC_0_APB_MASTER_PRDATA[18] ), .B(VCC), .C(VCC), 
        .IPA(\FIC_MSS_0/MSS_ADLIB_INST/F_HM0_RDATA_net[18] ), .IPB(), 
        .IPC());
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[1].REG_GEN.CONFIG_reg[1][5]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[5] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB15_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[1]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB5_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[1][5] ));
    CFG3 #( .INIT(8'hF2) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_233  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_13_[1]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_500 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_233_i ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[21].REG_GEN.CONFIG_reg[21][0]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[0] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB14_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[21]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB4_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[21][0] ));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_12_[7]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[7] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB6_rgbr_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_12__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_231_i ), .ADn(VCC), .SLn(
        VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_12_rs[7] ));
    IOTRI_OB_EB \FIC_MSS_0/MMUART_0_TXD_PAD/U_IOOUT  (.D(VCC), .E(VCC), 
        .DOUT(), .EOUT());
    RGB \FCCC_0/GL1_INST/U0_RGB1_RGB12  (.An(
        \FCCC_0/GL1_INST/U0_YNn_GSouth ), .ENn(GND), .YL(
        \FCCC_0/GL1_INST/U0_RGB1_RGB12_rgbl_net_1 ), .YR(
        \FCCC_0/GL1_INST/U0_RGB1_RGB12_rgbr_net_1 ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[13].REG_GEN.CONFIG_reg[13][7]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[7] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB13_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[13]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB3_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[13][7] ));
    sdf_IOPAD_TRI \GPIO_OUT_obuf[3]/U0/U_IOPAD  (.PAD(GPIO_OUT[3]), .D(
        \GPIO_OUT_obuf[3]/U0/DOUT ), .E(\GPIO_OUT_obuf[3]/U0/EOUT ));
    sdf_IOPAD_TRI \FIC_MSS_0/MDDR_ADDR_5_PAD/U_IOPAD  (.PAD(
        MDDR_ADDR[5]), .D(\FIC_MSS_0/DRAM_ADDR_net_0[5] ), .E(
        \FIC_MSS_0/MDDR_ADDR_5_PAD/EOUT ));
    IOTRI_OB_EB \GPIO_OUT_obuf[3]/U0/U_IOTRI  (.D(\GPIO_OUT_net_2[3] ), 
        .E(VCC), .DOUT(\GPIO_OUT_obuf[3]/U0/DOUT1 ), .EOUT(
        \GPIO_OUT_obuf[3]/U0/EOUT1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_194_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_35_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_194_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_194_rs_net_1 ));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/mem_15__RNIIISL[6]  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_63_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_255_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_15_rs[6] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_15_[6]_net_1 ));
    CFG4 #( .INIT(16'h0400) )  
        \CoreGPIO_0/xhdl1.GEN_BITS[0].REG_GEN.CONFIG_reg[0]2_0_a4_0_a2  
        (.A(\CoreAPB3_0_APBmslave3_PADDR[7] ), .B(\CoreGPIO_0/N_606 ), 
        .C(\CoreGPIO_0/N_243 ), .D(\CoreGPIO_0/INTR_reg21 ), .Y(
        \CoreGPIO_0/CONFIG_reg[0]2 ));
    CFG4 #( .INIT(16'hB383) )  \CoreGPIO_0/CONFIG_reg_o_2_31_am[2]  (
        .A(\CoreGPIO_0/CONFIG_reg_o_2_31_am_RNO[2]_net_1 ), .B(
        \CoreGPIO_0/CONFIG_reg_o_2_31_am_1[2] ), .C(
        \CoreAPB3_0_APBmslave3_PADDR[3] ), .D(
        \CoreGPIO_0/CONFIG_reg_o_2_31_am_RNO_0[2]_net_1 ), .Y(
        \CoreGPIO_0/CONFIG_reg_o_2_31_am[2]_net_1 ));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_16_set_RNI1UDI  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_16_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_222_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_12_rs[0] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_12_[0]_net_1 ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_39  (.A(GND), 
        .B(GND), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[22] ), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[29] ), .IPC());
    IOIN_IB \GPIO_IN_ibuf[4]/U0/U_IOIN  (.YIN(\GPIO_IN_ibuf[4]/U0/YIN )
        , .E(GND), .Y(\GPIO_IN_c[4] ));
    RGB \FCCC_0/GL1_INST/U0_RGB1_RGB11  (.An(
        \FCCC_0/GL1_INST/U0_YNn_GSouth ), .ENn(GND), .YL(
        \FCCC_0/GL1_INST/U0_RGB1_RGB11_rgbl_net_1 ), .YR(
        \FCCC_0/GL1_INST/U0_RGB1_RGB11_rgbr_net_1 ));
    INV_BA AFLSDF_INV_55 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_115_net_1 ), .Y(
        AFLSDF_INV_55_net_1));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_15_[0]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[0] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB6_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_15__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_248_i ), .ADn(VCC), .SLn(
        VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_15_rs[0] ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_81_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB4_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_0__1_sqmuxa ), .ALn(
        AFLSDF_INV_126_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_81_set_net_1 ));
    CFG4 #( .INIT(16'h1000) )  
        \CoreGPIO_0/xhdl1.GEN_BITS[16].REG_GEN.CONFIG_reg[16]2_0_a4_0_a2  
        (.A(\CoreAPB3_0_APBmslave3_PADDR[3] ), .B(
        \CoreAPB3_0_APBmslave3_PADDR[2] ), .C(\CoreGPIO_0/N_598 ), .D(
        \CoreGPIO_0/N_606 ), .Y(\CoreGPIO_0/CONFIG_reg[16]2 ));
    CFG4 #( .INIT(16'hAC0F) )  
        \CoreGPIO_0/CONFIG_reg_o_2_31_bm_RNO_0[0]  (.A(
        \CoreGPIO_0/CONFIG_reg[15][0] ), .B(
        \CoreGPIO_0/CONFIG_reg[31][0] ), .C(
        \CoreGPIO_0/CONFIG_reg_o_2_28_1_1[0] ), .D(
        \CoreAPB3_0_APBmslave3_PADDR[5] ), .Y(
        \CoreGPIO_0/CONFIG_reg_o_2_31_bm_RNO_0[0]_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_145_rs  (.D(VCC), .CLK(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_28_net_1 ), .EN(VCC), 
        .ALn(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_145_i ), .ADn(VCC), 
        .SLn(VCC), .SD(GND), .LAT(VCC), .Q(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_145_rs_net_1 ));
    CFG4 #( .INIT(16'hF2F3) )  
        \CoreGPIO_0/xhdl1.GEN_BITS[15].APB_32.INTR_reg_204_0_o2_1_0[15]  
        (.A(\CoreGPIO_0/CONFIG_reg[15][6] ), .B(
        \CoreGPIO_0/edge_neg[15] ), .C(
        \CoreGPIO_0/INTR_reg_204_0_o2_0[15] ), .D(
        \CoreGPIO_0/CONFIG_reg[15][5] ), .Y(
        \CoreGPIO_0/INTR_reg_204_0_o2_1[15] ));
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_14  (
        .A(\reg_apb_wrp_0/reg16x8_0/mem_1_[2]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_502 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_14_net_1 ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_50  (.A(GND), 
        .B(VCC), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_WDATA_net[4] ), .IPB(), .IPC());
    RGB \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB0  (.An(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_YNn_GSouth ), .ENn(GND), .YL()
        , .YR(\MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB0_rgbr_net_1 ));
    CFG4 #( .INIT(16'h7530) )  
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_4[4]  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_12_[4]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/mem_4_[4]_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/N_504 ), .D(
        \reg_apb_wrp_0/reg16x8_0/N_495 ), .Y(
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_4[4]_net_1 ));
    CFG4 #( .INIT(16'h0F35) )  
        \CoreGPIO_0/CONFIG_reg_o_2_31_bm_RNO_2[6]  (.A(
        \CoreGPIO_0/CONFIG_reg[7][6] ), .B(
        \CoreGPIO_0/CONFIG_reg[23][6] ), .C(
        \CoreAPB3_0_APBmslave3_PADDR[6] ), .D(
        \CoreAPB3_0_APBmslave3_PADDR[5] ), .Y(
        \CoreGPIO_0/CONFIG_reg_o_2_28_1_1[6] ));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_203_rs_RNIHO59  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_103_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_203_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_10_rs[6] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_10_[6]_net_1 ));
    CFG4 #( .INIT(16'h7350) )  
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_6[4]  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_8_[4]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/mem_0_[4]_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/N_499 ), .D(
        \reg_apb_wrp_0/reg16x8_0/N_496 ), .Y(
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_6[4]_net_1 ));
    CFG2 #( .INIT(4'h8) )  
        \reg_apb_wrp_0/reg16x8_0/mem_2__1_sqmuxa_0_a3  (.A(
        \reg_apb_wrp_0/reg16x8_0/N_501 ), .B(
        \reg_apb_wrp_0/wr_enable_net_1 ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_2__1_sqmuxa ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_166  (.A(VCC), 
        .B(VCC), .C(VCC), .IPA(), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/MGPIO11B_F2H_GPIN_net ), .IPC());
    CFG4 #( .INIT(16'h0F35) )  
        \CoreGPIO_0/CONFIG_reg_o_2_31_bm_RNO_2[7]  (.A(
        \CoreGPIO_0/CONFIG_reg[7][7] ), .B(
        \CoreGPIO_0/CONFIG_reg[23][7] ), .C(
        \CoreAPB3_0_APBmslave3_PADDR[6] ), .D(
        \CoreAPB3_0_APBmslave3_PADDR[5] ), .Y(
        \CoreGPIO_0/CONFIG_reg_o_2_28_1_1[7] ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[21].REG_GEN.CONFIG_reg[21][2]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[2] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB14_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[21]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB4_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[21][2] ));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_6_[5]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[5] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB11_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_6__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_198_i ), .ADn(VCC), .SLn(
        VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_6_rs[5] ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_76  (.A(VCC), 
        .B(VCC), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[10] ), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/PER2_FABRIC_PRDATA_net[17] ), .IPC());
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_68_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB18_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_8__1_sqmuxa ), .ALn(
        AFLSDF_INV_127_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_68_set_net_1 ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_40  (.A(GND), 
        .B(GND), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[23] ), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/F_FM0_ADDR_net[30] ), .IPC());
    CFG4 #( .INIT(16'hDC00) )  \CoreAPB3_0/u_mux_p_to_b3/PRDATA[26]  (
        .A(\CoreGPIO_0.N_247 ), .B(\CoreGPIO_0.N_533 ), .C(
        \CoreGPIO_0.xhdl1.GEN_BITS[26].APB_32.INTR_reg[26] ), .D(
        CoreAPB3_0_APBmslave5_PSELx), .Y(
        \FIC_MSS_0_FIC_0_APB_MASTER_PRDATA[26] ));
    CFG4 #( .INIT(16'hC480) )  
        \CoreGPIO_0/xhdl1.GEN_BITS[0].APB_32.INTR_reg_9_0_0_RNO[0]  (
        .A(\CoreGPIO_0/CONFIG_reg[0][7] ), .B(
        \CoreGPIO_0/CONFIG_reg[0][3] ), .C(
        \CoreGPIO_0/INTR_reg_9_0_0_50_tz_1 ), .D(
        \CoreGPIO_0/INTR_reg_9_0_0_m2[0] ), .Y(\CoreGPIO_0/N_1575_tz ));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_239_rs_RNIT0RQ  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_111_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_239_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_13_rs[7] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_13_[7]_net_1 ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[24].REG_GEN.CONFIG_reg[24][1]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[1] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB15_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[24]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB5_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[24][1] ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_24_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB16_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_1__1_sqmuxa ), .ALn(
        AFLSDF_INV_128_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_24_set_net_1 ));
    CFG4 #( .INIT(16'h7350) )  
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_0_3[5]  (.A(
        \reg_apb_wrp_0/reg16x8_0/mem_11_[5]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/mem_3_[5]_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/N_505 ), .D(
        \reg_apb_wrp_0/reg16x8_0/N_494 ), .Y(
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_0_3[5]_net_1 ));
    IP_INTERFACE \FCCC_0/CCC_INST/IP_INTERFACE_16  (.A(VCC), .B(VCC), 
        .C(VCC), .IPA(), .IPB(\FCCC_0/CCC_INST/GPD2_ARST_N_net ), .IPC(
        \FCCC_0/CCC_INST/PADDR_net[6] ));
    CFG4 #( .INIT(16'hEC00) )  \CoreAPB3_0/u_mux_p_to_b3/PRDATA[9]  (
        .A(\CoreGPIO_0.xhdl1.GEN_BITS[0].APB_32.GPOUT_reg9 ), .B(
        \CoreGPIO_0.N_568 ), .C(
        \CoreGPIO_0.xhdl1.GEN_BITS[9].APB_32.GPOUT_reg[9] ), .D(
        CoreAPB3_0_APBmslave5_PSELx), .Y(
        \FIC_MSS_0_FIC_0_APB_MASTER_PRDATA[9] ));
    sdf_IOPAD_IN \GPIO_IN_ibuf[0]/U0/U_IOPAD  (.PAD(GPIO_IN[0]), .Y(
        \GPIO_IN_ibuf[0]/U0/YIN1 ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[22].REG_GEN.CONFIG_reg[22][6]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[6] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB12_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[22]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB2_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[22][6] ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[2].REG_GEN.CONFIG_reg[2][6]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[6] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB17_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[2]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB7_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[2][6] ));
    SLE \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_32_set  (.D(
        CFG0_GND_INST_NET), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB8_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_2__1_sqmuxa ), .ALn(
        AFLSDF_INV_129_net_1), .ADn(GND), .SLn(VCC), .SD(GND), .LAT(
        GND), .Q(\reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_32_set_net_1 ));
    SLE \reg_apb_wrp_0/reg16x8_0/mem_12_[6]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[6] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB4_rgbl_net_1 ), .EN(
        \reg_apb_wrp_0/reg16x8_0/mem_12__1_sqmuxa ), .ALn(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_230_i ), .ADn(VCC), .SLn(
        VCC), .SD(GND), .LAT(GND), .Q(
        \reg_apb_wrp_0/reg16x8_0/mem_12_rs[6] ));
    INV_BA AFLSDF_INV_22 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_120_net_1 ), .Y(
        AFLSDF_INV_22_net_1));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_261  (.A(VCC), 
        .B(VCC), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[9] ), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[21] ), .IPC());
    CFG4 #( .INIT(16'hAC0F) )  
        \CoreGPIO_0/CONFIG_reg_o_2_31_bm_1_RNO_0[4]  (.A(
        \CoreGPIO_0/CONFIG_reg[9][4] ), .B(
        \CoreGPIO_0/CONFIG_reg[25][4] ), .C(
        \CoreGPIO_0/CONFIG_reg_o_2_18_1[4] ), .D(
        \CoreAPB3_0_APBmslave3_PADDR[5] ), .Y(
        \CoreGPIO_0/CONFIG_reg_o_2_31_bm_1_RNO_0[4]_net_1 ));
    INV_BA AFLSDF_INV_82 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_53_net_1 ), .Y(
        AFLSDF_INV_82_net_1));
    INV_BA AFLSDF_INV_109 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_52_net_1 ), .Y(
        AFLSDF_INV_109_net_1));
    CFG4 #( .INIT(16'hEC00) )  \CoreAPB3_0/u_mux_p_to_b3/PRDATA[17]  (
        .A(\CoreGPIO_0.xhdl1.GEN_BITS[0].APB_32.GPOUT_reg9 ), .B(
        \CoreGPIO_0.N_552 ), .C(
        \CoreGPIO_0.xhdl1.GEN_BITS[17].APB_32.GPOUT_reg[17] ), .D(
        CoreAPB3_0_APBmslave5_PSELx), .Y(
        \FIC_MSS_0_FIC_0_APB_MASTER_PRDATA[17] ));
    CFG4 #( .INIT(16'h330A) )  
        \CoreGPIO_0/xhdl1.GEN_BITS[23].APB_32.INTR_reg_308_0[23]  (.A(
        \CoreGPIO_0/INTR_reg[23] ), .B(
        \CoreGPIO_0/INTR_reg_308_0_o2_1[23] ), .C(
        \CoreAPB3_0_APBmslave3_PWDATA[23] ), .D(\CoreGPIO_0/N_248 ), 
        .Y(\CoreGPIO_0/INTR_reg_308[23] ));
    IP_INTERFACE \FCCC_0/CCC_INST/IP_INTERFACE_4  (.A(VCC), .B(VCC), 
        .C(VCC), .IPA(), .IPB(\FCCC_0/CCC_INST/NGMUX0_HOLD_N_net ), 
        .IPC(\FCCC_0/CCC_INST/PWDATA_net[2] ));
    CFG4 #( .INIT(16'h0F35) )  
        \CoreGPIO_0/CONFIG_reg_o_2_31_bm_RNO_1[7]  (.A(
        \CoreGPIO_0/CONFIG_reg[3][7] ), .B(
        \CoreGPIO_0/CONFIG_reg[19][7] ), .C(
        \CoreAPB3_0_APBmslave3_PADDR[6] ), .D(
        \CoreAPB3_0_APBmslave3_PADDR[5] ), .Y(
        \CoreGPIO_0/CONFIG_reg_o_2_25_1_1[7] ));
    SLE \CoreGPIO_0/xhdl1.GEN_BITS[17].REG_GEN.CONFIG_reg[17][5]  (.D(
        \CoreAPB3_0_APBmslave3_PWDATA[5] ), .CLK(
        \FCCC_0/GL1_INST/U0_RGB1_RGB15_rgbr_net_1 ), .EN(
        \CoreGPIO_0/CONFIG_reg[17]2 ), .ALn(
        \MSS_RESET_N_F2M_ibuf_RNIBBDD/U0_RGB1_RGB5_rgbr_net_1 ), .ADn(
        VCC), .SLn(VCC), .SD(GND), .LAT(GND), .Q(
        \CoreGPIO_0/CONFIG_reg[17][5] ));
    CFG3 #( .INIT(8'hF8) )  
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_142_rs_RNIO2KU  (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_45_set_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_142_rs_net_1 ), .C(
        \reg_apb_wrp_0/reg16x8_0/mem_1_rs[6] ), .Y(
        \reg_apb_wrp_0/reg16x8_0/mem_1_[6]_net_1 ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_163  (.A(VCC), 
        .B(VCC), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/SPI1_SDO_F2H_SCP_net ), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/SPI1_SS2_F2H_SCP_net ), .IPC());
    IOINFF_BYPASS \FIC_MSS_0/MDDR_DQ_8_PAD/U_IOINFF  (.A(
        \FIC_MSS_0/MDDR_DQ_8_PAD_Y ), .Y(\FIC_MSS_0/MDDR_DQ_8_PAD/YIN )
        );
    CFG2 #( .INIT(4'h6) )  
        \CoreGPIO_0/xhdl1.GEN_BITS[3].APB_32.edge_both_51_iv_0_x2[3]  
        (.A(\CoreGPIO_0/gpin2[3] ), .B(
        \CoreGPIO_0.xhdl1.GEN_BITS[3].gpin3[3] ), .Y(
        \CoreGPIO_0/N_253_i ));
    CFG4 #( .INIT(16'h0F35) )  
        \CoreGPIO_0/CONFIG_reg_o_2_31_am_1_RNO_1[1]  (.A(
        \CoreGPIO_0.xhdl1.GEN_BITS[4].REG_GEN.CONFIG_reg[4][1] ), .B(
        \CoreGPIO_0/CONFIG_reg[20][1] ), .C(
        \CoreAPB3_0_APBmslave3_PADDR[6] ), .D(
        \CoreAPB3_0_APBmslave3_PADDR[5] ), .Y(
        \CoreGPIO_0/CONFIG_reg_o_2_6_1[1] ));
    CFG2 #( .INIT(4'h2) )  
        \reg_apb_wrp_0/reg16x8_0/temp_data_2_15_i_a3_13[6]  (.A(
        \reg_apb_wrp_0/reg16x8_0/N_499 ), .B(
        \reg_apb_wrp_0/reg16x8_0/mem_8_[6]_net_1 ), .Y(
        \reg_apb_wrp_0/reg16x8_0/N_460 ));
    IP_INTERFACE \FIC_MSS_0/MSS_ADLIB_INST/IP_INTERFACE_255  (.A(VCC), 
        .B(VCC), .C(VCC), .IPA(
        \FIC_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[3] ), .IPB(
        \FIC_MSS_0/MSS_ADLIB_INST/F_ARADDR_HADDR1_net[15] ), .IPC());
    CFG2 #( .INIT(4'h4) )  \CoreGPIO_0/PRDATA_0_iv_0_a2_0[17]  (.A(
        \CoreGPIO_0.N_247 ), .B(\CoreGPIO_0/INTR_reg[17] ), .Y(
        \CoreGPIO_0.N_552 ));
    CFG4 #( .INIT(16'hAC0F) )  
        \CoreGPIO_0/CONFIG_reg_o_2_31_am_1_RNO_0[5]  (.A(
        \CoreGPIO_0/CONFIG_reg[8][5] ), .B(
        \CoreGPIO_0/CONFIG_reg[24][5] ), .C(
        \CoreGPIO_0/CONFIG_reg_o_2_3_1[5] ), .D(
        \CoreAPB3_0_APBmslave3_PADDR[5] ), .Y(
        \CoreGPIO_0/CONFIG_reg_o_2_31_am_1_RNO_0[5]_net_1 ));
    INV_BA AFLSDF_INV_33 (.A(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_8_net_1 ), .Y(
        AFLSDF_INV_33_net_1));
    CFG4 #( .INIT(16'h0F35) )  
        \CoreGPIO_0/CONFIG_reg_o_2_31_bm_1_RNO_2[6]  (.A(
        \CoreGPIO_0/CONFIG_reg[1][6] ), .B(
        \CoreGPIO_0/CONFIG_reg[17][6] ), .C(
        \CoreAPB3_0_APBmslave3_PADDR[6] ), .D(
        \CoreAPB3_0_APBmslave3_PADDR[5] ), .Y(
        \CoreGPIO_0/CONFIG_reg_o_2_18_1[6] ));
    CFG3 #( .INIT(8'h02) )  \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_109  
        (.A(\reg_apb_wrp_0/reg16x8_0/mem_13_[5]_net_1 ), .B(
        \reg_apb_wrp_0/reg16x8_0/N_500 ), .C(MSS_RESET_N_F2M_ibuf), .Y(
        \reg_apb_wrp_0/reg16x8_0/un1_mem_0_5_109_net_1 ));
    GND GND_power_inst1 (.Y(GND_power_net1));
    VCC VCC_power_inst1 (.Y(VCC_power_net1));
    
endmodule
