// ********************************************************************/
// Actel Corporation Proprietary and Confidential
//  Copyright 2011 Actel Corporation.  All rights reserved.
//
// ANY USE OR REDISTRIBUTION IN PART OR IN WHOLE MUST BE HANDLED IN
// ACCORDANCE WITH THE ACTEL LICENSE AGREEMENT AND MUST BE APPROVED
// IN ADVANCE IN WRITING.
//
// Description:  SRAM block, 4 byte wide, 512 to 35328 deep (in steps
//               of 512), used to construct the memory.
//
// Revision Information:
// Date     Description
//
// SVN Revision Information:
// SVN $Revision: 4805 $
// SVN $Date: 2008-11-27 17:48:48 +0530 (Thu, 27 Nov 2008) $
//
// Resolved SARs
// SAR      Date     Who   Description
//
// Notes:
//
// ********************************************************************/

`timescale 1ns/100ps

module FIC_COREAPBLSRAM_0_lsram_512to35328x32
(
    writeData,
    readData,
    wen,
    ren,
    writeAddr,
    readAddr,
    clk,
    resetn,
    lsram_512_BUSY_all
);

// ---------------------------------------------------------------------
// Parameters
// ---------------------------------------------------------------------
// DEPTH can range from 512 to 8192, in steps of 512
parameter DEPTH = 512;
parameter APB_DWIDTH = 32;

// ---------------------------------------------------------------------
// Port declarations
// ---------------------------------------------------------------------

   // ApbFabric interface
   // Inputs
   input [APB_DWIDTH-1:0] writeData;

   // AhbSramIf interface
   // Inputs
   input                  wen;
   input                  ren;
   input [17:0]           writeAddr;
   input [17:0]           readAddr;
   input                  clk;
   input                  resetn;

    // Output
   output                  lsram_512_BUSY_all;
   output [APB_DWIDTH-1:0] readData;

   reg [APB_DWIDTH-1:0]    readData;
   


// ---------------------------------------------------------------------
// Constant declarations
// ---------------------------------------------------------------------

// ---------------------------------------------------------------------
// Signal declarations
// ---------------------------------------------------------------------
        reg     [17:9]                  ckRdAddr;

        reg     [2:0]                   width0;
        reg     [2:0]                   width1;
        reg     [2:0]                   width2;
        reg     [2:0]                   width3;
        reg     [2:0]                   width4;
        reg     [2:0]                   width5;
        reg     [2:0]                   width6;
        reg     [2:0]                   width7;
        reg     [2:0]                   width8;
        reg     [2:0]                   width9;
        reg     [2:0]                   width10;
        reg     [2:0]                   width11;
        reg     [2:0]                   width12;
        reg     [2:0]                   width13;
        reg     [2:0]                   width14;
        reg     [2:0]                   width15;
        reg     [2:0]                   width16;
        reg     [2:0]                   width17;
        reg     [2:0]                   width18;
        reg     [2:0]                   width19;
        reg     [2:0]                   width20;
        reg     [2:0]                   width21;
        reg     [2:0]                   width22;
        reg     [2:0]                   width23;
        reg     [2:0]                   width24;
        reg     [2:0]                   width25;
        reg     [2:0]                   width26;
        reg     [2:0]                   width27;
        reg     [2:0]                   width28;
        reg     [2:0]                   width29;
        reg     [2:0]                   width30;
        reg     [2:0]                   width31;
        reg     [2:0]                   width32;
        reg     [2:0]                   width33;
        reg     [2:0]                   width34;
        reg     [2:0]                   width35;
        reg     [2:0]                   width36;
        reg     [2:0]                   width37;
        reg     [2:0]                   width38;
        reg     [2:0]                   width39;
        reg     [2:0]                   width40;
        reg     [2:0]                   width41;
        reg     [2:0]                   width42;
        reg     [2:0]                   width43;
        reg     [2:0]                   width44;
        reg     [2:0]                   width45;
        reg     [2:0]                   width46;
        reg     [2:0]                   width47;
        reg     [2:0]                   width48;
        reg     [2:0]                   width49;
        reg     [2:0]                   width50;
        reg     [2:0]                   width51;
        reg     [2:0]                   width52;
        reg     [2:0]                   width53;
        reg     [2:0]                   width54;
        reg     [2:0]                   width55;
        reg     [2:0]                   width56;
        reg     [2:0]                   width57;
        reg     [2:0]                   width58;
        reg     [2:0]                   width59;
        reg     [2:0]                   width60;
        reg     [2:0]                   width61;
        reg     [2:0]                   width62;
        reg     [2:0]                   width63;
        reg     [2:0]                   width64;
        reg     [2:0]                   width65;
        reg     [2:0]                   width66;
        reg     [2:0]                   width67;
        reg     [2:0]                   width68;


        reg     [1:0]                   wen_a0;
        reg     [1:0]                   wen_a1;
        reg     [1:0]                   wen_a2;
        reg     [1:0]                   wen_a3;
        reg     [1:0]                   wen_a4;
        reg     [1:0]                   wen_a5;
        reg     [1:0]                   wen_a6;
        reg     [1:0]                   wen_a7;
        reg     [1:0]                   wen_a8;
        reg     [1:0]                   wen_a9;
        reg     [1:0]                   wen_a10;
        reg     [1:0]                   wen_a11;
        reg     [1:0]                   wen_a12;
        reg     [1:0]                   wen_a13;
        reg     [1:0]                   wen_a14;
        reg     [1:0]                   wen_a15;
        reg     [1:0]                   wen_a16;
        reg     [1:0]                   wen_a17;
        reg     [1:0]                   wen_a18;
        reg     [1:0]                   wen_a19;
        reg     [1:0]                   wen_a20;
        reg     [1:0]                   wen_a21;
        reg     [1:0]                   wen_a22;
        reg     [1:0]                   wen_a23;
        reg     [1:0]                   wen_a24;
        reg     [1:0]                   wen_a25;
        reg     [1:0]                   wen_a26;
        reg     [1:0]                   wen_a27;
        reg     [1:0]                   wen_a28;
        reg     [1:0]                   wen_a29;
        reg     [1:0]                   wen_a30;
        reg     [1:0]                   wen_a31;
        reg     [1:0]                   wen_a32;
        reg     [1:0]                   wen_a33;
        reg     [1:0]                   wen_a34;
        reg     [1:0]                   wen_a35;
        reg     [1:0]                   wen_a36;
        reg     [1:0]                   wen_a37;
        reg     [1:0]                   wen_a38;
        reg     [1:0]                   wen_a39;
        reg     [1:0]                   wen_a40;
        reg     [1:0]                   wen_a41;
        reg     [1:0]                   wen_a42;
        reg     [1:0]                   wen_a43;
        reg     [1:0]                   wen_a44;
        reg     [1:0]                   wen_a45;
        reg     [1:0]                   wen_a46;
        reg     [1:0]                   wen_a47;
        reg     [1:0]                   wen_a48;
        reg     [1:0]                   wen_a49;
        reg     [1:0]                   wen_a50;
        reg     [1:0]                   wen_a51;
        reg     [1:0]                   wen_a52;
        reg     [1:0]                   wen_a53;
        reg     [1:0]                   wen_a54;
        reg     [1:0]                   wen_a55;
        reg     [1:0]                   wen_a56;
        reg     [1:0]                   wen_a57;
        reg     [1:0]                   wen_a58;
        reg     [1:0]                   wen_a59;
        reg     [1:0]                   wen_a60;
        reg     [1:0]                   wen_a61;
        reg     [1:0]                   wen_a62;
        reg     [1:0]                   wen_a63;
        reg     [1:0]                   wen_a64;
        reg     [1:0]                   wen_a65;
        reg     [1:0]                   wen_a66;
        reg     [1:0]                   wen_a67;
        reg     [1:0]                   wen_a68;

        reg     [1:0]                   wen_b0;
        reg     [1:0]                   wen_b1;
        reg     [1:0]                   wen_b2;
        reg     [1:0]                   wen_b3;
        reg     [1:0]                   wen_b4;
        reg     [1:0]                   wen_b5;
        reg     [1:0]                   wen_b6;
        reg     [1:0]                   wen_b7;
        reg     [1:0]                   wen_b8;
        reg     [1:0]                   wen_b9;
        reg     [1:0]                   wen_b10;
        reg     [1:0]                   wen_b11;
        reg     [1:0]                   wen_b12;
        reg     [1:0]                   wen_b13;
        reg     [1:0]                   wen_b14;
        reg     [1:0]                   wen_b15;
        reg     [1:0]                   wen_b16;
        reg     [1:0]                   wen_b17;
        reg     [1:0]                   wen_b18;
        reg     [1:0]                   wen_b19;
        reg     [1:0]                   wen_b20;
        reg     [1:0]                   wen_b21;
        reg     [1:0]                   wen_b22;
        reg     [1:0]                   wen_b23;
        reg     [1:0]                   wen_b24;
        reg     [1:0]                   wen_b25;
        reg     [1:0]                   wen_b26;
        reg     [1:0]                   wen_b27;
        reg     [1:0]                   wen_b28;
        reg     [1:0]                   wen_b29;
        reg     [1:0]                   wen_b30;
        reg     [1:0]                   wen_b31;
        reg     [1:0]                   wen_b32;
        reg     [1:0]                   wen_b33;
        reg     [1:0]                   wen_b34;
        reg     [1:0]                   wen_b35;
        reg     [1:0]                   wen_b36;
        reg     [1:0]                   wen_b37;
        reg     [1:0]                   wen_b38;
        reg     [1:0]                   wen_b39;
        reg     [1:0]                   wen_b40;
        reg     [1:0]                   wen_b41;
        reg     [1:0]                   wen_b42;
        reg     [1:0]                   wen_b43;
        reg     [1:0]                   wen_b44;
        reg     [1:0]                   wen_b45;
        reg     [1:0]                   wen_b46;
        reg     [1:0]                   wen_b47;
        reg     [1:0]                   wen_b48;
        reg     [1:0]                   wen_b49;
        reg     [1:0]                   wen_b50;
        reg     [1:0]                   wen_b51;
        reg     [1:0]                   wen_b52;
        reg     [1:0]                   wen_b53;
        reg     [1:0]                   wen_b54;
        reg     [1:0]                   wen_b55;
        reg     [1:0]                   wen_b56;
        reg     [1:0]                   wen_b57;
        reg     [1:0]                   wen_b58;
        reg     [1:0]                   wen_b59;
        reg     [1:0]                   wen_b60;
        reg     [1:0]                   wen_b61;
        reg     [1:0]                   wen_b62;
        reg     [1:0]                   wen_b63;
        reg     [1:0]                   wen_b64;
        reg     [1:0]                   wen_b65;
        reg     [1:0]                   wen_b66;
        reg     [1:0]                   wen_b67;
        reg     [1:0]                   wen_b68;

        reg     [35:0]                   writeData0;
        reg     [17:0]                   writeData1;
        reg     [17:0]                   writeData2;
        reg     [17:0]                   writeData3;
        reg     [17:0]                   writeData4;
        reg     [17:0]                   writeData5;
        reg     [17:0]                   writeData6;
        reg     [17:0]                   writeData7;
        reg     [17:0]                   writeData8;
        reg     [17:0]                   writeData9;
        reg     [17:0]                   writeData10;
        reg     [17:0]                   writeData11;
        reg     [17:0]                   writeData12;
        reg     [17:0]                   writeData13;
        reg     [17:0]                   writeData14;
        reg     [17:0]                   writeData15;
        reg     [17:0]                   writeData16;
        reg     [17:0]                   writeData17;
        reg     [17:0]                   writeData18;
        reg     [17:0]                   writeData19;
        reg     [17:0]                   writeData20;
        reg     [17:0]                   writeData21;
        reg     [17:0]                   writeData22;
        reg     [17:0]                   writeData23;
        reg     [17:0]                   writeData24;
        reg     [17:0]                   writeData25;
        reg     [17:0]                   writeData26;
        reg     [17:0]                   writeData27;
        reg     [17:0]                   writeData28;
        reg     [17:0]                   writeData29;
        reg     [17:0]                   writeData30;
        reg     [17:0]                   writeData31;
        reg     [17:0]                   writeData32;
        reg     [17:0]                   writeData33;
        reg     [17:0]                   writeData34;
        reg     [17:0]                   writeData35;
        reg     [17:0]                   writeData36;
        reg     [17:0]                   writeData37;
        reg     [17:0]                   writeData38;
        reg     [17:0]                   writeData39;
        reg     [17:0]                   writeData40;
        reg     [17:0]                   writeData41;
        reg     [17:0]                   writeData42;
        reg     [17:0]                   writeData43;
        reg     [17:0]                   writeData44;
        reg     [17:0]                   writeData45;
        reg     [17:0]                   writeData46;
        reg     [17:0]                   writeData47;
        reg     [17:0]                   writeData48;
        reg     [17:0]                   writeData49;
        reg     [17:0]                   writeData50;
        reg     [17:0]                   writeData51;
        reg     [17:0]                   writeData52;
        reg     [17:0]                   writeData53;
        reg     [17:0]                   writeData54;
        reg     [17:0]                   writeData55;
        reg     [17:0]                   writeData56;
        reg     [17:0]                   writeData57;
        reg     [17:0]                   writeData58;
        reg     [17:0]                   writeData59;
        reg     [17:0]                   writeData60;
        reg     [17:0]                   writeData61;
        reg     [17:0]                   writeData62;
        reg     [17:0]                   writeData63;
        reg     [17:0]                   writeData64;
        reg     [17:0]                   writeData65;
        reg     [17:0]                   writeData66;
        reg     [17:0]                   writeData67;
        reg     [17:0]                   writeData68;

        wire    [35:0]                   readData0;
        wire    [17:0]                   readData1;
        wire    [17:0]                   readData2;
        wire    [17:0]                   readData3;
        wire    [17:0]                   readData4;
        wire    [17:0]                   readData5;
        wire    [17:0]                   readData6;
        wire    [17:0]                   readData7;
        wire    [17:0]                   readData8;
        wire    [17:0]                   readData9;
        wire    [17:0]                   readData10;
        wire    [17:0]                   readData11;
        wire    [17:0]                   readData12;
        wire    [17:0]                   readData13;
        wire    [17:0]                   readData14;
        wire    [17:0]                   readData15;
        wire    [17:0]                   readData16;
        wire    [17:0]                   readData17;
        wire    [17:0]                   readData18;
        wire    [17:0]                   readData19;
        wire    [17:0]                   readData20;
        wire    [17:0]                   readData21;
        wire    [17:0]                   readData22;
        wire    [17:0]                   readData23;
        wire    [17:0]                   readData24;
        wire    [17:0]                   readData25;
        wire    [17:0]                   readData26;
        wire    [17:0]                   readData27;
        wire    [17:0]                   readData28;
        wire    [17:0]                   readData29;
        wire    [17:0]                   readData30;
        wire    [17:0]                   readData31;
        wire    [17:0]                   readData32;
        wire    [17:0]                   readData33;
        wire    [17:0]                   readData34;
        wire    [17:0]                   readData35;
        wire    [17:0]                   readData36;
        wire    [17:0]                   readData37;
        wire    [17:0]                   readData38;
        wire    [17:0]                   readData39;
        wire    [17:0]                   readData40;
        wire    [17:0]                   readData41;
        wire    [17:0]                   readData42;
        wire    [17:0]                   readData43;
        wire    [17:0]                   readData44;
        wire    [17:0]                   readData45;
        wire    [17:0]                   readData46;
        wire    [17:0]                   readData47;
        wire    [17:0]                   readData48;
        wire    [17:0]                   readData49;
        wire    [17:0]                   readData50;
        wire    [17:0]                   readData51;
        wire    [17:0]                   readData52;
        wire    [17:0]                   readData53;
        wire    [17:0]                   readData54;
        wire    [17:0]                   readData55;
        wire    [17:0]                   readData56;
        wire    [17:0]                   readData57;
        wire    [17:0]                   readData58;
        wire    [17:0]                   readData59;
        wire    [17:0]                   readData60;
        wire    [17:0]                   readData61;
        wire    [17:0]                   readData62;
        wire    [17:0]                   readData63;
        wire    [17:0]                   readData64;
        wire    [17:0]                   readData65;
        wire    [17:0]                   readData66;
        wire    [17:0]                   readData67;
        wire    [17:0]                   readData68;

        reg     [13:0]                  writeAddr0;
        reg     [13:0]                  writeAddr1;
        reg     [13:0]                  writeAddr2;
        reg     [13:0]                  writeAddr3;
        reg     [13:0]                  writeAddr4;
        reg     [13:0]                  writeAddr5;
        reg     [13:0]                  writeAddr6;
        reg     [13:0]                  writeAddr7;
        reg     [13:0]                  writeAddr8;
        reg     [13:0]                  writeAddr9;
        reg     [13:0]                  writeAddr10;
        reg     [13:0]                  writeAddr11;
        reg     [13:0]                  writeAddr12;
        reg     [13:0]                  writeAddr13;
        reg     [13:0]                  writeAddr14;
        reg     [13:0]                  writeAddr15;
        reg     [13:0]                  writeAddr16;
        reg     [13:0]                  writeAddr17;
        reg     [13:0]                  writeAddr18;
        reg     [13:0]                  writeAddr19;
        reg     [13:0]                  writeAddr20;
        reg     [13:0]                  writeAddr21;
        reg     [13:0]                  writeAddr22;
        reg     [13:0]                  writeAddr23;
        reg     [13:0]                  writeAddr24;
        reg     [13:0]                  writeAddr25;
        reg     [13:0]                  writeAddr26;
        reg     [13:0]                  writeAddr27;
        reg     [13:0]                  writeAddr28;
        reg     [13:0]                  writeAddr29;
        reg     [13:0]                  writeAddr30;
        reg     [13:0]                  writeAddr31;
        reg     [13:0]                  writeAddr32;
        reg     [13:0]                  writeAddr33;
        reg     [13:0]                  writeAddr34;
        reg     [13:0]                  writeAddr35;
        reg     [13:0]                  writeAddr36;
        reg     [13:0]                  writeAddr37;
        reg     [13:0]                  writeAddr38;
        reg     [13:0]                  writeAddr39;
        reg     [13:0]                  writeAddr40;
        reg     [13:0]                  writeAddr41;
        reg     [13:0]                  writeAddr42;
        reg     [13:0]                  writeAddr43;
        reg     [13:0]                  writeAddr44;
        reg     [13:0]                  writeAddr45;
        reg     [13:0]                  writeAddr46;
        reg     [13:0]                  writeAddr47;
        reg     [13:0]                  writeAddr48;
        reg     [13:0]                  writeAddr49;
        reg     [13:0]                  writeAddr50;
        reg     [13:0]                  writeAddr51;
        reg     [13:0]                  writeAddr52;
        reg     [13:0]                  writeAddr53;
        reg     [13:0]                  writeAddr54;
        reg     [13:0]                  writeAddr55;
        reg     [13:0]                  writeAddr56;
        reg     [13:0]                  writeAddr57;
        reg     [13:0]                  writeAddr58;
        reg     [13:0]                  writeAddr59;
        reg     [13:0]                  writeAddr60;
        reg     [13:0]                  writeAddr61;
        reg     [13:0]                  writeAddr62;
        reg     [13:0]                  writeAddr63;
        reg     [13:0]                  writeAddr64;
        reg     [13:0]                  writeAddr65;
        reg     [13:0]                  writeAddr66;
        reg     [13:0]                  writeAddr67;
        reg     [13:0]                  writeAddr68;

        reg     [13:0]                  readAddr0;
        reg     [13:0]                  readAddr1;
        reg     [13:0]                  readAddr2;
        reg     [13:0]                  readAddr3;
        reg     [13:0]                  readAddr4;
        reg     [13:0]                  readAddr5;
        reg     [13:0]                  readAddr6;
        reg     [13:0]                  readAddr7;
        reg     [13:0]                  readAddr8;
        reg     [13:0]                  readAddr9;
        reg     [13:0]                  readAddr10;
        reg     [13:0]                  readAddr11;
        reg     [13:0]                  readAddr12;
        reg     [13:0]                  readAddr13;
        reg     [13:0]                  readAddr14;
        reg     [13:0]                  readAddr15;
        reg     [13:0]                  readAddr16;
        reg     [13:0]                  readAddr17;
        reg     [13:0]                  readAddr18;
        reg     [13:0]                  readAddr19;
        reg     [13:0]                  readAddr20;
        reg     [13:0]                  readAddr21;
        reg     [13:0]                  readAddr22;
        reg     [13:0]                  readAddr23;
        reg     [13:0]                  readAddr24;
        reg     [13:0]                  readAddr25;
        reg     [13:0]                  readAddr26;
        reg     [13:0]                  readAddr27;
        reg     [13:0]                  readAddr28;
        reg     [13:0]                  readAddr29;
        reg     [13:0]                  readAddr30;
        reg     [13:0]                  readAddr31;
        reg     [13:0]                  readAddr32;
        reg     [13:0]                  readAddr33;
        reg     [13:0]                  readAddr34;
        reg     [13:0]                  readAddr35;
        reg     [13:0]                  readAddr36;
        reg     [13:0]                  readAddr37;
        reg     [13:0]                  readAddr38;
        reg     [13:0]                  readAddr39;
        reg     [13:0]                  readAddr40;
        reg     [13:0]                  readAddr41;
        reg     [13:0]                  readAddr42;
        reg     [13:0]                  readAddr43;
        reg     [13:0]                  readAddr44;
        reg     [13:0]                  readAddr45;
        reg     [13:0]                  readAddr46;
        reg     [13:0]                  readAddr47;
        reg     [13:0]                  readAddr48;
        reg     [13:0]                  readAddr49;
        reg     [13:0]                  readAddr50;
        reg     [13:0]                  readAddr51;
        reg     [13:0]                  readAddr52;
        reg     [13:0]                  readAddr53;
        reg     [13:0]                  readAddr54;
        reg     [13:0]                  readAddr55;
        reg     [13:0]                  readAddr56;
        reg     [13:0]                  readAddr57;
        reg     [13:0]                  readAddr58;
        reg     [13:0]                  readAddr59;
        reg     [13:0]                  readAddr60;
        reg     [13:0]                  readAddr61;
        reg     [13:0]                  readAddr62;
        reg     [13:0]                  readAddr63;
        reg     [13:0]                  readAddr64;
        reg     [13:0]                  readAddr65;
        reg     [13:0]                  readAddr66;
        reg     [13:0]                  readAddr67;
        reg     [11:0]                  readAddr68;


   wire                                 lsram_512_BUSY_all;
   wire                                 lsram_512_BUSY_68;
   wire                                 lsram_512_BUSY_67;
   wire                                 lsram_512_BUSY_66;
   wire                                 lsram_512_BUSY_65;
   wire                                 lsram_512_BUSY_64;
   wire                                 lsram_512_BUSY_63;
   wire                                 lsram_512_BUSY_62;
   wire                                 lsram_512_BUSY_61;
   wire                                 lsram_512_BUSY_60;
   wire                                 lsram_512_BUSY_59;
   wire                                 lsram_512_BUSY_58;
   wire                                 lsram_512_BUSY_57;
   wire                                 lsram_512_BUSY_56;
   wire                                 lsram_512_BUSY_55;
   wire                                 lsram_512_BUSY_54;
   wire                                 lsram_512_BUSY_53;
   wire                                 lsram_512_BUSY_52;
   wire                                 lsram_512_BUSY_51;
   wire                                 lsram_512_BUSY_50;
   wire                                 lsram_512_BUSY_49;
   wire                                 lsram_512_BUSY_48;
   wire                                 lsram_512_BUSY_47;
   wire                                 lsram_512_BUSY_46;
   wire                                 lsram_512_BUSY_45;
   wire                                 lsram_512_BUSY_44;
   wire                                 lsram_512_BUSY_43;
   wire                                 lsram_512_BUSY_42;
   wire                                 lsram_512_BUSY_41;
   wire                                 lsram_512_BUSY_40;
   wire                                 lsram_512_BUSY_39;
   wire                                 lsram_512_BUSY_38;
   wire                                 lsram_512_BUSY_37;
   wire                                 lsram_512_BUSY_36;
   wire                                 lsram_512_BUSY_35;
   wire                                 lsram_512_BUSY_34;
   wire                                 lsram_512_BUSY_33;
   wire                                 lsram_512_BUSY_32;
   wire                                 lsram_512_BUSY_31;
   wire                                 lsram_512_BUSY_30;
   wire                                 lsram_512_BUSY_29;
   wire                                 lsram_512_BUSY_28;
   wire                                 lsram_512_BUSY_27;
   wire                                 lsram_512_BUSY_26;
   wire                                 lsram_512_BUSY_25;
   wire                                 lsram_512_BUSY_24;
   wire                                 lsram_512_BUSY_23;
   wire                                 lsram_512_BUSY_22;
   wire                                 lsram_512_BUSY_21;
   wire                                 lsram_512_BUSY_20;
   wire                                 lsram_512_BUSY_19;
   wire                                 lsram_512_BUSY_18;
   wire                                 lsram_512_BUSY_17;
   wire                                 lsram_512_BUSY_16;
   wire                                 lsram_512_BUSY_15;
   wire                                 lsram_512_BUSY_14;
   wire                                 lsram_512_BUSY_13;
   wire                                 lsram_512_BUSY_12;
   wire                                 lsram_512_BUSY_11;
   wire                                 lsram_512_BUSY_10;
   wire                                 lsram_512_BUSY_9;
   wire                                 lsram_512_BUSY_8;
   wire                                 lsram_512_BUSY_7;
   wire                                 lsram_512_BUSY_6;
   wire                                 lsram_512_BUSY_5;
   wire                                 lsram_512_BUSY_4;
   wire                                 lsram_512_BUSY_3;
   wire                                 lsram_512_BUSY_2;
   wire                                 lsram_512_BUSY_1;
   wire                                 lsram_512_BUSY_0;
   

//----------------------------------------------------------------------
// Main body of code
//----------------------------------------------------------------------

    always @ (posedge clk or negedge resetn)
    begin
        if (!resetn)
            ckRdAddr[15:9] <= 7'b0000000;
        else
            ckRdAddr[15:9] <= readAddr[15:9];
    end

    //----------------------------------------------------------------------------------------
    // Assign values to various signals based on DEPTH and RAM4K9_WIDTH settings.
    // Default is to build the (byte wide) memory from RAM blocks which are configured to
    // be tall and narrow.
    //----------------------------------------------------------------------------------------
    always @(*)
    begin
       readData = {APB_DWIDTH{1'b0}};
        width0  = 2'b0;
        width1  = 2'b0;
        width2  = 2'b0;
        width3  = 2'b0;
        width4  = 2'b0;
        width5  = 2'b0;
        width6  = 2'b0;
        width7  = 2'b0;
        width8  = 2'b0;
        width9  = 2'b0;
        width10 = 2'b0;
        width11 = 2'b0;
        width12 = 2'b0;
        width13 = 2'b0;
        width14 = 2'b0;
        width15 = 2'b0;
        width16 = 2'b0;
        width17 = 2'b0;
        width18 = 2'b0;
        width19 = 2'b0;
        width20 = 2'b0;
        width21 = 2'b0;
        width22 = 2'b0;
        width23 = 2'b0;
        width24 = 2'b0;
        width25 = 2'b0;
        width26 = 2'b0;
        width27 = 2'b0;
        width28 = 2'b0;
        width29 = 2'b0;
        width30 = 2'b0;
        width31 = 2'b0;
        width32 = 2'b0;
        width33 = 2'b0;
        width34 = 2'b0;
        width35 = 2'b0;
        width36 = 2'b0;
        width37 = 2'b0;
        width38 = 2'b0;
        width39 = 2'b0;
        width40 = 2'b0;
        width41 = 2'b0;
        width42 = 2'b0;
        width43 = 2'b0;
        width44 = 2'b0;
        width45 = 2'b0;
        width46 = 2'b0;
        width47 = 2'b0;
        width48 = 2'b0;
        width49 = 2'b0;
        width50 = 2'b0;
        width51 = 2'b0;
        width52 = 2'b0;
        width53 = 2'b0;
        width54 = 2'b0;
        width55 = 2'b0;
        width56 = 2'b0;
        width57 = 2'b0;
        width58 = 2'b0;
        width59 = 2'b0;
        width60 = 2'b0;
        width61 = 2'b0;
        width62 = 2'b0;
        width63 = 2'b0;
        width64 = 2'b0;
        width65 = 2'b0;
        width66 = 2'b0;
        width67 = 2'b0;
        width68 = 2'b0;

        wen_a0  = 2'b0;
        wen_a1  = 2'b0;
        wen_a2  = 2'b0;
        wen_a3  = 2'b0;
        wen_a4  = 2'b0;
        wen_a5  = 2'b0;
        wen_a6  = 2'b0;
        wen_a7  = 2'b0;
        wen_a8  = 2'b0;
        wen_a9  = 2'b0;
        wen_a10 = 2'b0;
        wen_a11 = 2'b0;
        wen_a12 = 2'b0;
        wen_a13 = 2'b0;
        wen_a14 = 2'b0;
        wen_a15 = 2'b0;
        wen_a16 = 2'b0;
        wen_a17 = 2'b0;
        wen_a18 = 2'b0;
        wen_a19 = 2'b0;
        wen_a20 = 2'b0;
        wen_a21 = 2'b0;
        wen_a22 = 2'b0;
        wen_a23 = 2'b0;
        wen_a24 = 2'b0;
        wen_a25 = 2'b0;
        wen_a26 = 2'b0;
        wen_a27 = 2'b0;
        wen_a28 = 2'b0;
        wen_a29 = 2'b0;
        wen_a30 = 2'b0;
        wen_a31 = 2'b0;
        wen_a32 = 2'b0;
        wen_a33 = 2'b0;
        wen_a34 = 2'b0;
        wen_a35 = 2'b0;
        wen_a36 = 2'b0;
        wen_a37 = 2'b0;
        wen_a38 = 2'b0;
        wen_a39 = 2'b0;
        wen_a40 = 2'b0;
        wen_a41 = 2'b0;
        wen_a42 = 2'b0;
        wen_a43 = 2'b0;
        wen_a44 = 2'b0;
        wen_a45 = 2'b0;
        wen_a46 = 2'b0;
        wen_a47 = 2'b0;
        wen_a48 = 2'b0;
        wen_a49 = 2'b0;
        wen_a50 = 2'b0;
        wen_a51 = 2'b0;
        wen_a52 = 2'b0;
        wen_a53 = 2'b0;
        wen_a54 = 2'b0;
        wen_a55 = 2'b0;
        wen_a56 = 2'b0;
        wen_a57 = 2'b0;
        wen_a58 = 2'b0;
        wen_a59 = 2'b0;
        wen_a60 = 2'b0;
        wen_a61 = 2'b0;
        wen_a62 = 2'b0;
        wen_a63 = 2'b0;
        wen_a64 = 2'b0;
        wen_a65 = 2'b0;
        wen_a66 = 2'b0;
        wen_a67 = 2'b0;
        wen_a68 = 2'b0;

        wen_b0  = 2'b0;
        wen_b1  = 2'b0;
        wen_b2  = 2'b0;
        wen_b3  = 2'b0;
        wen_b4  = 2'b0;
        wen_b5  = 2'b0;
        wen_b6  = 2'b0;
        wen_b7  = 2'b0;
        wen_b8  = 2'b0;
        wen_b9  = 2'b0;
        wen_b10 = 2'b0;
        wen_b11 = 2'b0;
        wen_b12 = 2'b0;
        wen_b13 = 2'b0;
        wen_b14 = 2'b0;
        wen_b15 = 2'b0;
        wen_b16 = 2'b0;
        wen_b17 = 2'b0;
        wen_b18 = 2'b0;
        wen_b19 = 2'b0;
        wen_b20 = 2'b0;
        wen_b21 = 2'b0;
        wen_b22 = 2'b0;
        wen_b23 = 2'b0;
        wen_b24 = 2'b0;
        wen_b25 = 2'b0;
        wen_b26 = 2'b0;
        wen_b27 = 2'b0;
        wen_b28 = 2'b0;
        wen_b29 = 2'b0;
        wen_b30 = 2'b0;
        wen_b31 = 2'b0;
        wen_b32 = 2'b0;
        wen_b33 = 2'b0;
        wen_b34 = 2'b0;
        wen_b35 = 2'b0;
        wen_b36 = 2'b0;
        wen_b37 = 2'b0;
        wen_b38 = 2'b0;
        wen_b39 = 2'b0;
        wen_b40 = 2'b0;
        wen_b41 = 2'b0;
        wen_b42 = 2'b0;
        wen_b43 = 2'b0;
        wen_b44 = 2'b0;
        wen_b45 = 2'b0;
        wen_b46 = 2'b0;
        wen_b47 = 2'b0;
        wen_b48 = 2'b0;
        wen_b49 = 2'b0;
        wen_b50 = 2'b0;
        wen_b51 = 2'b0;
        wen_b52 = 2'b0;
        wen_b53 = 2'b0;
        wen_b54 = 2'b0;
        wen_b55 = 2'b0;
        wen_b56 = 2'b0;
        wen_b57 = 2'b0;
        wen_b58 = 2'b0;
        wen_b59 = 2'b0;
        wen_b60 = 2'b0;
        wen_b61 = 2'b0;
        wen_b62 = 2'b0;
        wen_b63 = 2'b0;
        wen_b64 = 2'b0;
        wen_b65 = 2'b0;
        wen_b66 = 2'b0;
        wen_b67 = 2'b0;
        wen_b68 = 2'b0;

        writeData0  = 36'b0;
        writeData1  = 18'b0;
        writeData2  = 18'b0;
        writeData3  = 18'b0;
        writeData4  = 18'b0;
        writeData5  = 18'b0;
        writeData6  = 18'b0;
        writeData7  = 18'b0;
        writeData8  = 18'b0;
        writeData9  = 18'b0;
        writeData10 = 18'b0;
        writeData11 = 18'b0;
        writeData12 = 18'b0;
        writeData13 = 18'b0;
        writeData14 = 18'b0;
        writeData15 = 18'b0;
        writeData16 = 18'b0;
        writeData17 = 18'b0;
        writeData18 = 18'b0;
        writeData19 = 18'b0;
        writeData20 = 18'b0;
        writeData21 = 18'b0;
        writeData22 = 18'b0;
        writeData23 = 18'b0;
        writeData24 = 18'b0;
        writeData25 = 18'b0;
        writeData26 = 18'b0;
        writeData27 = 18'b0;
        writeData28 = 18'b0;
        writeData29 = 18'b0;
        writeData30 = 18'b0;
        writeData31 = 18'b0;
        writeData32 = 18'b0;
        writeData33 = 18'b0;
        writeData34 = 18'b0;
        writeData35 = 18'b0;
        writeData36 = 18'b0;
        writeData37 = 18'b0;
        writeData38 = 18'b0;
        writeData39 = 18'b0;
        writeData40 = 18'b0;
        writeData41 = 18'b0;
        writeData42 = 18'b0;
        writeData43 = 18'b0;
        writeData44 = 18'b0;
        writeData45 = 18'b0;
        writeData46 = 18'b0;
        writeData47 = 18'b0;
        writeData48 = 18'b0;
        writeData49 = 18'b0;
        writeData50 = 18'b0;
        writeData51 = 18'b0;
        writeData52 = 18'b0;
        writeData53 = 18'b0;
        writeData54 = 18'b0;
        writeData55 = 18'b0;
        writeData56 = 18'b0;
        writeData57 = 18'b0;
        writeData58 = 18'b0;
        writeData59 = 18'b0;
        writeData60 = 18'b0;
        writeData61 = 18'b0;
        writeData62 = 18'b0;
        writeData63 = 18'b0;
        writeData64 = 18'b0;
        writeData65 = 18'b0;
        writeData66 = 18'b0;
        writeData67 = 18'b0;
        writeData68 = 18'b0;

        writeAddr0  = 14'b0;
        writeAddr1  = 14'b0;
        writeAddr2  = 14'b0;
        writeAddr3  = 14'b0;
        writeAddr4  = 14'b0;
        writeAddr5  = 14'b0;
        writeAddr6  = 14'b0;
        writeAddr7  = 14'b0;
        writeAddr8  = 14'b0;
        writeAddr9  = 14'b0;
        writeAddr10 = 14'b0;
        writeAddr11 = 14'b0;
        writeAddr12 = 14'b0;
        writeAddr13 = 14'b0;
        writeAddr14 = 14'b0;
        writeAddr15 = 14'b0;
        writeAddr16 = 14'b0;
        writeAddr17 = 14'b0;
        writeAddr18 = 14'b0;
        writeAddr19 = 14'b0;
        writeAddr20 = 14'b0;
        writeAddr21 = 14'b0;
        writeAddr22 = 14'b0;
        writeAddr23 = 14'b0;
        writeAddr24 = 14'b0;
        writeAddr25 = 14'b0;
        writeAddr26 = 14'b0;
        writeAddr27 = 14'b0;
        writeAddr28 = 14'b0;
        writeAddr29 = 14'b0;
        writeAddr30 = 14'b0;
        writeAddr31 = 14'b0;
        writeAddr32 = 14'b0;
        writeAddr33 = 14'b0;
        writeAddr34 = 14'b0;
        writeAddr35 = 14'b0;
        writeAddr36 = 14'b0;
        writeAddr37 = 14'b0;
        writeAddr38 = 14'b0;
        writeAddr39 = 14'b0;
        writeAddr40 = 14'b0;
        writeAddr41 = 14'b0;
        writeAddr42 = 14'b0;
        writeAddr43 = 14'b0;
        writeAddr44 = 14'b0;
        writeAddr45 = 14'b0;
        writeAddr46 = 14'b0;
        writeAddr47 = 14'b0;
        writeAddr48 = 14'b0;
        writeAddr49 = 14'b0;
        writeAddr50 = 14'b0;
        writeAddr51 = 14'b0;
        writeAddr52 = 14'b0;
        writeAddr53 = 14'b0;
        writeAddr54 = 14'b0;
        writeAddr55 = 14'b0;
        writeAddr56 = 14'b0;
        writeAddr57 = 14'b0;
        writeAddr58 = 14'b0;
        writeAddr59 = 14'b0;
        writeAddr60 = 14'b0;
        writeAddr61 = 14'b0;
        writeAddr62 = 14'b0;
        writeAddr63 = 14'b0;
        writeAddr64 = 14'b0;
        writeAddr65 = 14'b0;
        writeAddr66 = 14'b0;
        writeAddr67 = 14'b0;
        writeAddr68 = 14'b0;

        readAddr0  = 14'b0;
        readAddr1  = 14'b0;
        readAddr2  = 14'b0;
        readAddr3  = 14'b0;
        readAddr4  = 14'b0;
        readAddr5  = 14'b0;
        readAddr6  = 14'b0;
        readAddr7  = 14'b0;
        readAddr8  = 14'b0;
        readAddr9  = 14'b0;
        readAddr10 = 14'b0;
        readAddr11 = 14'b0;
        readAddr12 = 14'b0;
        readAddr13 = 14'b0;
        readAddr14 = 14'b0;
        readAddr15 = 14'b0;
        readAddr16 = 14'b0;
        readAddr17 = 14'b0;
        readAddr18 = 14'b0;
        readAddr19 = 14'b0;
        readAddr20 = 14'b0;
        readAddr21 = 14'b0;
        readAddr22 = 14'b0;
        readAddr23 = 14'b0;
        readAddr24 = 14'b0;
        readAddr25 = 14'b0;
        readAddr26 = 14'b0;
        readAddr27 = 14'b0;
        readAddr28 = 14'b0;
        readAddr29 = 14'b0;
        readAddr30 = 14'b0;
        readAddr31 = 14'b0;
        readAddr32 = 14'b0;
        readAddr33 = 14'b0;
        readAddr34 = 14'b0;
        readAddr35 = 14'b0;
        readAddr36 = 14'b0;
        readAddr37 = 14'b0;
        readAddr38 = 14'b0;
        readAddr39 = 14'b0;
        readAddr40 = 14'b0;
        readAddr41 = 14'b0;
        readAddr42 = 14'b0;
        readAddr43 = 14'b0;
        readAddr44 = 14'b0;
        readAddr45 = 14'b0;
        readAddr46 = 14'b0;
        readAddr47 = 14'b0;
        readAddr48 = 14'b0;
        readAddr49 = 14'b0;
        readAddr50 = 14'b0;
        readAddr51 = 14'b0;
        readAddr52 = 14'b0;
        readAddr53 = 14'b0;
        readAddr54 = 14'b0;
        readAddr55 = 14'b0;
        readAddr56 = 14'b0;
        readAddr57 = 14'b0;
        readAddr58 = 14'b0;
        readAddr59 = 14'b0;
        readAddr60 = 14'b0;
        readAddr61 = 14'b0;
        readAddr62 = 14'b0;
        readAddr63 = 14'b0;
        readAddr64 = 14'b0;
        readAddr65 = 14'b0;
        readAddr66 = 14'b0;
        readAddr67 = 14'b0;
        readAddr68 = 14'b0;

        case (DEPTH)
            512: begin
                width0 = 3'b101;
                writeAddr0 = {writeAddr[8:0], 5'b0};
                readAddr0  = {readAddr[8:0],  5'b0};
                writeData0 = {1'b0, writeData[31:24], 1'b0, writeData[23:16], 1'b0, writeData[15:8], 1'b0, writeData[7:0]};
                wen_a0 = {wen, wen};
                wen_b0 = {wen, wen};
                readData = {readData0[34:27],readData0[25:18],readData0[16:9],readData0[7:0]};
            end
            1024: begin
                width2 = 3'b100;
                width1 = 3'b100;
                writeAddr2 = {writeAddr[9:0], 4'b0};
                writeAddr1 = {writeAddr[9:0], 4'b0};
                readAddr2  = {readAddr[9:0],  4'b0};
                readAddr1  = {readAddr[9:0],  4'b0};
                writeData2 = {1'b0, writeData[31:24], 1'b0, writeData[23:16]};
                writeData1 = {1'b0, writeData[15:8], 1'b0, writeData[7:0]};
                wen_a2 = {wen, wen};
                wen_a1 = {wen, wen};
                readData = {readData2[16:9],readData2[7:0],readData1[16:9],readData1[7:0]};
            end
            1536: begin
                width2 = 3'b100;
                width1 = 3'b100;
                width0 = 3'b101;
                writeAddr2 = {writeAddr[9:0], 4'b0};
                writeAddr1 = {writeAddr[9:0], 4'b0};
                writeAddr0 = {writeAddr[8:0], 5'b0};
                readAddr2  = {readAddr[9:0],  4'b0};
                readAddr1  = {readAddr[9:0],  4'b0};
                readAddr0  = {readAddr[8:0],  5'b0};
                writeData2 = {1'b0, writeData[31:24], 1'b0, writeData[23:16]};
                writeData1 = {1'b0, writeData[15:8], 1'b0, writeData[7:0]};
                writeData0 = {1'b0, writeData[31:24], 1'b0, writeData[23:16], 1'b0, writeData[15:8], 1'b0, writeData[7:0]};
                case (writeAddr[10:9])
                    2'b00, 2'b01 : {wen_a2, wen_a1, wen_a0, wen_b0} = {wen,  wen,  wen,  wen,  1'b0, 1'b0, 1'b0, 1'b0};
                    2'b10: {wen_a2, wen_a1, wen_a0, wen_b0} = {1'b0, 1'b0, 1'b0, 1'b0, wen,  wen, wen, wen};
                    default: {wen_a2, wen_a1, wen_a0, wen_b0} = {1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0};
                endcase
                case (ckRdAddr[10:9])
                    2'b00, 2'b01: readData = {readData2[16:9],readData2[7:0],readData1[16:9],readData1[7:0]};
                    2'b10: readData = {readData0[34:27],readData0[25:18],readData0[16:9],readData0[7:0]};
                    default: readData = 32'b0;
                endcase
            end
            2048: begin
                width4 = 3'b011;
                width3 = 3'b011;
                width2 = 3'b011;
                width1 = 3'b011;

                writeAddr4 = {writeAddr[10:0], 3'b0};
                writeAddr3 = {writeAddr[10:0], 3'b0};
                writeAddr2 = {writeAddr[10:0], 3'b0};
                writeAddr1 = {writeAddr[10:0], 3'b0};

                readAddr4  = {readAddr[10:0],  3'b0};
                readAddr3  = {readAddr[10:0],  3'b0};
                readAddr2  = {readAddr[10:0],  3'b0};
                readAddr1  = {readAddr[10:0],  3'b0};

                writeData4 = {10'b0, writeData[31:24]};
                writeData3 = {10'b0, writeData[23:16]};
                writeData2 = {10'b0, writeData[15:8]};
                writeData1 = {10'b0, writeData[7:0]};

                wen_a4 = {1'b0, wen};
                wen_a3 = {1'b0, wen};
                wen_a2 = {1'b0, wen};
                wen_a1 = {1'b0, wen};
                readData = {readData4[7:0],readData3[7:0],readData2[7:0],readData1[7:0]};
            end
            2560: begin
                width4 = 3'b011;
                width3 = 3'b011;
                width2 = 3'b011;
                width1 = 3'b011;
                width0 = 3'b101;

                writeAddr4 = {writeAddr[10:0], 3'b0};
                writeAddr3 = {writeAddr[10:0], 3'b0};
                writeAddr2 = {writeAddr[10:0], 3'b0};
                writeAddr1 = {writeAddr[10:0], 3'b0};
                writeAddr0 = {writeAddr[8:0], 5'b0};

                readAddr4  = {readAddr[10:0],  3'b0};
                readAddr3  = {readAddr[10:0],  3'b0};
                readAddr2  = {readAddr[10:0],  3'b0};
                readAddr1  = {readAddr[10:0],  3'b0};
                readAddr0  = {readAddr[8:0],  5'b0};

                writeData4 = {10'b0, writeData[31:24]};
                writeData3 = {10'b0, writeData[23:16]};
                writeData2 = {10'b0, writeData[15:8]};
                writeData1 = {10'b0, writeData[7:0]};
                writeData0 = {1'b0, writeData[31:24], 1'b0, writeData[23:16], 1'b0, writeData[15:8], 1'b0, writeData[7:0]};

                case (writeAddr[11:9])
                    3'b000 , 3'b001, 3'b010, 3'b011 : begin
                        wen_a4 = {1'b0, wen};
                        wen_a3 = {1'b0, wen};
                        wen_a2 = {1'b0, wen};
                        wen_a1 = {1'b0, wen};
                        wen_a0 = {1'b0, 1'b0};
                        wen_b0 = {1'b0, 1'b0};
                    end
                    3'b100 : begin
                        wen_a4 = {1'b0, 1'b0};
                        wen_a3 = {1'b0, 1'b0};
                        wen_a2 = {1'b0, 1'b0};
                        wen_a1 = {1'b0, 1'b0};
                        wen_a0 = {wen,  wen};
                        wen_b0 = {wen,  wen};
                    end
                    default: begin
                        wen_a4 = {1'b0, 1'b0};
                        wen_a3 = {1'b0, 1'b0};
                        wen_a2 = {1'b0, 1'b0};
                        wen_a1 = {1'b0, 1'b0};
                        wen_a0 = {1'b0, 1'b0};
                        wen_b0 = {1'b0, 1'b0};
                    end
                endcase
                case (ckRdAddr[11:9])
                    3'b000 , 3'b001, 3'b010, 3'b011 : begin
                        readData = {readData4[7:0],readData3[7:0],readData2[7:0],readData1[7:0]};
                    end
                    3'b100 : begin
                        readData = {readData0[34:27],readData0[25:18],readData0[16:9],readData0[7:0]};
                    end
                    default : begin
                        readData = 32'b0;
                    end
                endcase
            end
            3072: begin
                width6 = 3'b011;
                width5 = 3'b011;
                width4 = 3'b011;
                width3 = 3'b011;
                width2 = 3'b100;
                width1 = 3'b100;

                writeAddr6 = {writeAddr[10:0], 3'b0};
                writeAddr5 = {writeAddr[10:0], 3'b0};
                writeAddr4 = {writeAddr[10:0], 3'b0};
                writeAddr3 = {writeAddr[10:0], 3'b0};
                writeAddr2 = {writeAddr[9:0], 4'b0};
                writeAddr1 = {writeAddr[9:0], 4'b0};

                readAddr6  = {readAddr[10:0],  3'b0};
                readAddr5  = {readAddr[10:0],  3'b0};
                readAddr4  = {readAddr[10:0],  3'b0};
                readAddr3  = {readAddr[10:0],  3'b0};
                readAddr2  = {readAddr[9:0],  4'b0};
                readAddr1  = {readAddr[9:0],  4'b0};

                writeData6 = {10'b0, writeData[31:24]};
                writeData5 = {10'b0, writeData[23:16]};
                writeData4 = {10'b0, writeData[15:8]};
                writeData3 = {10'b0, writeData[7:0]};
                writeData2 = {1'b0, writeData[31:24], 1'b0, writeData[23:16]};
                writeData1 = {1'b0, writeData[15:8], 1'b0, writeData[7:0]};

                case (writeAddr[11:10])
                    2'b00, 2'b01 : begin
                        wen_a6 = {1'b0, wen};
                        wen_a5 = {1'b0, wen};
                        wen_a4 = {1'b0, wen};
                        wen_a3 = {1'b0, wen};
                        wen_a2 = {1'b0, 1'b0};
                        wen_a1 = {1'b0, 1'b0};
                    end
                    2'b10 : begin
                        wen_a6 = {1'b0, 1'b0};
                        wen_a5 = {1'b0, 1'b0};
                        wen_a4 = {1'b0, 1'b0};
                        wen_a3 = {1'b0, 1'b0};
                        wen_a2 = {wen, wen};
                        wen_a1 = {wen, wen};
                    end
                    2'b11 : begin
                        wen_a6 = {1'b0, 1'b0};
                        wen_a5 = {1'b0, 1'b0};
                        wen_a4 = {1'b0, 1'b0};
                        wen_a3 = {1'b0, 1'b0};
                        wen_a2 = {1'b0, 1'b0};
                        wen_a1 = {1'b0, 1'b0};
                    end
                endcase
                case (ckRdAddr[11:10])
                    2'b00, 2'b01 : begin
                        readData = {readData6[7:0],readData5[7:0],readData4[7:0],readData3[7:0]};
                    end
                    2'b10 : begin
                        readData = {readData2[16:9],readData2[7:0],readData1[16:9],readData1[7:0]};
                    end
                    2'b11 : begin
                        readData = 32'b0;
                    end
                endcase
            end
            3584: begin
                width6 = 3'b011;
                width5 = 3'b011;
                width4 = 3'b011;
                width3 = 3'b011;
                width2 = 3'b100;
                width1 = 3'b100;
                width0 = 3'b101;

                writeAddr6 = {writeAddr[10:0], 3'b0};
                writeAddr5 = {writeAddr[10:0], 3'b0};
                writeAddr4 = {writeAddr[10:0], 3'b0};
                writeAddr3 = {writeAddr[10:0], 3'b0};
                writeAddr2 = {writeAddr[9:0], 4'b0};
                writeAddr1 = {writeAddr[9:0], 4'b0};
                writeAddr0 = {writeAddr[8:0], 5'b0};

                readAddr6  = {readAddr[10:0],  3'b0};
                readAddr5  = {readAddr[10:0],  3'b0};
                readAddr4  = {readAddr[10:0],  3'b0};
                readAddr3  = {readAddr[10:0],  3'b0};
                readAddr2  = {readAddr[9:0],  4'b0};
                readAddr1  = {readAddr[9:0],  4'b0};
                readAddr0  = {readAddr[8:0],  5'b0};

                writeData6 = {10'b0, writeData[31:24]};
                writeData5 = {10'b0, writeData[23:16]};
                writeData4 = {10'b0, writeData[15:8]};
                writeData3 = {10'b0, writeData[7:0]};
                writeData2 = {1'b0, writeData[31:24], 1'b0, writeData[23:16]};
                writeData1 = {1'b0, writeData[15:8], 1'b0, writeData[7:0]};
                writeData0 = {1'b0, writeData[31:24], 1'b0, writeData[23:16], 1'b0, writeData[15:8], 1'b0, writeData[7:0]};

                case (writeAddr[11:9])
                    3'b000, 3'b001, 3'b010, 3'b011 : begin
                        wen_a6 = {1'b0, wen};
                        wen_a5 = {1'b0, wen};
                        wen_a4 = {1'b0, wen};
                        wen_a3 = {1'b0, wen};
                        wen_a2 = {1'b0, 1'b0};
                        wen_a1 = {1'b0, 1'b0};
                        wen_a0 = {1'b0, 1'b0};
                        wen_b0 = {1'b0, 1'b0};
                    end
                    3'b100, 3'b101 : begin
                        wen_a6 = {1'b0, 1'b0};
                        wen_a5 = {1'b0, 1'b0};
                        wen_a4 = {1'b0, 1'b0};
                        wen_a3 = {1'b0, 1'b0};
                        wen_a2 = {wen, wen};
                        wen_a1 = {wen, wen};
                        wen_a0 = {1'b0, 1'b0};
                        wen_b0 = {1'b0, 1'b0};
                    end
                    3'b110 : begin
                        wen_a6 = {1'b0, 1'b0};
                        wen_a5 = {1'b0, 1'b0};
                        wen_a4 = {1'b0, 1'b0};
                        wen_a3 = {1'b0, 1'b0};
                        wen_a2 = {1'b0, 1'b0};
                        wen_a1 = {1'b0, 1'b0};
                        wen_a0 = {wen, wen};
                        wen_b0 = {wen, wen};
                    end
                    3'b111 : begin
                        wen_a6 = {1'b0, 1'b0};
                        wen_a5 = {1'b0, 1'b0};
                        wen_a4 = {1'b0, 1'b0};
                        wen_a3 = {1'b0, 1'b0};
                        wen_a2 = {1'b0, 1'b0};
                        wen_a1 = {1'b0, 1'b0};
                        wen_a0 = {1'b0, 1'b0};
                        wen_b0 = {1'b0, 1'b0};
                    end
                endcase
                case (ckRdAddr[11:9])
                    3'b000, 3'b001, 3'b010, 3'b011 : begin
                        readData = {readData6[7:0],readData5[7:0],readData4[7:0],readData3[7:0]};
                    end
                    3'b100, 3'b101 : begin
                        readData = {readData2[16:9],readData2[7:0],readData1[16:9],readData1[7:0]};
                    end
                    3'b110 : begin
                        readData = {readData0[34:27],readData0[25:18],readData0[16:9],readData0[7:0]};
                    end
                    3'b111 : begin
                        readData = 32'b0;
                    end
                endcase
            end
            4096: begin
                width8 = 3'b010;
                width7 = 3'b010;
                width6 = 3'b010;
                width5 = 3'b010;
                width4 = 3'b010;
                width3 = 3'b010;
                width2 = 3'b010;
                width1 = 3'b010;

                writeAddr8 = {writeAddr[11:0], 2'b0};
                writeAddr7 = {writeAddr[11:0], 2'b0};
                writeAddr6 = {writeAddr[11:0], 2'b0};
                writeAddr5 = {writeAddr[11:0], 2'b0};
                writeAddr4 = {writeAddr[11:0], 2'b0};
                writeAddr3 = {writeAddr[11:0], 2'b0};
                writeAddr2 = {writeAddr[11:0], 2'b0};
                writeAddr1 = {writeAddr[11:0], 2'b0};

                readAddr8  = {readAddr[11:0],  2'b0};
                readAddr7  = {readAddr[11:0],  2'b0};
                readAddr6  = {readAddr[11:0],  2'b0};
                readAddr5  = {readAddr[11:0],  2'b0};
                readAddr4  = {readAddr[11:0],  2'b0};
                readAddr3  = {readAddr[11:0],  2'b0};
                readAddr2  = {readAddr[11:0],  2'b0};
                readAddr1  = {readAddr[11:0],  2'b0};

                writeData8 = {14'b0, writeData[31:28]};
                writeData7 = {14'b0, writeData[27:24]};
                writeData6 = {14'b0, writeData[23:20]};
                writeData5 = {14'b0, writeData[19:16]};
                writeData4 = {14'b0, writeData[15:12]};
                writeData3 = {14'b0, writeData[11:8]};
                writeData2 = {14'b0, writeData[7:4]};
                writeData1 = {14'b0, writeData[3:0]};

                wen_a8 = {1'b0, wen};
                wen_a7 = {1'b0, wen};
                wen_a6 = {1'b0, wen};
                wen_a5 = {1'b0, wen};
                wen_a4 = {1'b0, wen};
                wen_a3 = {1'b0, wen};
                wen_a2 = {1'b0, wen};
                wen_a1 = {1'b0, wen};

                readData = {
                                readData8[3:0],
                                readData7[3:0],
                                readData6[3:0],
                                readData5[3:0],
                                readData4[3:0],
                                readData3[3:0],
                                readData2[3:0],
                                readData1[3:0]
                };
            end
            4608: begin
                width8 = 3'b010;
                width7 = 3'b010;
                width6 = 3'b010;
                width5 = 3'b010;
                width4 = 3'b010;
                width3 = 3'b010;
                width2 = 3'b010;
                width1 = 3'b010;
                width0 = 3'b101;

                writeAddr8 = {writeAddr[11:0], 2'b0};
                writeAddr7 = {writeAddr[11:0], 2'b0};
                writeAddr6 = {writeAddr[11:0], 2'b0};
                writeAddr5 = {writeAddr[11:0], 2'b0};
                writeAddr4 = {writeAddr[11:0], 2'b0};
                writeAddr3 = {writeAddr[11:0], 2'b0};
                writeAddr2 = {writeAddr[11:0], 2'b0};
                writeAddr1 = {writeAddr[11:0], 2'b0};
                writeAddr0 = {writeAddr[8:0], 5'b0};

                readAddr8  = {readAddr[11:0],  2'b0};
                readAddr7  = {readAddr[11:0],  2'b0};
                readAddr6  = {readAddr[11:0],  2'b0};
                readAddr5  = {readAddr[11:0],  2'b0};
                readAddr4  = {readAddr[11:0],  2'b0};
                readAddr3  = {readAddr[11:0],  2'b0};
                readAddr2  = {readAddr[11:0],  2'b0};
                readAddr1  = {readAddr[11:0],  2'b0};
                readAddr0  = {readAddr[8:0],  5'b0};

                writeData8 = {14'b0, writeData[31:28]};
                writeData7 = {14'b0, writeData[27:24]};
                writeData6 = {14'b0, writeData[23:20]};
                writeData5 = {14'b0, writeData[19:16]};
                writeData4 = {14'b0, writeData[15:12]};
                writeData3 = {14'b0, writeData[11:8]};
                writeData2 = {14'b0, writeData[7:4]};
                writeData1 = {14'b0, writeData[3:0]};
                writeData0 = {1'b0, writeData[31:24], 1'b0, writeData[23:16], 1'b0, writeData[15:8], 1'b0, writeData[7:0]};

                case (writeAddr[12:9])
                    4'b0000, 4'b0001, 4'b0010, 4'b0011,
                    4'b0100, 4'b0101, 4'b0110, 4'b0111 : begin
                        wen_a8 = {1'b0, wen};
                        wen_a7 = {1'b0, wen};
                        wen_a6 = {1'b0, wen};
                        wen_a5 = {1'b0, wen};
                        wen_a4 = {1'b0, wen};
                        wen_a3 = {1'b0, wen};
                        wen_a2 = {1'b0, wen};
                        wen_a1 = {1'b0, wen};
                        wen_a0 = {1'b0, 1'b0};
                        wen_b0 = {1'b0, 1'b0};
                    end
                    4'b1000 : begin
                        wen_a8 = {1'b0, 1'b0};
                        wen_a7 = {1'b0, 1'b0};
                        wen_a6 = {1'b0, 1'b0};
                        wen_a5 = {1'b0, 1'b0};
                        wen_a4 = {1'b0, 1'b0};
                        wen_a3 = {1'b0, 1'b0};
                        wen_a2 = {1'b0, 1'b0};
                        wen_a1 = {1'b0, 1'b0};
                        wen_a0 = {wen, wen};
                        wen_b0 = {wen, wen};
                    end
                    default : begin
                        wen_a8 = {1'b0, 1'b0};
                        wen_a7 = {1'b0, 1'b0};
                        wen_a6 = {1'b0, 1'b0};
                        wen_a5 = {1'b0, 1'b0};
                        wen_a4 = {1'b0, 1'b0};
                        wen_a3 = {1'b0, 1'b0};
                        wen_a2 = {1'b0, 1'b0};
                        wen_a1 = {1'b0, 1'b0};
                        wen_a0 = {1'b0, 1'b0};
                        wen_b0 = {1'b0, 1'b0};
                    end
                endcase
                case (ckRdAddr[12:9])
                    4'b0000, 4'b0001, 4'b0010, 4'b0011,
                    4'b0100, 4'b0101, 4'b0110, 4'b0111 : begin
                        readData = {
                                        readData8[3:0],
                                        readData7[3:0],
                                        readData6[3:0],
                                        readData5[3:0],
                                        readData4[3:0],
                                        readData3[3:0],
                                        readData2[3:0],
                                        readData1[3:0]
                        };
                    end
                    4'b1000 : begin
                        readData = {readData0[34:27],readData0[25:18],readData0[16:9],readData0[7:0]};
                    end
                    default : begin
                        readData = 32'b0;
                    end
                endcase
            end
            5120: begin
                width10 = 3'b010;
                width9 = 3'b010;
                width8 = 3'b010;
                width7 = 3'b010;
                width6 = 3'b010;
                width5 = 3'b010;
                width4 = 3'b010;
                width3 = 3'b010;
                width2 = 3'b100;
                width1 = 3'b100;
                writeAddr10 = {writeAddr[11:0], 2'b0};
                writeAddr9 = {writeAddr[11:0], 2'b0};
                writeAddr8 = {writeAddr[11:0], 2'b0};
                writeAddr7 = {writeAddr[11:0], 2'b0};
                writeAddr6 = {writeAddr[11:0], 2'b0};
                writeAddr5 = {writeAddr[11:0], 2'b0};
                writeAddr4 = {writeAddr[11:0], 2'b0};
                writeAddr3 = {writeAddr[11:0], 2'b0};
                writeAddr2 = {writeAddr[9:0], 4'b0};
                writeAddr1 = {writeAddr[9:0], 4'b0};
                readAddr10  = {readAddr[11:0],  2'b0};
                readAddr9  = {readAddr[11:0],  2'b0};
                readAddr8  = {readAddr[11:0],  2'b0};
                readAddr7  = {readAddr[11:0],  2'b0};
                readAddr6  = {readAddr[11:0],  2'b0};
                readAddr5  = {readAddr[11:0],  2'b0};
                readAddr4  = {readAddr[11:0],  2'b0};
                readAddr3  = {readAddr[11:0],  2'b0};
                readAddr2  = {readAddr[9:0],  4'b0};
                readAddr1  = {readAddr[9:0],  4'b0};
                writeData10 = {14'b0, writeData[31:28]};
                writeData9 = {14'b0, writeData[27:24]};
                writeData8 = {14'b0, writeData[23:20]};
                writeData7 = {14'b0, writeData[19:16]};
                writeData6 = {14'b0, writeData[15:12]};
                writeData5 = {14'b0, writeData[11:8]};
                writeData4 = {14'b0, writeData[7:4]};
                writeData3 = {14'b0, writeData[3:0]};
                writeData2 = {1'b0, writeData[31:24], 1'b0, writeData[23:16]};
                writeData1 = {1'b0, writeData[15:8], 1'b0, writeData[7:0]};
                case (writeAddr[12:9])
                    4'b0000, 4'b0001, 4'b0010, 4'b0011,
                    4'b0100, 4'b0101, 4'b0110, 4'b0111 : begin
                        wen_a10 = {1'b0, wen};
                        wen_a9 = {1'b0, wen};
                        wen_a8 = {1'b0, wen};
                        wen_a7 = {1'b0, wen};
                        wen_a6 = {1'b0, wen};
                        wen_a5 = {1'b0, wen};
                        wen_a4 = {1'b0, wen};
                        wen_a3 = {1'b0, wen};
                        wen_a2 = {1'b0, 1'b0};
                        wen_a1 = {1'b0, 1'b0};
                    end
                    4'b1000, 4'b1001 : begin
                        wen_a10 = {1'b0, 1'b0};
                        wen_a9 = {1'b0, 1'b0};
                        wen_a8 = {1'b0, 1'b0};
                        wen_a7 = {1'b0, 1'b0};
                        wen_a6 = {1'b0, 1'b0};
                        wen_a5 = {1'b0, 1'b0};
                        wen_a4 = {1'b0, 1'b0};
                        wen_a3 = {1'b0, 1'b0};
                        wen_a2 = {wen, wen};
                        wen_a1 = {wen, wen};
                    end
                    default : begin
                        wen_a10 = {1'b0, 1'b0};
                        wen_a9 = {1'b0, 1'b0};
                        wen_a8 = {1'b0, 1'b0};
                        wen_a7 = {1'b0, 1'b0};
                        wen_a6 = {1'b0, 1'b0};
                        wen_a5 = {1'b0, 1'b0};
                        wen_a4 = {1'b0, 1'b0};
                        wen_a3 = {1'b0, 1'b0};
                        wen_a2 = {1'b0, 1'b0};
                        wen_a1 = {1'b0, 1'b0};
                    end
                endcase
                case (ckRdAddr[12:9])
                    4'b0000, 4'b0001, 4'b0010, 4'b0011,
                    4'b0100, 4'b0101, 4'b0110, 4'b0111 : begin
                        readData = {
                                        readData10[3:0],
                                        readData9[3:0],
                                        readData8[3:0],
                                        readData7[3:0],
                                        readData6[3:0],
                                        readData5[3:0],
                                        readData4[3:0],
                                        readData3[3:0]
                        };
                    end
                    4'b1000, 4'b1001 : begin
                        readData = {readData2[16:9],readData2[7:0],readData1[16:9],readData1[7:0]};
                    end
                    default : begin
                        readData = 32'b0;
                    end
                endcase
            end
            5632: begin
                width10 = 3'b010;
                width9 = 3'b010;
                width8 = 3'b010;
                width7 = 3'b010;
                width6 = 3'b010;
                width5 = 3'b010;
                width4 = 3'b010;
                width3 = 3'b010;
                width2 = 3'b100;
                width1 = 3'b100;
                width0 = 3'b101;
                writeAddr10 = {writeAddr[11:0], 2'b0};
                writeAddr9 = {writeAddr[11:0], 2'b0};
                writeAddr8 = {writeAddr[11:0], 2'b0};
                writeAddr7 = {writeAddr[11:0], 2'b0};
                writeAddr6 = {writeAddr[11:0], 2'b0};
                writeAddr5 = {writeAddr[11:0], 2'b0};
                writeAddr4 = {writeAddr[11:0], 2'b0};
                writeAddr3 = {writeAddr[11:0], 2'b0};
                writeAddr2 = {writeAddr[9:0], 4'b0};
                writeAddr1 = {writeAddr[9:0], 4'b0};
                writeAddr0 = {writeAddr[8:0], 5'b0};
                readAddr10  = {readAddr[11:0],  2'b0};
                readAddr9  = {readAddr[11:0],  2'b0};
                readAddr8  = {readAddr[11:0],  2'b0};
                readAddr7  = {readAddr[11:0],  2'b0};
                readAddr6  = {readAddr[11:0],  2'b0};
                readAddr5  = {readAddr[11:0],  2'b0};
                readAddr4  = {readAddr[11:0],  2'b0};
                readAddr3  = {readAddr[11:0],  2'b0};
                readAddr2  = {readAddr[9:0],  4'b0};
                readAddr1  = {readAddr[9:0],  4'b0};
                readAddr0  = {readAddr[8:0],  5'b0};
                writeData10 = {14'b0, writeData[31:28]};
                writeData9 = {14'b0, writeData[27:24]};
                writeData8 = {14'b0, writeData[23:20]};
                writeData7 = {14'b0, writeData[19:16]};
                writeData6 = {14'b0, writeData[15:12]};
                writeData5 = {14'b0, writeData[11:8]};
                writeData4 = {14'b0, writeData[7:4]};
                writeData3 = {14'b0, writeData[3:0]};
                writeData2 = {1'b0, writeData[31:24], 1'b0, writeData[23:16]};
                writeData1 = {1'b0, writeData[15:8], 1'b0, writeData[7:0]};
                writeData0 = {1'b0, writeData[31:24], 1'b0, writeData[23:16], 1'b0, writeData[15:8], 1'b0, writeData[7:0]};
                case (writeAddr[12:9])
                    4'b0000, 4'b0001, 4'b0010, 4'b0011,
                    4'b0100, 4'b0101, 4'b0110, 4'b0111 : begin
                        wen_a10 = {1'b0, wen};
                        wen_a9 = {1'b0, wen};
                        wen_a8 = {1'b0, wen};
                        wen_a7 = {1'b0, wen};
                        wen_a6 = {1'b0, wen};
                        wen_a5 = {1'b0, wen};
                        wen_a4 = {1'b0, wen};
                        wen_a3 = {1'b0, wen};
                        wen_a2 = {1'b0, 1'b0};
                        wen_a1 = {1'b0, 1'b0};
                        wen_a0 = {1'b0, 1'b0};
                        wen_b0 = {1'b0, 1'b0};
                    end
                    4'b1000, 4'b1001 : begin
                        wen_a10 = {1'b0, 1'b0};
                        wen_a9 = {1'b0, 1'b0};
                        wen_a8 = {1'b0, 1'b0};
                        wen_a7 = {1'b0, 1'b0};
                        wen_a6 = {1'b0, 1'b0};
                        wen_a5 = {1'b0, 1'b0};
                        wen_a4 = {1'b0, 1'b0};
                        wen_a3 = {1'b0, 1'b0};
                        wen_a2 = {wen, wen};
                        wen_a1 = {wen, wen};
                        wen_a0 = {1'b0, 1'b0};
                        wen_b0 = {1'b0, 1'b0};
                    end
                    4'b1010 : begin
                        wen_a10 = {1'b0, 1'b0};
                        wen_a9 = {1'b0, 1'b0};
                        wen_a8 = {1'b0, 1'b0};
                        wen_a7 = {1'b0, 1'b0};
                        wen_a6 = {1'b0, 1'b0};
                        wen_a5 = {1'b0, 1'b0};
                        wen_a4 = {1'b0, 1'b0};
                        wen_a3 = {1'b0, 1'b0};
                        wen_a0 = {wen,  wen};
                        wen_b0 = {wen,  wen};
                    end
                    default : begin
                        wen_a10 = {1'b0, 1'b0};
                        wen_a9 = {1'b0, 1'b0};
                        wen_a8 = {1'b0, 1'b0};
                        wen_a7 = {1'b0, 1'b0};
                        wen_a6 = {1'b0, 1'b0};
                        wen_a5 = {1'b0, 1'b0};
                        wen_a4 = {1'b0, 1'b0};
                        wen_a3 = {1'b0, 1'b0};
                        wen_a2 = {1'b0, 1'b0};
                        wen_a1 = {1'b0, 1'b0};
                        wen_a0 = {1'b0, 1'b0};
                        wen_b0 = {1'b0, 1'b0};
                    end
                endcase
                case (ckRdAddr[12:9])
                    4'b0000, 4'b0001, 4'b0010, 4'b0011,
                    4'b0100, 4'b0101, 4'b0110, 4'b0111 : begin
                        readData = {
                                        readData10[3:0],
                                        readData9[3:0],
                                        readData8[3:0],
                                        readData7[3:0],
                                        readData6[3:0],
                                        readData5[3:0],
                                        readData4[3:0],
                                        readData3[3:0]
                        };
                    end
                    4'b1000, 4'b1001 : begin
                        readData = {readData2[16:9],readData2[7:0],readData1[16:9],readData1[7:0]};
                    end
                    4'b1010 : begin
                        readData = {readData0[34:27],readData0[25:18],readData0[16:9],readData0[7:0]};
                    end
                    default : begin
                        readData = 32'b0;
                    end
                endcase
            end
            6144: begin
                width12 = 3'b010;
                width11 = 3'b010;
                width10 = 3'b010;
                width9 = 3'b010;
                width8 = 3'b010;
                width7 = 3'b010;
                width6 = 3'b010;
                width5 = 3'b010;
                width4 = 3'b011;
                width3 = 3'b011;
                width2 = 3'b011;
                width1 = 3'b011;
                writeAddr12 = {writeAddr[11:0], 2'b0};
                writeAddr11 = {writeAddr[11:0], 2'b0};
                writeAddr10 = {writeAddr[11:0], 2'b0};
                writeAddr9 = {writeAddr[11:0], 2'b0};
                writeAddr8 = {writeAddr[11:0], 2'b0};
                writeAddr7 = {writeAddr[11:0], 2'b0};
                writeAddr6 = {writeAddr[11:0], 2'b0};
                writeAddr5 = {writeAddr[11:0], 2'b0};
                writeAddr4 = {writeAddr[10:0], 3'b0};
                writeAddr3 = {writeAddr[10:0], 3'b0};
                writeAddr2 = {writeAddr[10:0], 3'b0};
                writeAddr1 = {writeAddr[10:0], 3'b0};
                readAddr12  = {readAddr[11:0],  2'b0};
                readAddr11  = {readAddr[11:0],  2'b0};
                readAddr10  = {readAddr[11:0],  2'b0};
                readAddr9  = {readAddr[11:0],  2'b0};
                readAddr8  = {readAddr[11:0],  2'b0};
                readAddr7  = {readAddr[11:0],  2'b0};
                readAddr6  = {readAddr[11:0],  2'b0};
                readAddr5  = {readAddr[11:0],  2'b0};
                readAddr4  = {readAddr[10:0],  3'b0};
                readAddr3  = {readAddr[10:0],  3'b0};
                readAddr2  = {readAddr[10:0],  3'b0};
                readAddr1  = {readAddr[10:0],  3'b0};
                writeData12 = {14'b0, writeData[31:28]};
                writeData11 = {14'b0, writeData[27:24]};
                writeData10 = {14'b0, writeData[23:20]};
                writeData9 = {14'b0, writeData[19:16]};
                writeData8 = {14'b0, writeData[15:12]};
                writeData7 = {14'b0, writeData[11:8]};
                writeData6 = {14'b0, writeData[7:4]};
                writeData5 = {14'b0, writeData[3:0]};
                writeData4 = {10'b0, writeData[31:24]};
                writeData3 = {10'b0, writeData[23:16]};
                writeData2 = {10'b0, writeData[15:8]};
                writeData1 = {10'b0, writeData[7:0]};
                case (writeAddr[12:9])
                    4'b0000, 4'b0001, 4'b0010, 4'b0011,
                    4'b0100, 4'b0101, 4'b0110, 4'b0111 : begin
                        wen_a12 = {1'b0, wen};
                        wen_a11 = {1'b0, wen};
                        wen_a10 = {1'b0, wen};
                        wen_a9 = {1'b0, wen};
                        wen_a8 = {1'b0, wen};
                        wen_a7 = {1'b0, wen};
                        wen_a6 = {1'b0, wen};
                        wen_a5 = {1'b0, wen};
                        wen_a4 = {1'b0, 1'b0};
                        wen_a3 = {1'b0, 1'b0};
                        wen_a2 = {1'b0, 1'b0};
                        wen_a1 = {1'b0, 1'b0};
                    end
                    4'b1000, 4'b1001, 4'b1010, 4'b1011 : begin
                        wen_a12 = {1'b0, 1'b0};
                        wen_a11 = {1'b0, 1'b0};
                        wen_a10 = {1'b0, 1'b0};
                        wen_a9 = {1'b0, 1'b0};
                        wen_a8 = {1'b0, 1'b0};
                        wen_a7 = {1'b0, 1'b0};
                        wen_a6 = {1'b0, 1'b0};
                        wen_a5 = {1'b0, 1'b0};
                        wen_a4 = {1'b0, wen};
                        wen_a3 = {1'b0, wen};
                        wen_a2 = {1'b0, wen};
                        wen_a1 = {1'b0, wen};
                    end
                    default : begin
                        wen_a12 = {1'b0, 1'b0};
                        wen_a11 = {1'b0, 1'b0};
                        wen_a10 = {1'b0, 1'b0};
                        wen_a9 = {1'b0, 1'b0};
                        wen_a8 = {1'b0, 1'b0};
                        wen_a7 = {1'b0, 1'b0};
                        wen_a6 = {1'b0, 1'b0};
                        wen_a5 = {1'b0, 1'b0};
                        wen_a4 = {1'b0, 1'b0};
                        wen_a3 = {1'b0, 1'b0};
                        wen_a2 = {1'b0, 1'b0};
                        wen_a1 = {1'b0, 1'b0};
                    end
                endcase
                case (ckRdAddr[12:9])
                    4'b0000, 4'b0001, 4'b0010, 4'b0011,
                    4'b0100, 4'b0101, 4'b0110, 4'b0111 : begin
                        readData = {
                                        readData12[3:0],
                                        readData11[3:0],
                                        readData10[3:0],
                                        readData9[3:0],
                                        readData8[3:0],
                                        readData7[3:0],
                                        readData6[3:0],
                                        readData5[3:0]
                        };
                    end
                    4'b1000, 4'b1001, 4'b1010, 4'b1011 : begin
                        readData = {readData4[7:0],readData3[7:0],readData2[7:0],readData1[7:0]};
                    end
                    default : begin
                        readData = 32'b0;
                    end
                endcase
            end
            6656: begin
                width12 = 3'b010;
                width11 = 3'b010;
                width10 = 3'b010;
                width9 = 3'b010;
                width8 = 3'b010;
                width7 = 3'b010;
                width6 = 3'b010;
                width5 = 3'b010;
                width4 = 3'b011;
                width3 = 3'b011;
                width2 = 3'b011;
                width1 = 3'b011;
                width0 = 3'b101;
                writeAddr12 = {writeAddr[11:0], 2'b0};
                writeAddr11 = {writeAddr[11:0], 2'b0};
                writeAddr10 = {writeAddr[11:0], 2'b0};
                writeAddr9 = {writeAddr[11:0], 2'b0};
                writeAddr8 = {writeAddr[11:0], 2'b0};
                writeAddr7 = {writeAddr[11:0], 2'b0};
                writeAddr6 = {writeAddr[11:0], 2'b0};
                writeAddr5 = {writeAddr[11:0], 2'b0};
                writeAddr4 = {writeAddr[10:0], 3'b0};
                writeAddr3 = {writeAddr[10:0], 3'b0};
                writeAddr2 = {writeAddr[10:0], 3'b0};
                writeAddr1 = {writeAddr[10:0], 3'b0};
                writeAddr0 = {writeAddr[8:0], 5'b0};
                readAddr12  = {readAddr[11:0],  2'b0};
                readAddr11  = {readAddr[11:0],  2'b0};
                readAddr10  = {readAddr[11:0],  2'b0};
                readAddr9  = {readAddr[11:0],  2'b0};
                readAddr8  = {readAddr[11:0],  2'b0};
                readAddr7  = {readAddr[11:0],  2'b0};
                readAddr6  = {readAddr[11:0],  2'b0};
                readAddr5  = {readAddr[11:0],  2'b0};
                readAddr4  = {readAddr[10:0],  3'b0};
                readAddr3  = {readAddr[10:0],  3'b0};
                readAddr2  = {readAddr[10:0],  3'b0};
                readAddr1  = {readAddr[10:0],  3'b0};
                readAddr0  = {readAddr[8:0],  5'b0};
                writeData12 = {14'b0, writeData[31:28]};
                writeData11 = {14'b0, writeData[27:24]};
                writeData10 = {14'b0, writeData[23:20]};
                writeData9 = {14'b0, writeData[19:16]};
                writeData8 = {14'b0, writeData[15:12]};
                writeData7 = {14'b0, writeData[11:8]};
                writeData6 = {14'b0, writeData[7:4]};
                writeData5 = {14'b0, writeData[3:0]};
                writeData4 = {10'b0, writeData[31:24]};
                writeData3 = {10'b0, writeData[23:16]};
                writeData2 = {10'b0, writeData[15:8]};
                writeData1 = {10'b0, writeData[7:0]};
                writeData0 = {1'b0, writeData[31:24], 1'b0, writeData[23:16], 1'b0, writeData[15:8], 1'b0, writeData[7:0]};
                case (writeAddr[12:9])
                    4'b0000, 4'b0001, 4'b0010, 4'b0011,
                    4'b0100, 4'b0101, 4'b0110, 4'b0111 : begin
                        wen_a12 = {1'b0, wen};
                        wen_a11 = {1'b0, wen};
                        wen_a10 = {1'b0, wen};
                        wen_a9 = {1'b0, wen};
                        wen_a8 = {1'b0, wen};
                        wen_a7 = {1'b0, wen};
                        wen_a6 = {1'b0, wen};
                        wen_a5 = {1'b0, wen};
                        wen_a4 = {1'b0, 1'b0};
                        wen_a3 = {1'b0, 1'b0};
                        wen_a2 = {1'b0, 1'b0};
                        wen_a1 = {1'b0, 1'b0};
                        wen_a0 = {1'b0, 1'b0};
                        wen_b0 = {1'b0, 1'b0};
                    end
                    4'b1000, 4'b1001, 4'b1010, 4'b1011 : begin
                        wen_a12 = {1'b0, 1'b0};
                        wen_a11 = {1'b0, 1'b0};
                        wen_a10 = {1'b0, 1'b0};
                        wen_a9 = {1'b0, 1'b0};
                        wen_a8 = {1'b0, 1'b0};
                        wen_a7 = {1'b0, 1'b0};
                        wen_a6 = {1'b0, 1'b0};
                        wen_a5 = {1'b0, 1'b0};
                        wen_a4 = {1'b0, wen};
                        wen_a3 = {1'b0, wen};
                        wen_a2 = {1'b0, wen};
                        wen_a1 = {1'b0, wen};
                        wen_a0 = {1'b0, 1'b0};
                        wen_b0 = {1'b0, 1'b0};
                    end
                    4'b1100 : begin
                        wen_a12 = {1'b0, 1'b0};
                        wen_a11 = {1'b0, 1'b0};
                        wen_a10 = {1'b0, 1'b0};
                        wen_a9 = {1'b0, 1'b0};
                        wen_a8 = {1'b0, 1'b0};
                        wen_a7 = {1'b0, 1'b0};
                        wen_a6 = {1'b0, 1'b0};
                        wen_a5 = {1'b0, 1'b0};
                        wen_a4 = {1'b0, 1'b0};
                        wen_a3 = {1'b0, 1'b0};
                        wen_a2 = {1'b0, 1'b0};
                        wen_a1 = {1'b0, 1'b0};
                        wen_a0 = {wen, wen};
                        wen_b0 = {wen, wen};
                    end
                    default : begin
                        wen_a12 = {1'b0, 1'b0};
                        wen_a11 = {1'b0, 1'b0};
                        wen_a10 = {1'b0, 1'b0};
                        wen_a9 = {1'b0, 1'b0};
                        wen_a8 = {1'b0, 1'b0};
                        wen_a7 = {1'b0, 1'b0};
                        wen_a6 = {1'b0, 1'b0};
                        wen_a5 = {1'b0, 1'b0};
                        wen_a4 = {1'b0, 1'b0};
                        wen_a3 = {1'b0, 1'b0};
                        wen_a2 = {1'b0, 1'b0};
                        wen_a1 = {1'b0, 1'b0};
                        wen_a0 = {1'b0, 1'b0};
                        wen_b0 = {1'b0, 1'b0};
                    end
                endcase
                case (ckRdAddr[12:9])
                    4'b0000, 4'b0001, 4'b0010, 4'b0011,
                    4'b0100, 4'b0101, 4'b0110, 4'b0111 : begin
                        readData = {
                                        readData12[3:0],
                                        readData11[3:0],
                                        readData10[3:0],
                                        readData9[3:0],
                                        readData8[3:0],
                                        readData7[3:0],
                                        readData6[3:0],
                                        readData5[3:0]
                        };
                    end
                    4'b1000, 4'b1001, 4'b1010, 4'b1011 : begin
                        readData = {readData4[7:0],readData3[7:0],readData2[7:0],readData1[7:0]};
                    end
                    4'b1100 : begin
                        readData = {readData0[34:27],readData0[25:18],readData0[16:9],readData0[7:0]};
                    end
                    default : begin
                        readData = 32'b0;
                    end
                endcase
            end
            7168: begin
                width14 = 3'b010;
                width13 = 3'b010;
                width12 = 3'b010;
                width11 = 3'b010;
                width10 = 3'b010;
                width9 = 3'b010;
                width8 = 3'b010;
                width7 = 3'b010;
                width6 = 3'b011;
                width5 = 3'b011;
                width4 = 3'b011;
                width3 = 3'b011;
                width2 = 3'b100;
                width1 = 3'b100;

                writeAddr14 = {writeAddr[11:0], 2'b0};
                writeAddr13 = {writeAddr[11:0], 2'b0};
                writeAddr12 = {writeAddr[11:0], 2'b0};
                writeAddr11 = {writeAddr[11:0], 2'b0};
                writeAddr10 = {writeAddr[11:0], 2'b0};
                writeAddr9 = {writeAddr[11:0], 2'b0};
                writeAddr8 = {writeAddr[11:0], 2'b0};
                writeAddr7 = {writeAddr[11:0], 2'b0};
                writeAddr6 = {writeAddr[10:0], 3'b0};
                writeAddr5 = {writeAddr[10:0], 3'b0};
                writeAddr4 = {writeAddr[10:0], 3'b0};
                writeAddr3 = {writeAddr[10:0], 3'b0};
                writeAddr2 = {writeAddr[9:0], 4'b0};
                writeAddr1 = {writeAddr[9:0], 4'b0};

                readAddr14  = {readAddr[11:0],  2'b0};
                readAddr13  = {readAddr[11:0],  2'b0};
                readAddr12  = {readAddr[11:0],  2'b0};
                readAddr11  = {readAddr[11:0],  2'b0};
                readAddr10  = {readAddr[11:0],  2'b0};
                readAddr9  = {readAddr[11:0],  2'b0};
                readAddr8  = {readAddr[11:0],  2'b0};
                readAddr7  = {readAddr[11:0],  2'b0};
                readAddr6  = {readAddr[10:0],  3'b0};
                readAddr5  = {readAddr[10:0],  3'b0};
                readAddr4  = {readAddr[10:0],  3'b0};
                readAddr3  = {readAddr[10:0],  3'b0};
                readAddr2  = {readAddr[9:0],  4'b0};
                readAddr1  = {readAddr[9:0],  4'b0};

                writeData14 = {14'b0, writeData[31:28]};
                writeData13 = {14'b0, writeData[27:24]};
                writeData12 = {14'b0, writeData[23:20]};
                writeData11 = {14'b0, writeData[19:16]};
                writeData10 = {14'b0, writeData[15:12]};
                writeData9 = {14'b0, writeData[11:8]};
                writeData8 = {14'b0, writeData[7:4]};
                writeData7 = {14'b0, writeData[3:0]};
                writeData6 = {10'b0, writeData[31:24]};
                writeData5 = {10'b0, writeData[23:16]};
                writeData4 = {10'b0, writeData[15:8]};
                writeData3 = {10'b0, writeData[7:0]};
                writeData2 = {1'b0, writeData[31:24], 1'b0, writeData[23:16]};
                writeData1 = {1'b0, writeData[15:8], 1'b0, writeData[7:0]};

                case (writeAddr[12:9])
                    4'b0000, 4'b0001, 4'b0010, 4'b0011,
                    4'b0100, 4'b0101, 4'b0110, 4'b0111 : begin
                        wen_a14 = {1'b0, wen};
                        wen_a13 = {1'b0, wen};
                        wen_a12 = {1'b0, wen};
                        wen_a11 = {1'b0, wen};
                        wen_a10 = {1'b0, wen};
                        wen_a9 = {1'b0, wen};
                        wen_a8 = {1'b0, wen};
                        wen_a7 = {1'b0, wen};
                        wen_a6 = {1'b0, 1'b0};
                        wen_a5 = {1'b0, 1'b0};
                        wen_a4 = {1'b0, 1'b0};
                        wen_a3 = {1'b0, 1'b0};
                        wen_a2 = {1'b0, 1'b0};
                        wen_a1 = {1'b0, 1'b0};
                    end
                    4'b1000, 4'b1001, 4'b1010, 4'b1011 : begin
                        wen_a14 = {1'b0, 1'b0};
                        wen_a13 = {1'b0, 1'b0};
                        wen_a12 = {1'b0, 1'b0};
                        wen_a11 = {1'b0, 1'b0};
                        wen_a10 = {1'b0, 1'b0};
                        wen_a9 = {1'b0, 1'b0};
                        wen_a8 = {1'b0, 1'b0};
                        wen_a7 = {1'b0, 1'b0};
                        wen_a6 = {1'b0, wen};
                        wen_a5 = {1'b0, wen};
                        wen_a4 = {1'b0, wen};
                        wen_a3 = {1'b0, wen};
                        wen_a2 = {1'b0, 1'b0};
                        wen_a1 = {1'b0, 1'b0};
                    end
                    4'b1100, 4'b1101 : begin
                        wen_a14 = {1'b0, 1'b0};
                        wen_a13 = {1'b0, 1'b0};
                        wen_a12 = {1'b0, 1'b0};
                        wen_a11 = {1'b0, 1'b0};
                        wen_a10 = {1'b0, 1'b0};
                        wen_a9 = {1'b0, 1'b0};
                        wen_a8 = {1'b0, 1'b0};
                        wen_a7 = {1'b0, 1'b0};
                        wen_a6 = {1'b0, 1'b0};
                        wen_a5 = {1'b0, 1'b0};
                        wen_a4 = {1'b0, 1'b0};
                        wen_a3 = {1'b0, 1'b0};
                        wen_a2 = {wen, wen};
                        wen_a1 = {wen, wen};
                    end
                    default : begin
                        wen_a14 = {1'b0, 1'b0};
                        wen_a13 = {1'b0, 1'b0};
                        wen_a12 = {1'b0, 1'b0};
                        wen_a11 = {1'b0, 1'b0};
                        wen_a10 = {1'b0, 1'b0};
                        wen_a9 = {1'b0, 1'b0};
                        wen_a8 = {1'b0, 1'b0};
                        wen_a7 = {1'b0, 1'b0};
                        wen_a6 = {1'b0, 1'b0};
                        wen_a5 = {1'b0, 1'b0};
                        wen_a4 = {1'b0, 1'b0};
                        wen_a3 = {1'b0, 1'b0};
                        wen_a2 = {1'b0, 1'b0};
                        wen_a1 = {1'b0, 1'b0};
                    end
                endcase
                case (ckRdAddr[12:9])
                    4'b0000, 4'b0001, 4'b0010, 4'b0011,
                    4'b0100, 4'b0101, 4'b0110, 4'b0111 : begin
                        readData = {
                                        readData14[3:0],
                                        readData13[3:0],
                                        readData12[3:0],
                                        readData11[3:0],
                                        readData10[3:0],
                                        readData9[3:0],
                                        readData8[3:0],
                                        readData7[3:0]
                        };
                    end
                    4'b1000, 4'b1001, 4'b1010, 4'b1011 : begin
                        readData = {readData6[7:0],readData5[7:0],readData4[7:0],readData3[7:0]};
                    end
                    4'b1100, 4'b1101 : begin
                        readData = {readData2[16:9],readData2[7:0],readData1[16:9],readData1[7:0]};
                    end
                    default : begin
                        readData = 32'b0;
                    end
                endcase
            end
            7680: begin
                width14 = 3'b010;
                width13 = 3'b010;
                width12 = 3'b010;
                width11 = 3'b010;
                width10 = 3'b010;
                width9 = 3'b010;
                width8 = 3'b010;
                width7 = 3'b010;
                width6 = 3'b011;
                width5 = 3'b011;
                width4 = 3'b011;
                width3 = 3'b011;
                width2 = 3'b100;
                width1 = 3'b100;
                width0 = 3'b101;

                writeAddr14 = {writeAddr[11:0], 2'b0};
                writeAddr13 = {writeAddr[11:0], 2'b0};
                writeAddr12 = {writeAddr[11:0], 2'b0};
                writeAddr11 = {writeAddr[11:0], 2'b0};
                writeAddr10 = {writeAddr[11:0], 2'b0};
                writeAddr9 = {writeAddr[11:0], 2'b0};
                writeAddr8 = {writeAddr[11:0], 2'b0};
                writeAddr7 = {writeAddr[11:0], 2'b0};
                writeAddr6 = {writeAddr[10:0], 3'b0};
                writeAddr5 = {writeAddr[10:0], 3'b0};
                writeAddr4 = {writeAddr[10:0], 3'b0};
                writeAddr3 = {writeAddr[10:0], 3'b0};
                writeAddr2 = {writeAddr[9:0], 4'b0};
                writeAddr1 = {writeAddr[9:0], 4'b0};
                writeAddr0 = {writeAddr[8:0], 5'b0};

                readAddr14  = {readAddr[11:0],  2'b0};
                readAddr13  = {readAddr[11:0],  2'b0};
                readAddr12  = {readAddr[11:0],  2'b0};
                readAddr11  = {readAddr[11:0],  2'b0};
                readAddr10  = {readAddr[11:0],  2'b0};
                readAddr9  = {readAddr[11:0],  2'b0};
                readAddr8  = {readAddr[11:0],  2'b0};
                readAddr7  = {readAddr[11:0],  2'b0};
                readAddr6  = {readAddr[10:0],  3'b0};
                readAddr5  = {readAddr[10:0],  3'b0};
                readAddr4  = {readAddr[10:0],  3'b0};
                readAddr3  = {readAddr[10:0],  3'b0};
                readAddr2  = {readAddr[9:0],  4'b0};
                readAddr1  = {readAddr[9:0],  4'b0};
                readAddr0  = {readAddr[8:0],  5'b0};

                writeData14 = {14'b0, writeData[31:28]};
                writeData13 = {14'b0, writeData[27:24]};
                writeData12 = {14'b0, writeData[23:20]};
                writeData11 = {14'b0, writeData[19:16]};
                writeData10 = {14'b0, writeData[15:12]};
                writeData9 = {14'b0, writeData[11:8]};
                writeData8 = {14'b0, writeData[7:4]};
                writeData7 = {14'b0, writeData[3:0]};
                writeData6 = {10'b0, writeData[31:24]};
                writeData5 = {10'b0, writeData[23:16]};
                writeData4 = {10'b0, writeData[15:8]};
                writeData3 = {10'b0, writeData[7:0]};
                writeData2 = {1'b0, writeData[31:24], 1'b0, writeData[23:16]};
                writeData1 = {1'b0, writeData[15:8], 1'b0, writeData[7:0]};
                writeData0 = {1'b0, writeData[31:24], 1'b0, writeData[23:16], 1'b0, writeData[15:8], 1'b0, writeData[7:0]};

                case (writeAddr[12:9])
                    4'b0000, 4'b0001, 4'b0010, 4'b0011,
                    4'b0100, 4'b0101, 4'b0110, 4'b0111 : begin
                        wen_a14 = {1'b0, wen};
                        wen_a13 = {1'b0, wen};
                        wen_a12 = {1'b0, wen};
                        wen_a11 = {1'b0, wen};
                        wen_a10 = {1'b0, wen};
                        wen_a9 = {1'b0, wen};
                        wen_a8 = {1'b0, wen};
                        wen_a7 = {1'b0, wen};
                        wen_a6 = {1'b0, 1'b0};
                        wen_a5 = {1'b0, 1'b0};
                        wen_a4 = {1'b0, 1'b0};
                        wen_a3 = {1'b0, 1'b0};
                        wen_a2 = {1'b0, 1'b0};
                        wen_a1 = {1'b0, 1'b0};
                        wen_a0 = {1'b0, 1'b0};
                        wen_b0 = {1'b0, 1'b0};
                    end
                    4'b1000, 4'b1001, 4'b1010, 4'b1011 : begin
                        wen_a14 = {1'b0, 1'b0};
                        wen_a13 = {1'b0, 1'b0};
                        wen_a12 = {1'b0, 1'b0};
                        wen_a11 = {1'b0, 1'b0};
                        wen_a10 = {1'b0, 1'b0};
                        wen_a9 = {1'b0, 1'b0};
                        wen_a8 = {1'b0, 1'b0};
                        wen_a7 = {1'b0, 1'b0};
                        wen_a6 = {1'b0, wen};
                        wen_a5 = {1'b0, wen};
                        wen_a4 = {1'b0, wen};
                        wen_a3 = {1'b0, wen};
                        wen_a2 = {1'b0, 1'b0};
                        wen_a1 = {1'b0, 1'b0};
                        wen_a0 = {1'b0, 1'b0};
                        wen_b0 = {1'b0, 1'b0};
                    end
                    4'b1100, 4'b1101 : begin
                        wen_a14 = {1'b0, 1'b0};
                        wen_a13 = {1'b0, 1'b0};
                        wen_a12 = {1'b0, 1'b0};
                        wen_a11 = {1'b0, 1'b0};
                        wen_a10 = {1'b0, 1'b0};
                        wen_a9 = {1'b0, 1'b0};
                        wen_a8 = {1'b0, 1'b0};
                        wen_a7 = {1'b0, 1'b0};
                        wen_a6 = {1'b0, 1'b0};
                        wen_a5 = {1'b0, 1'b0};
                        wen_a4 = {1'b0, 1'b0};
                        wen_a3 = {1'b0, 1'b0};
                        wen_a2 = {wen, wen};
                        wen_a1 = {wen, wen};
                        wen_a0 = {1'b0, 1'b0};
                        wen_b0 = {1'b0, 1'b0};
                    end
                    4'b1110 : begin
                        wen_a14 = {1'b0, 1'b0};
                        wen_a13 = {1'b0, 1'b0};
                        wen_a12 = {1'b0, 1'b0};
                        wen_a11 = {1'b0, 1'b0};
                        wen_a10 = {1'b0, 1'b0};
                        wen_a9 = {1'b0, 1'b0};
                        wen_a8 = {1'b0, 1'b0};
                        wen_a7 = {1'b0, 1'b0};
                        wen_a6 = {1'b0, 1'b0};
                        wen_a5 = {1'b0, 1'b0};
                        wen_a4 = {1'b0, 1'b0};
                        wen_a3 = {1'b0, 1'b0};
                        wen_a2 = {1'b0, 1'b0};
                        wen_a1 = {1'b0, 1'b0};
                        wen_a0 = {wen, wen};
                        wen_b0 = {wen, wen};
                    end
                    default : begin
                        wen_a14 = {1'b0, 1'b0};
                        wen_a13 = {1'b0, 1'b0};
                        wen_a12 = {1'b0, 1'b0};
                        wen_a11 = {1'b0, 1'b0};
                        wen_a10 = {1'b0, 1'b0};
                        wen_a9 = {1'b0, 1'b0};
                        wen_a8 = {1'b0, 1'b0};
                        wen_a7 = {1'b0, 1'b0};
                        wen_a6 = {1'b0, 1'b0};
                        wen_a5 = {1'b0, 1'b0};
                        wen_a4 = {1'b0, 1'b0};
                        wen_a3 = {1'b0, 1'b0};
                        wen_a2 = {1'b0, 1'b0};
                        wen_a1 = {1'b0, 1'b0};
                        wen_a0 = {1'b0, 1'b0};
                        wen_b0 = {1'b0, 1'b0};
                    end
                endcase
                case (ckRdAddr[12:9])
                    4'b0000, 4'b0001, 4'b0010, 4'b0011,
                    4'b0100, 4'b0101, 4'b0110, 4'b0111 : begin
                        readData = {
                                        readData14[3:0],
                                        readData13[3:0],
                                        readData12[3:0],
                                        readData11[3:0],
                                        readData10[3:0],
                                        readData9[3:0],
                                        readData8[3:0],
                                        readData7[3:0]
                        };
                    end
                    4'b1000, 4'b1001, 4'b1010, 4'b1011 : begin
                        readData = {readData6[7:0],readData5[7:0],readData4[7:0],readData3[7:0]};
                    end
                    4'b1100, 4'b1101 : begin
                        readData = {readData2[16:9],readData2[7:0],readData1[16:9],readData1[7:0]};
                    end
                    4'b1110 : begin
                        readData = {readData0[34:27],readData0[25:18],readData0[16:9],readData0[7:0]};
                    end
                    default : begin
                        readData = 32'b0;
                    end
                endcase
            end
            8192: begin
                width16 = 3'b001;
                width15 = 3'b001;
                width14 = 3'b001;
                width13 = 3'b001;
                width12 = 3'b001;
                width11 = 3'b001;
                width10 = 3'b001;
                width9 = 3'b001;
                width8 = 3'b001;
                width7 = 3'b001;
                width6 = 3'b001;
                width5 = 3'b001;
                width4 = 3'b001;
                width3 = 3'b001;
                width2 = 3'b001;
                width1 = 3'b001;

                writeAddr16 = {writeAddr[12:0], 1'b0};
                writeAddr15 = {writeAddr[12:0], 1'b0};
                writeAddr14 = {writeAddr[12:0], 1'b0};
                writeAddr13 = {writeAddr[12:0], 1'b0};
                writeAddr12 = {writeAddr[12:0], 1'b0};
                writeAddr11 = {writeAddr[12:0], 1'b0};
                writeAddr10 = {writeAddr[12:0], 1'b0};
                writeAddr9 = {writeAddr[12:0], 1'b0};
                writeAddr8 = {writeAddr[12:0], 1'b0};
                writeAddr7 = {writeAddr[12:0], 1'b0};
                writeAddr6 = {writeAddr[12:0], 1'b0};
                writeAddr5 = {writeAddr[12:0], 1'b0};
                writeAddr4 = {writeAddr[12:0], 1'b0};
                writeAddr3 = {writeAddr[12:0], 1'b0};
                writeAddr2 = {writeAddr[12:0], 1'b0};
                writeAddr1 = {writeAddr[12:0], 1'b0};

                readAddr16  = {readAddr[12:0],  1'b0};
                readAddr15  = {readAddr[12:0],  1'b0};
                readAddr14  = {readAddr[12:0],  1'b0};
                readAddr13  = {readAddr[12:0],  1'b0};
                readAddr12  = {readAddr[12:0],  1'b0};
                readAddr11  = {readAddr[12:0],  1'b0};
                readAddr10  = {readAddr[12:0],  1'b0};
                readAddr9  = {readAddr[12:0],  1'b0};
                readAddr8  = {readAddr[12:0],  1'b0};
                readAddr7  = {readAddr[12:0],  1'b0};
                readAddr6  = {readAddr[12:0],  1'b0};
                readAddr5  = {readAddr[12:0],  1'b0};
                readAddr4  = {readAddr[12:0],  1'b0};
                readAddr3  = {readAddr[12:0],  1'b0};
                readAddr2  = {readAddr[12:0],  1'b0};
                readAddr1  = {readAddr[12:0],  1'b0};

                writeData16 = {16'b0, writeData[31:30]};
                writeData15 = {16'b0, writeData[29:28]};
                writeData14 = {16'b0, writeData[27:26]};
                writeData13 = {16'b0, writeData[25:24]};
                writeData12 = {16'b0, writeData[23:22]};
                writeData11 = {16'b0, writeData[21:20]};
                writeData10 = {16'b0, writeData[19:18]};
                writeData9 = {16'b0, writeData[17:16]};
                writeData8 = {16'b0, writeData[15:14]};
                writeData7 = {16'b0, writeData[13:12]};
                writeData6 = {16'b0, writeData[11:10]};
                writeData5 = {16'b0, writeData[9:8]};
                writeData4 = {16'b0, writeData[7:6]};
                writeData3 = {16'b0, writeData[5:4]};
                writeData2 = {16'b0, writeData[3:2]};
                writeData1 = {16'b0, writeData[1:0]};

                wen_a16 = {1'b0, wen};
                wen_a15 = {1'b0, wen};
                wen_a14 = {1'b0, wen};
                wen_a13 = {1'b0, wen};
                wen_a12 = {1'b0, wen};
                wen_a11 = {1'b0, wen};
                wen_a10 = {1'b0, wen};
                wen_a9 = {1'b0, wen};
                wen_a8 = {1'b0, wen};
                wen_a7 = {1'b0, wen};
                wen_a6 = {1'b0, wen};
                wen_a5 = {1'b0, wen};
                wen_a4 = {1'b0, wen};
                wen_a3 = {1'b0, wen};
                wen_a2 = {1'b0, wen};
                wen_a1 = {1'b0, wen};

                readData = {
                                readData16[1:0],
                                readData15[1:0],
                                readData14[1:0],
                                readData13[1:0],
                                readData12[1:0],
                                readData11[1:0],
                                readData10[1:0],
                                readData9[1:0],
                                readData8[1:0],
                                readData7[1:0],
                                readData6[1:0],
                                readData5[1:0],
                                readData4[1:0],
                                readData3[1:0],
                                readData2[1:0],
                                readData1[1:0]
                };
            end
            8704: begin
                width16 = 3'b001;
                width15 = 3'b001;
                width14 = 3'b001;
                width13 = 3'b001;
                width12 = 3'b001;
                width11 = 3'b001;
                width10 = 3'b001;
                width9 = 3'b001;
                width8 = 3'b001;
                width7 = 3'b001;
                width6 = 3'b001;
                width5 = 3'b001;
                width4 = 3'b001;
                width3 = 3'b001;
                width2 = 3'b001;
                width1 = 3'b001;
                width0 = 3'b101;

                writeAddr16 = {writeAddr[12:0], 1'b0};
                writeAddr15 = {writeAddr[12:0], 1'b0};
                writeAddr14 = {writeAddr[12:0], 1'b0};
                writeAddr13 = {writeAddr[12:0], 1'b0};
                writeAddr12 = {writeAddr[12:0], 1'b0};
                writeAddr11 = {writeAddr[12:0], 1'b0};
                writeAddr10 = {writeAddr[12:0], 1'b0};
                writeAddr9 = {writeAddr[12:0], 1'b0};
                writeAddr8 = {writeAddr[12:0], 1'b0};
                writeAddr7 = {writeAddr[12:0], 1'b0};
                writeAddr6 = {writeAddr[12:0], 1'b0};
                writeAddr5 = {writeAddr[12:0], 1'b0};
                writeAddr4 = {writeAddr[12:0], 1'b0};
                writeAddr3 = {writeAddr[12:0], 1'b0};
                writeAddr2 = {writeAddr[12:0], 1'b0};
                writeAddr1 = {writeAddr[12:0], 1'b0};
                writeAddr0 = {writeAddr[8:0], 5'b0};

                readAddr16  = {readAddr[12:0],  1'b0};
                readAddr15  = {readAddr[12:0],  1'b0};
                readAddr14  = {readAddr[12:0],  1'b0};
                readAddr13  = {readAddr[12:0],  1'b0};
                readAddr12  = {readAddr[12:0],  1'b0};
                readAddr11  = {readAddr[12:0],  1'b0};
                readAddr10  = {readAddr[12:0],  1'b0};
                readAddr9  = {readAddr[12:0],  1'b0};
                readAddr8  = {readAddr[12:0],  1'b0};
                readAddr7  = {readAddr[12:0],  1'b0};
                readAddr6  = {readAddr[12:0],  1'b0};
                readAddr5  = {readAddr[12:0],  1'b0};
                readAddr4  = {readAddr[12:0],  1'b0};
                readAddr3  = {readAddr[12:0],  1'b0};
                readAddr2  = {readAddr[12:0],  1'b0};
                readAddr1  = {readAddr[12:0],  1'b0};
                readAddr0  = {readAddr[8:0],  5'b0};

                writeData16 = {16'b0, writeData[31:30]};
                writeData15 = {16'b0, writeData[29:28]};
                writeData14 = {16'b0, writeData[27:26]};
                writeData13 = {16'b0, writeData[25:24]};
                writeData12 = {16'b0, writeData[23:22]};
                writeData11 = {16'b0, writeData[21:20]};
                writeData10 = {16'b0, writeData[19:18]};
                writeData9 = {16'b0, writeData[17:16]};
                writeData8 = {16'b0, writeData[15:14]};
                writeData7 = {16'b0, writeData[13:12]};
                writeData6 = {16'b0, writeData[11:10]};
                writeData5 = {16'b0, writeData[9:8]};
                writeData4 = {16'b0, writeData[7:6]};
                writeData3 = {16'b0, writeData[5:4]};
                writeData2 = {16'b0, writeData[3:2]};
                writeData1 = {16'b0, writeData[1:0]};
                writeData0 = {1'b0, writeData[31:24], 1'b0, writeData[23:16], 1'b0, writeData[15:8], 1'b0, writeData[7:0]};

                case (writeAddr[13:9])
                    5'b00000, 5'b00001, 5'b00010, 5'b00011,
                    5'b00100, 5'b00101, 5'b00110, 5'b00111,
                    5'b01000, 5'b01001, 5'b01010, 5'b01011,
                    5'b01100, 5'b01101, 5'b01110, 5'b01111 : begin
                        wen_a16 = {1'b0, wen};
                        wen_a15 = {1'b0, wen};
                        wen_a14 = {1'b0, wen};
                        wen_a13 = {1'b0, wen};
                        wen_a12 = {1'b0, wen};
                        wen_a11 = {1'b0, wen};
                        wen_a10 = {1'b0, wen};
                        wen_a9 = {1'b0, wen};
                        wen_a8 = {1'b0, wen};
                        wen_a7 = {1'b0, wen};
                        wen_a6 = {1'b0, wen};
                        wen_a5 = {1'b0, wen};
                        wen_a4 = {1'b0, wen};
                        wen_a3 = {1'b0, wen};
                        wen_a2 = {1'b0, wen};
                        wen_a1 = {1'b0, wen};
                        wen_a0 = {1'b0, 1'b0};
                        wen_b0 = {1'b0, 1'b0};
                    end
                    5'b10000 : begin
                        wen_a16 = {1'b0, 1'b0};
                        wen_a15 = {1'b0, 1'b0};
                        wen_a14 = {1'b0, 1'b0};
                        wen_a13 = {1'b0, 1'b0};
                        wen_a12 = {1'b0, 1'b0};
                        wen_a11 = {1'b0, 1'b0};
                        wen_a10 = {1'b0, 1'b0};
                        wen_a9 = {1'b0, 1'b0};
                        wen_a8 = {1'b0, 1'b0};
                        wen_a7 = {1'b0, 1'b0};
                        wen_a6 = {1'b0, 1'b0};
                        wen_a5 = {1'b0, 1'b0};
                        wen_a4 = {1'b0, 1'b0};
                        wen_a3 = {1'b0, 1'b0};
                        wen_a2 = {1'b0, 1'b0};
                        wen_a1 = {1'b0, 1'b0};
                        wen_a0 = {wen, wen};
                        wen_b0 = {wen, wen};
                    end
                    default : begin
                        wen_a16 = {1'b0, 1'b0};
                        wen_a15 = {1'b0, 1'b0};
                        wen_a14 = {1'b0, 1'b0};
                        wen_a13 = {1'b0, 1'b0};
                        wen_a12 = {1'b0, 1'b0};
                        wen_a11 = {1'b0, 1'b0};
                        wen_a10 = {1'b0, 1'b0};
                        wen_a9 = {1'b0, 1'b0};
                        wen_a8 = {1'b0, 1'b0};
                        wen_a7 = {1'b0, 1'b0};
                        wen_a6 = {1'b0, 1'b0};
                        wen_a5 = {1'b0, 1'b0};
                        wen_a4 = {1'b0, 1'b0};
                        wen_a3 = {1'b0, 1'b0};
                        wen_a2 = {1'b0, 1'b0};
                        wen_a1 = {1'b0, 1'b0};
                        wen_a0 = {1'b0, 1'b0};
                        wen_b0 = {1'b0, 1'b0};
                    end
                endcase
                case (ckRdAddr[13:9])
                    5'b00000, 5'b00001, 5'b00010, 5'b00011,
                    5'b00100, 5'b00101, 5'b00110, 5'b00111,
                    5'b01000, 5'b01001, 5'b01010, 5'b01011,
                    5'b01100, 5'b01101, 5'b01110, 5'b01111 : begin
                        readData = {
                                        readData16[1:0],
                                        readData15[1:0],
                                        readData14[1:0],
                                        readData13[1:0],
                                        readData12[1:0],
                                        readData11[1:0],
                                        readData10[1:0],
                                        readData9[1:0],
                                        readData8[1:0],
                                        readData7[1:0],
                                        readData6[1:0],
                                        readData5[1:0],
                                        readData4[1:0],
                                        readData3[1:0],
                                        readData2[1:0],
                                        readData1[1:0]
                        };
                    end
                    5'b10000 : begin
                        readData = {readData0[34:27],readData0[25:18],readData0[16:9],readData0[7:0]};
                    end
                    default : begin
                        readData = 32'b0;
                    end
                endcase
            end
            9216: begin
                width18 = 3'b001;
                width17 = 3'b001;
                width16 = 3'b001;
                width15 = 3'b001;
                width14 = 3'b001;
                width13 = 3'b001;
                width12 = 3'b001;
                width11 = 3'b001;
                width10 = 3'b001;
                width9 = 3'b001;
                width8 = 3'b001;
                width7 = 3'b001;
                width6 = 3'b001;
                width5 = 3'b001;
                width4 = 3'b001;
                width3 = 3'b001;
                width2 = 3'b100;
                width1 = 3'b100;

                writeAddr18 = {writeAddr[12:0], 1'b0};
                writeAddr17 = {writeAddr[12:0], 1'b0};
                writeAddr16 = {writeAddr[12:0], 1'b0};
                writeAddr15 = {writeAddr[12:0], 1'b0};
                writeAddr14 = {writeAddr[12:0], 1'b0};
                writeAddr13 = {writeAddr[12:0], 1'b0};
                writeAddr12 = {writeAddr[12:0], 1'b0};
                writeAddr11 = {writeAddr[12:0], 1'b0};
                writeAddr10 = {writeAddr[12:0], 1'b0};
                writeAddr9 = {writeAddr[12:0], 1'b0};
                writeAddr8 = {writeAddr[12:0], 1'b0};
                writeAddr7 = {writeAddr[12:0], 1'b0};
                writeAddr6 = {writeAddr[12:0], 1'b0};
                writeAddr5 = {writeAddr[12:0], 1'b0};
                writeAddr4 = {writeAddr[12:0], 1'b0};
                writeAddr3 = {writeAddr[12:0], 1'b0};
                writeAddr2 = {writeAddr[9:0], 4'b0};
                writeAddr1 = {writeAddr[9:0], 4'b0};

                readAddr18  = {readAddr[12:0],  1'b0};
                readAddr17  = {readAddr[12:0],  1'b0};
                readAddr16  = {readAddr[12:0],  1'b0};
                readAddr15  = {readAddr[12:0],  1'b0};
                readAddr14  = {readAddr[12:0],  1'b0};
                readAddr13  = {readAddr[12:0],  1'b0};
                readAddr12  = {readAddr[12:0],  1'b0};
                readAddr11  = {readAddr[12:0],  1'b0};
                readAddr10  = {readAddr[12:0],  1'b0};
                readAddr9  = {readAddr[12:0],  1'b0};
                readAddr8  = {readAddr[12:0],  1'b0};
                readAddr7  = {readAddr[12:0],  1'b0};
                readAddr6  = {readAddr[12:0],  1'b0};
                readAddr5  = {readAddr[12:0],  1'b0};
                readAddr4  = {readAddr[12:0],  1'b0};
                readAddr3  = {readAddr[12:0],  1'b0};
                readAddr2  = {readAddr[9:0],  4'b0};
                readAddr1  = {readAddr[9:0],  4'b0};

                writeData18 = {16'b0, writeData[31:30]};
                writeData17 = {16'b0, writeData[29:28]};
                writeData16 = {16'b0, writeData[27:26]};
                writeData15 = {16'b0, writeData[25:24]};
                writeData14 = {16'b0, writeData[23:22]};
                writeData13 = {16'b0, writeData[21:20]};
                writeData12 = {16'b0, writeData[19:18]};
                writeData11 = {16'b0, writeData[17:16]};
                writeData10 = {16'b0, writeData[15:14]};
                writeData9 = {16'b0, writeData[13:12]};
                writeData8 = {16'b0, writeData[11:10]};
                writeData7 = {16'b0, writeData[9:8]};
                writeData6 = {16'b0, writeData[7:6]};
                writeData5 = {16'b0, writeData[5:4]};
                writeData4 = {16'b0, writeData[3:2]};
                writeData3 = {16'b0, writeData[1:0]};
                writeData2 = {1'b0, writeData[31:24], 1'b0, writeData[23:16]};
                writeData1 = {1'b0, writeData[15:8], 1'b0, writeData[7:0]};

                case (writeAddr[13:9])
                    5'b00000, 5'b00001, 5'b00010, 5'b00011,
                    5'b00100, 5'b00101, 5'b00110, 5'b00111,
                    5'b01000, 5'b01001, 5'b01010, 5'b01011,
                    5'b01100, 5'b01101, 5'b01110, 5'b01111 : begin
                        wen_a18 = {1'b0, wen};
                        wen_a17 = {1'b0, wen};
                        wen_a16 = {1'b0, wen};
                        wen_a15 = {1'b0, wen};
                        wen_a14 = {1'b0, wen};
                        wen_a13 = {1'b0, wen};
                        wen_a12 = {1'b0, wen};
                        wen_a11 = {1'b0, wen};
                        wen_a10 = {1'b0, wen};
                        wen_a9 = {1'b0, wen};
                        wen_a8 = {1'b0, wen};
                        wen_a7 = {1'b0, wen};
                        wen_a6 = {1'b0, wen};
                        wen_a5 = {1'b0, wen};
                        wen_a4 = {1'b0, wen};
                        wen_a3 = {1'b0, wen};
                        wen_a2 = {1'b0, 1'b0};
                        wen_a1 = {1'b0, 1'b0};
                    end
                    5'b10000, 5'b10001 : begin
                        wen_a18 = {1'b0, 1'b0};
                        wen_a17 = {1'b0, 1'b0};
                        wen_a16 = {1'b0, 1'b0};
                        wen_a15 = {1'b0, 1'b0};
                        wen_a14 = {1'b0, 1'b0};
                        wen_a13 = {1'b0, 1'b0};
                        wen_a12 = {1'b0, 1'b0};
                        wen_a11 = {1'b0, 1'b0};
                        wen_a10 = {1'b0, 1'b0};
                        wen_a9 = {1'b0, 1'b0};
                        wen_a8 = {1'b0, 1'b0};
                        wen_a7 = {1'b0, 1'b0};
                        wen_a6 = {1'b0, 1'b0};
                        wen_a5 = {1'b0, 1'b0};
                        wen_a4 = {1'b0, 1'b0};
                        wen_a3 = {1'b0, 1'b0};
                        wen_a2 = {wen, wen};
                        wen_a1 = {wen, wen};
                    end
                    default : begin
                        wen_a18 = {1'b0, 1'b0};
                        wen_a17 = {1'b0, 1'b0};
                        wen_a16 = {1'b0, 1'b0};
                        wen_a15 = {1'b0, 1'b0};
                        wen_a14 = {1'b0, 1'b0};
                        wen_a13 = {1'b0, 1'b0};
                        wen_a12 = {1'b0, 1'b0};
                        wen_a11 = {1'b0, 1'b0};
                        wen_a10 = {1'b0, 1'b0};
                        wen_a9 = {1'b0, 1'b0};
                        wen_a8 = {1'b0, 1'b0};
                        wen_a7 = {1'b0, 1'b0};
                        wen_a6 = {1'b0, 1'b0};
                        wen_a5 = {1'b0, 1'b0};
                        wen_a4 = {1'b0, 1'b0};
                        wen_a3 = {1'b0, 1'b0};
                        wen_a2 = {1'b0, 1'b0};
                        wen_a1 = {1'b0, 1'b0};
                    end
                endcase
                case (ckRdAddr[13:9])
                    5'b00000, 5'b00001, 5'b00010, 5'b00011,
                    5'b00100, 5'b00101, 5'b00110, 5'b00111,
                    5'b01000, 5'b01001, 5'b01010, 5'b01011,
                    5'b01100, 5'b01101, 5'b01110, 5'b01111 : begin
                        readData = {
                                        readData18[1:0],
                                        readData17[1:0],
                                        readData16[1:0],
                                        readData15[1:0],
                                        readData14[1:0],
                                        readData13[1:0],
                                        readData12[1:0],
                                        readData11[1:0],
                                        readData10[1:0],
                                        readData9[1:0],
                                        readData8[1:0],
                                        readData7[1:0],
                                        readData6[1:0],
                                        readData5[1:0],
                                        readData4[1:0],
                                        readData3[1:0]
                        };
                    end
                    5'b10000, 5'b10001 : begin
                        readData = {readData2[16:9],readData2[7:0],readData1[16:9],readData1[7:0]};
                    end
                    default : begin
                        readData = 32'b0;
                    end
                endcase
            end
            9728: begin
                width18 = 3'b001;
                width17 = 3'b001;
                width16 = 3'b001;
                width15 = 3'b001;
                width14 = 3'b001;
                width13 = 3'b001;
                width12 = 3'b001;
                width11 = 3'b001;
                width10 = 3'b001;
                width9 = 3'b001;
                width8 = 3'b001;
                width7 = 3'b001;
                width6 = 3'b001;
                width5 = 3'b001;
                width4 = 3'b001;
                width3 = 3'b001;
                width2 = 3'b100;
                width1 = 3'b100;
                width0 = 3'b101;

                writeAddr18 = {writeAddr[12:0], 1'b0};
                writeAddr17 = {writeAddr[12:0], 1'b0};
                writeAddr16 = {writeAddr[12:0], 1'b0};
                writeAddr15 = {writeAddr[12:0], 1'b0};
                writeAddr14 = {writeAddr[12:0], 1'b0};
                writeAddr13 = {writeAddr[12:0], 1'b0};
                writeAddr12 = {writeAddr[12:0], 1'b0};
                writeAddr11 = {writeAddr[12:0], 1'b0};
                writeAddr10 = {writeAddr[12:0], 1'b0};
                writeAddr9 = {writeAddr[12:0], 1'b0};
                writeAddr8 = {writeAddr[12:0], 1'b0};
                writeAddr7 = {writeAddr[12:0], 1'b0};
                writeAddr6 = {writeAddr[12:0], 1'b0};
                writeAddr5 = {writeAddr[12:0], 1'b0};
                writeAddr4 = {writeAddr[12:0], 1'b0};
                writeAddr3 = {writeAddr[12:0], 1'b0};
                writeAddr2 = {writeAddr[9:0], 4'b0};
                writeAddr1 = {writeAddr[9:0], 4'b0};
                writeAddr0 = {writeAddr[8:0], 5'b0};

                readAddr18  = {readAddr[12:0],  1'b0};
                readAddr17  = {readAddr[12:0],  1'b0};
                readAddr16  = {readAddr[12:0],  1'b0};
                readAddr15  = {readAddr[12:0],  1'b0};
                readAddr14  = {readAddr[12:0],  1'b0};
                readAddr13  = {readAddr[12:0],  1'b0};
                readAddr12  = {readAddr[12:0],  1'b0};
                readAddr11  = {readAddr[12:0],  1'b0};
                readAddr10  = {readAddr[12:0],  1'b0};
                readAddr9  = {readAddr[12:0],  1'b0};
                readAddr8  = {readAddr[12:0],  1'b0};
                readAddr7  = {readAddr[12:0],  1'b0};
                readAddr6  = {readAddr[12:0],  1'b0};
                readAddr5  = {readAddr[12:0],  1'b0};
                readAddr4  = {readAddr[12:0],  1'b0};
                readAddr3  = {readAddr[12:0],  1'b0};
                readAddr2  = {readAddr[9:0],  4'b0};
                readAddr1  = {readAddr[9:0],  4'b0};
                readAddr0  = {readAddr[8:0],  5'b0};

                writeData18 = {16'b0, writeData[31:30]};
                writeData17 = {16'b0, writeData[29:28]};
                writeData16 = {16'b0, writeData[27:26]};
                writeData15 = {16'b0, writeData[25:24]};
                writeData14 = {16'b0, writeData[23:22]};
                writeData13 = {16'b0, writeData[21:20]};
                writeData12 = {16'b0, writeData[19:18]};
                writeData11 = {16'b0, writeData[17:16]};
                writeData10 = {16'b0, writeData[15:14]};
                writeData9 = {16'b0, writeData[13:12]};
                writeData8 = {16'b0, writeData[11:10]};
                writeData7 = {16'b0, writeData[9:8]};
                writeData6 = {16'b0, writeData[7:6]};
                writeData5 = {16'b0, writeData[5:4]};
                writeData4 = {16'b0, writeData[3:2]};
                writeData3 = {16'b0, writeData[1:0]};
                writeData2 = {1'b0, writeData[31:24], 1'b0, writeData[23:16]};
                writeData1 = {1'b0, writeData[15:8], 1'b0, writeData[7:0]};
                writeData0 = {1'b0, writeData[31:24], 1'b0, writeData[23:16], 1'b0, writeData[15:8], 1'b0, writeData[7:0]};

                case (writeAddr[13:9])
                    5'b00000, 5'b00001, 5'b00010, 5'b00011,
                    5'b00100, 5'b00101, 5'b00110, 5'b00111,
                    5'b01000, 5'b01001, 5'b01010, 5'b01011,
                    5'b01100, 5'b01101, 5'b01110, 5'b01111 : begin
                        wen_a18 = {1'b0, wen};
                        wen_a17 = {1'b0, wen};
                        wen_a16 = {1'b0, wen};
                        wen_a15 = {1'b0, wen};
                        wen_a14 = {1'b0, wen};
                        wen_a13 = {1'b0, wen};
                        wen_a12 = {1'b0, wen};
                        wen_a11 = {1'b0, wen};
                        wen_a10 = {1'b0, wen};
                        wen_a9 = {1'b0, wen};
                        wen_a8 = {1'b0, wen};
                        wen_a7 = {1'b0, wen};
                        wen_a6 = {1'b0, wen};
                        wen_a5 = {1'b0, wen};
                        wen_a4 = {1'b0, wen};
                        wen_a3 = {1'b0, wen};
                        wen_a2 = {1'b0, 1'b0};
                        wen_a1 = {1'b0, 1'b0};
                        wen_a0 = {1'b0, 1'b0};
                        wen_b0 = {1'b0, 1'b0};
                    end
                    5'b10000, 5'b10001 : begin
                        wen_a18 = {1'b0, 1'b0};
                        wen_a17 = {1'b0, 1'b0};
                        wen_a16 = {1'b0, 1'b0};
                        wen_a15 = {1'b0, 1'b0};
                        wen_a14 = {1'b0, 1'b0};
                        wen_a13 = {1'b0, 1'b0};
                        wen_a12 = {1'b0, 1'b0};
                        wen_a11 = {1'b0, 1'b0};
                        wen_a10 = {1'b0, 1'b0};
                        wen_a9 = {1'b0, 1'b0};
                        wen_a8 = {1'b0, 1'b0};
                        wen_a7 = {1'b0, 1'b0};
                        wen_a6 = {1'b0, 1'b0};
                        wen_a5 = {1'b0, 1'b0};
                        wen_a4 = {1'b0, 1'b0};
                        wen_a3 = {1'b0, 1'b0};
                        wen_a2 = {wen, wen};
                        wen_a1 = {wen, wen};
                        wen_a0 = {1'b0, 1'b0};
                        wen_b0 = {1'b0, 1'b0};
                    end
                    5'b10010 : begin
                        wen_a18 = {1'b0, 1'b0};
                        wen_a17 = {1'b0, 1'b0};
                        wen_a16 = {1'b0, 1'b0};
                        wen_a15 = {1'b0, 1'b0};
                        wen_a14 = {1'b0, 1'b0};
                        wen_a13 = {1'b0, 1'b0};
                        wen_a12 = {1'b0, 1'b0};
                        wen_a11 = {1'b0, 1'b0};
                        wen_a10 = {1'b0, 1'b0};
                        wen_a9 = {1'b0, 1'b0};
                        wen_a8 = {1'b0, 1'b0};
                        wen_a7 = {1'b0, 1'b0};
                        wen_a6 = {1'b0, 1'b0};
                        wen_a5 = {1'b0, 1'b0};
                        wen_a4 = {1'b0, 1'b0};
                        wen_a3 = {1'b0, 1'b0};
                        wen_a2 = {1'b0, 1'b0};
                        wen_a1 = {1'b0, 1'b0};
                        wen_a0 = {wen, wen};
                        wen_b0 = {wen, wen};
                    end
                    default : begin
                        wen_a18 = {1'b0, 1'b0};
                        wen_a17 = {1'b0, 1'b0};
                        wen_a16 = {1'b0, 1'b0};
                        wen_a15 = {1'b0, 1'b0};
                        wen_a14 = {1'b0, 1'b0};
                        wen_a13 = {1'b0, 1'b0};
                        wen_a12 = {1'b0, 1'b0};
                        wen_a11 = {1'b0, 1'b0};
                        wen_a10 = {1'b0, 1'b0};
                        wen_a9 = {1'b0, 1'b0};
                        wen_a8 = {1'b0, 1'b0};
                        wen_a7 = {1'b0, 1'b0};
                        wen_a6 = {1'b0, 1'b0};
                        wen_a5 = {1'b0, 1'b0};
                        wen_a4 = {1'b0, 1'b0};
                        wen_a3 = {1'b0, 1'b0};
                        wen_a2 = {1'b0, 1'b0};
                        wen_a1 = {1'b0, 1'b0};
                        wen_a0 = {1'b0, 1'b0};
                        wen_b0 = {1'b0, 1'b0};
                    end
                endcase
                case (ckRdAddr[13:9])
                    5'b00000, 5'b00001, 5'b00010, 5'b00011,
                    5'b00100, 5'b00101, 5'b00110, 5'b00111,
                    5'b01000, 5'b01001, 5'b01010, 5'b01011,
                    5'b01100, 5'b01101, 5'b01110, 5'b01111 : begin
                        readData = {
                                        readData18[1:0],
                                        readData17[1:0],
                                        readData16[1:0],
                                        readData15[1:0],
                                        readData14[1:0],
                                        readData13[1:0],
                                        readData12[1:0],
                                        readData11[1:0],
                                        readData10[1:0],
                                        readData9[1:0],
                                        readData8[1:0],
                                        readData7[1:0],
                                        readData6[1:0],
                                        readData5[1:0],
                                        readData4[1:0],
                                        readData3[1:0]
                        };
                    end
                    5'b10000, 5'b10001 : begin
                        readData = {readData2[16:9],readData2[7:0],readData1[16:9],readData1[7:0]};
                    end
                    5'b10010 : begin
                        readData = {readData0[34:27],readData0[25:18],readData0[16:9],readData0[7:0]};
                    end
                    default : begin
                        readData = 32'b0;
                    end
                endcase
            end
            10240: begin
                width20 = 3'b001;
                width19 = 3'b001;
                width18 = 3'b001;
                width17 = 3'b001;
                width16 = 3'b001;
                width15 = 3'b001;
                width14 = 3'b001;
                width13 = 3'b001;
                width12 = 3'b001;
                width11 = 3'b001;
                width10 = 3'b001;
                width9 = 3'b001;
                width8 = 3'b001;
                width7 = 3'b001;
                width6 = 3'b001;
                width5 = 3'b001;
                width4 = 3'b011;
                width3 = 3'b011;
                width2 = 3'b011;
                width1 = 3'b011;

                writeAddr20 = {writeAddr[12:0], 1'b0};
                writeAddr19 = {writeAddr[12:0], 1'b0};
                writeAddr18 = {writeAddr[12:0], 1'b0};
                writeAddr17 = {writeAddr[12:0], 1'b0};
                writeAddr16 = {writeAddr[12:0], 1'b0};
                writeAddr15 = {writeAddr[12:0], 1'b0};
                writeAddr14 = {writeAddr[12:0], 1'b0};
                writeAddr13 = {writeAddr[12:0], 1'b0};
                writeAddr12 = {writeAddr[12:0], 1'b0};
                writeAddr11 = {writeAddr[12:0], 1'b0};
                writeAddr10 = {writeAddr[12:0], 1'b0};
                writeAddr9 = {writeAddr[12:0], 1'b0};
                writeAddr8 = {writeAddr[12:0], 1'b0};
                writeAddr7 = {writeAddr[12:0], 1'b0};
                writeAddr6 = {writeAddr[12:0], 1'b0};
                writeAddr5 = {writeAddr[12:0], 1'b0};
                writeAddr4 = {writeAddr[10:0], 3'b0};
                writeAddr3 = {writeAddr[10:0], 3'b0};
                writeAddr2 = {writeAddr[10:0], 3'b0};
                writeAddr1 = {writeAddr[10:0], 3'b0};

                readAddr20  = {readAddr[12:0],  1'b0};
                readAddr19  = {readAddr[12:0],  1'b0};
                readAddr18  = {readAddr[12:0],  1'b0};
                readAddr17  = {readAddr[12:0],  1'b0};
                readAddr16  = {readAddr[12:0],  1'b0};
                readAddr15  = {readAddr[12:0],  1'b0};
                readAddr14  = {readAddr[12:0],  1'b0};
                readAddr13  = {readAddr[12:0],  1'b0};
                readAddr12  = {readAddr[12:0],  1'b0};
                readAddr11  = {readAddr[12:0],  1'b0};
                readAddr10  = {readAddr[12:0],  1'b0};
                readAddr9  = {readAddr[12:0],  1'b0};
                readAddr8  = {readAddr[12:0],  1'b0};
                readAddr7  = {readAddr[12:0],  1'b0};
                readAddr6  = {readAddr[12:0],  1'b0};
                readAddr5  = {readAddr[12:0],  1'b0};
                readAddr4  = {readAddr[10:0],  3'b0};
                readAddr3  = {readAddr[10:0],  3'b0};
                readAddr2  = {readAddr[10:0],  3'b0};
                readAddr1  = {readAddr[10:0],  3'b0};

                writeData20 = {16'b0, writeData[31:30]};
                writeData19 = {16'b0, writeData[29:28]};
                writeData18 = {16'b0, writeData[27:26]};
                writeData17 = {16'b0, writeData[25:24]};
                writeData16 = {16'b0, writeData[23:22]};
                writeData15 = {16'b0, writeData[21:20]};
                writeData14 = {16'b0, writeData[19:18]};
                writeData13 = {16'b0, writeData[17:16]};
                writeData12 = {16'b0, writeData[15:14]};
                writeData11 = {16'b0, writeData[13:12]};
                writeData10 = {16'b0, writeData[11:10]};
                writeData9 = {16'b0, writeData[9:8]};
                writeData8 = {16'b0, writeData[7:6]};
                writeData7 = {16'b0, writeData[5:4]};
                writeData6 = {16'b0, writeData[3:2]};
                writeData5 = {16'b0, writeData[1:0]};
                writeData4 = {10'b0, writeData[31:24]};
                writeData3 = {10'b0, writeData[23:16]};
                writeData2 = {10'b0, writeData[15:8]};
                writeData1 = {10'b0, writeData[7:0]};

                case (writeAddr[13:9])
                    5'b00000, 5'b00001, 5'b00010, 5'b00011,
                    5'b00100, 5'b00101, 5'b00110, 5'b00111,
                    5'b01000, 5'b01001, 5'b01010, 5'b01011,
                    5'b01100, 5'b01101, 5'b01110, 5'b01111 : begin
                        wen_a20 = {1'b0, wen};
                        wen_a19 = {1'b0, wen};
                        wen_a18 = {1'b0, wen};
                        wen_a17 = {1'b0, wen};
                        wen_a16 = {1'b0, wen};
                        wen_a15 = {1'b0, wen};
                        wen_a14 = {1'b0, wen};
                        wen_a13 = {1'b0, wen};
                        wen_a12 = {1'b0, wen};
                        wen_a11 = {1'b0, wen};
                        wen_a10 = {1'b0, wen};
                        wen_a9 = {1'b0, wen};
                        wen_a8 = {1'b0, wen};
                        wen_a7 = {1'b0, wen};
                        wen_a6 = {1'b0, wen};
                        wen_a5 = {1'b0, wen};
                        wen_a4 = {1'b0, 1'b0};
                        wen_a3 = {1'b0, 1'b0};
                        wen_a2 = {1'b0, 1'b0};
                        wen_a1 = {1'b0, 1'b0};
                    end
                    5'b10000, 5'b10001, 5'b10010, 5'b10011 : begin
                        wen_a20 = {1'b0, 1'b0};
                        wen_a19 = {1'b0, 1'b0};
                        wen_a18 = {1'b0, 1'b0};
                        wen_a17 = {1'b0, 1'b0};
                        wen_a16 = {1'b0, 1'b0};
                        wen_a15 = {1'b0, 1'b0};
                        wen_a14 = {1'b0, 1'b0};
                        wen_a13 = {1'b0, 1'b0};
                        wen_a12 = {1'b0, 1'b0};
                        wen_a11 = {1'b0, 1'b0};
                        wen_a10 = {1'b0, 1'b0};
                        wen_a9 = {1'b0, 1'b0};
                        wen_a8 = {1'b0, 1'b0};
                        wen_a7 = {1'b0, 1'b0};
                        wen_a6 = {1'b0, 1'b0};
                        wen_a5 = {1'b0, 1'b0};
                        wen_a4 = {1'b0, wen};
                        wen_a3 = {1'b0, wen};
                        wen_a2 = {1'b0, wen};
                        wen_a1 = {1'b0, wen};
                    end
                    default : begin
                        wen_a20 = {1'b0, 1'b0};
                        wen_a19 = {1'b0, 1'b0};
                        wen_a18 = {1'b0, 1'b0};
                        wen_a17 = {1'b0, 1'b0};
                        wen_a16 = {1'b0, 1'b0};
                        wen_a15 = {1'b0, 1'b0};
                        wen_a14 = {1'b0, 1'b0};
                        wen_a13 = {1'b0, 1'b0};
                        wen_a12 = {1'b0, 1'b0};
                        wen_a11 = {1'b0, 1'b0};
                        wen_a10 = {1'b0, 1'b0};
                        wen_a9 = {1'b0, 1'b0};
                        wen_a8 = {1'b0, 1'b0};
                        wen_a7 = {1'b0, 1'b0};
                        wen_a6 = {1'b0, 1'b0};
                        wen_a5 = {1'b0, 1'b0};
                        wen_a4 = {1'b0, 1'b0};
                        wen_a3 = {1'b0, 1'b0};
                        wen_a2 = {1'b0, 1'b0};
                        wen_a1 = {1'b0, 1'b0};
                    end
                endcase
                case (ckRdAddr[13:9])
                    5'b00000, 5'b00001, 5'b00010, 5'b00011,
                    5'b00100, 5'b00101, 5'b00110, 5'b00111,
                    5'b01000, 5'b01001, 5'b01010, 5'b01011,
                    5'b01100, 5'b01101, 5'b01110, 5'b01111 : begin
                        readData = {
                                        readData20[1:0],
                                        readData19[1:0],
                                        readData18[1:0],
                                        readData17[1:0],
                                        readData16[1:0],
                                        readData15[1:0],
                                        readData14[1:0],
                                        readData13[1:0],
                                        readData12[1:0],
                                        readData11[1:0],
                                        readData10[1:0],
                                        readData9[1:0],
                                        readData8[1:0],
                                        readData7[1:0],
                                        readData6[1:0],
                                        readData5[1:0]
                        };
                    end
                    5'b10000, 5'b10001, 5'b10010, 5'b10011 : begin
                        readData = {readData4[7:0],readData3[7:0],readData2[7:0],readData1[7:0]};
                    end
                    default : begin
                        readData = 32'b0;
                    end
                endcase
            end
            10752: begin
                width20 = 3'b001;
                width19 = 3'b001;
                width18 = 3'b001;
                width17 = 3'b001;
                width16 = 3'b001;
                width15 = 3'b001;
                width14 = 3'b001;
                width13 = 3'b001;
                width12 = 3'b001;
                width11 = 3'b001;
                width10 = 3'b001;
                width9 = 3'b001;
                width8 = 3'b001;
                width7 = 3'b001;
                width6 = 3'b001;
                width5 = 3'b001;
                width4 = 3'b011;
                width3 = 3'b011;
                width2 = 3'b011;
                width1 = 3'b011;
                width0 = 3'b101;

                writeAddr20 = {writeAddr[12:0], 1'b0};
                writeAddr19 = {writeAddr[12:0], 1'b0};
                writeAddr18 = {writeAddr[12:0], 1'b0};
                writeAddr17 = {writeAddr[12:0], 1'b0};
                writeAddr16 = {writeAddr[12:0], 1'b0};
                writeAddr15 = {writeAddr[12:0], 1'b0};
                writeAddr14 = {writeAddr[12:0], 1'b0};
                writeAddr13 = {writeAddr[12:0], 1'b0};
                writeAddr12 = {writeAddr[12:0], 1'b0};
                writeAddr11 = {writeAddr[12:0], 1'b0};
                writeAddr10 = {writeAddr[12:0], 1'b0};
                writeAddr9 = {writeAddr[12:0], 1'b0};
                writeAddr8 = {writeAddr[12:0], 1'b0};
                writeAddr7 = {writeAddr[12:0], 1'b0};
                writeAddr6 = {writeAddr[12:0], 1'b0};
                writeAddr5 = {writeAddr[12:0], 1'b0};
                writeAddr4 = {writeAddr[10:0], 3'b0};
                writeAddr3 = {writeAddr[10:0], 3'b0};
                writeAddr2 = {writeAddr[10:0], 3'b0};
                writeAddr1 = {writeAddr[10:0], 3'b0};
                writeAddr0 = {writeAddr[8:0], 5'b0};

                readAddr20  = {readAddr[12:0],  1'b0};
                readAddr19  = {readAddr[12:0],  1'b0};
                readAddr18  = {readAddr[12:0],  1'b0};
                readAddr17  = {readAddr[12:0],  1'b0};
                readAddr16  = {readAddr[12:0],  1'b0};
                readAddr15  = {readAddr[12:0],  1'b0};
                readAddr14  = {readAddr[12:0],  1'b0};
                readAddr13  = {readAddr[12:0],  1'b0};
                readAddr12  = {readAddr[12:0],  1'b0};
                readAddr11  = {readAddr[12:0],  1'b0};
                readAddr10  = {readAddr[12:0],  1'b0};
                readAddr9  = {readAddr[12:0],  1'b0};
                readAddr8  = {readAddr[12:0],  1'b0};
                readAddr7  = {readAddr[12:0],  1'b0};
                readAddr6  = {readAddr[12:0],  1'b0};
                readAddr5  = {readAddr[12:0],  1'b0};
                readAddr4  = {readAddr[10:0],  3'b0};
                readAddr3  = {readAddr[10:0],  3'b0};
                readAddr2  = {readAddr[10:0],  3'b0};
                readAddr1  = {readAddr[10:0],  3'b0};
                readAddr0  = {readAddr[8:0],  5'b0};

                writeData20 = {16'b0, writeData[31:30]};
                writeData19 = {16'b0, writeData[29:28]};
                writeData18 = {16'b0, writeData[27:26]};
                writeData17 = {16'b0, writeData[25:24]};
                writeData16 = {16'b0, writeData[23:22]};
                writeData15 = {16'b0, writeData[21:20]};
                writeData14 = {16'b0, writeData[19:18]};
                writeData13 = {16'b0, writeData[17:16]};
                writeData12 = {16'b0, writeData[15:14]};
                writeData11 = {16'b0, writeData[13:12]};
                writeData10 = {16'b0, writeData[11:10]};
                writeData9 = {16'b0, writeData[9:8]};
                writeData8 = {16'b0, writeData[7:6]};
                writeData7 = {16'b0, writeData[5:4]};
                writeData6 = {16'b0, writeData[3:2]};
                writeData5 = {16'b0, writeData[1:0]};
                writeData4 = {10'b0, writeData[31:24]};
                writeData3 = {10'b0, writeData[23:16]};
                writeData2 = {10'b0, writeData[15:8]};
                writeData1 = {10'b0, writeData[7:0]};
                writeData0 = {1'b0, writeData[31:24], 1'b0, writeData[23:16], 1'b0, writeData[15:8], 1'b0, writeData[7:0]};

                case (writeAddr[13:9])
                    5'b00000, 5'b00001, 5'b00010, 5'b00011,
                    5'b00100, 5'b00101, 5'b00110, 5'b00111,
                    5'b01000, 5'b01001, 5'b01010, 5'b01011,
                    5'b01100, 5'b01101, 5'b01110, 5'b01111 : begin
                        wen_a20 = {1'b0, wen};
                        wen_a19 = {1'b0, wen};
                        wen_a18 = {1'b0, wen};
                        wen_a17 = {1'b0, wen};
                        wen_a16 = {1'b0, wen};
                        wen_a15 = {1'b0, wen};
                        wen_a14 = {1'b0, wen};
                        wen_a13 = {1'b0, wen};
                        wen_a12 = {1'b0, wen};
                        wen_a11 = {1'b0, wen};
                        wen_a10 = {1'b0, wen};
                        wen_a9 = {1'b0, wen};
                        wen_a8 = {1'b0, wen};
                        wen_a7 = {1'b0, wen};
                        wen_a6 = {1'b0, wen};
                        wen_a5 = {1'b0, wen};
                        wen_a4 = {1'b0, 1'b0};
                        wen_a3 = {1'b0, 1'b0};
                        wen_a2 = {1'b0, 1'b0};
                        wen_a1 = {1'b0, 1'b0};
                        wen_a0 = {1'b0, 1'b0};
                        wen_b0 = {1'b0, 1'b0};
                    end
                    5'b10000, 5'b10001, 5'b10010, 5'b10011 : begin
                        wen_a20 = {1'b0, 1'b0};
                        wen_a19 = {1'b0, 1'b0};
                        wen_a18 = {1'b0, 1'b0};
                        wen_a17 = {1'b0, 1'b0};
                        wen_a16 = {1'b0, 1'b0};
                        wen_a15 = {1'b0, 1'b0};
                        wen_a14 = {1'b0, 1'b0};
                        wen_a13 = {1'b0, 1'b0};
                        wen_a12 = {1'b0, 1'b0};
                        wen_a11 = {1'b0, 1'b0};
                        wen_a10 = {1'b0, 1'b0};
                        wen_a9 = {1'b0, 1'b0};
                        wen_a8 = {1'b0, 1'b0};
                        wen_a7 = {1'b0, 1'b0};
                        wen_a6 = {1'b0, 1'b0};
                        wen_a5 = {1'b0, 1'b0};
                        wen_a4 = {1'b0, wen};
                        wen_a3 = {1'b0, wen};
                        wen_a2 = {1'b0, wen};
                        wen_a1 = {1'b0, wen};
                        wen_a0 = {1'b0, 1'b0};
                        wen_b0 = {1'b0, 1'b0};
                    end
                    5'b10100 : begin
                        wen_a20 = {1'b0, 1'b0};
                        wen_a19 = {1'b0, 1'b0};
                        wen_a18 = {1'b0, 1'b0};
                        wen_a17 = {1'b0, 1'b0};
                        wen_a16 = {1'b0, 1'b0};
                        wen_a15 = {1'b0, 1'b0};
                        wen_a14 = {1'b0, 1'b0};
                        wen_a13 = {1'b0, 1'b0};
                        wen_a12 = {1'b0, 1'b0};
                        wen_a11 = {1'b0, 1'b0};
                        wen_a10 = {1'b0, 1'b0};
                        wen_a9 = {1'b0, 1'b0};
                        wen_a8 = {1'b0, 1'b0};
                        wen_a7 = {1'b0, 1'b0};
                        wen_a6 = {1'b0, 1'b0};
                        wen_a5 = {1'b0, 1'b0};
                        wen_a4 = {1'b0, 1'b0};
                        wen_a3 = {1'b0, 1'b0};
                        wen_a2 = {1'b0, 1'b0};
                        wen_a1 = {1'b0, 1'b0};
                        wen_a0 = {wen,  wen};
                        wen_b0 = {wen,  wen};
                    end
                    default : begin
                        wen_a20 = {1'b0, 1'b0};
                        wen_a19 = {1'b0, 1'b0};
                        wen_a18 = {1'b0, 1'b0};
                        wen_a17 = {1'b0, 1'b0};
                        wen_a16 = {1'b0, 1'b0};
                        wen_a15 = {1'b0, 1'b0};
                        wen_a14 = {1'b0, 1'b0};
                        wen_a13 = {1'b0, 1'b0};
                        wen_a12 = {1'b0, 1'b0};
                        wen_a11 = {1'b0, 1'b0};
                        wen_a10 = {1'b0, 1'b0};
                        wen_a9 = {1'b0, 1'b0};
                        wen_a8 = {1'b0, 1'b0};
                        wen_a7 = {1'b0, 1'b0};
                        wen_a6 = {1'b0, 1'b0};
                        wen_a5 = {1'b0, 1'b0};
                        wen_a4 = {1'b0, 1'b0};
                        wen_a3 = {1'b0, 1'b0};
                        wen_a2 = {1'b0, 1'b0};
                        wen_a1 = {1'b0, 1'b0};
                        wen_a0 = {1'b0, 1'b0};
                        wen_b0 = {1'b0, 1'b0};
                    end
                endcase
                case (ckRdAddr[13:9])
                    5'b00000, 5'b00001, 5'b00010, 5'b00011,
                    5'b00100, 5'b00101, 5'b00110, 5'b00111,
                    5'b01000, 5'b01001, 5'b01010, 5'b01011,
                    5'b01100, 5'b01101, 5'b01110, 5'b01111 : begin
                        readData = {
                                        readData20[1:0],
                                        readData19[1:0],
                                        readData18[1:0],
                                        readData17[1:0],
                                        readData16[1:0],
                                        readData15[1:0],
                                        readData14[1:0],
                                        readData13[1:0],
                                        readData12[1:0],
                                        readData11[1:0],
                                        readData10[1:0],
                                        readData9[1:0],
                                        readData8[1:0],
                                        readData7[1:0],
                                        readData6[1:0],
                                        readData5[1:0]
                        };
                    end
                    5'b10000, 5'b10001, 5'b10010, 5'b10011 : begin
                        readData = {readData4[7:0],readData3[7:0],readData2[7:0],readData1[7:0]};
                    end
                    5'b10100 : begin
                        readData = {readData0[34:27],readData0[25:18],readData0[16:9],readData0[7:0]};
                    end
                    default : begin
                        readData = 32'b0;
                    end
                endcase
            end
            11264: begin
                width22 = 3'b001;
                width21 = 3'b001;
                width20 = 3'b001;
                width19 = 3'b001;
                width18 = 3'b001;
                width17 = 3'b001;
                width16 = 3'b001;
                width15 = 3'b001;
                width14 = 3'b001;
                width13 = 3'b001;
                width12 = 3'b001;
                width11 = 3'b001;
                width10 = 3'b001;
                width9 = 3'b001;
                width8 = 3'b001;
                width7 = 3'b001;
                width6 = 3'b011;
                width5 = 3'b011;
                width4 = 3'b011;
                width3 = 3'b011;
                width2 = 3'b100;
                width1 = 3'b100;

                writeAddr22 = {writeAddr[12:0], 1'b0};
                writeAddr21 = {writeAddr[12:0], 1'b0};
                writeAddr20 = {writeAddr[12:0], 1'b0};
                writeAddr19 = {writeAddr[12:0], 1'b0};
                writeAddr18 = {writeAddr[12:0], 1'b0};
                writeAddr17 = {writeAddr[12:0], 1'b0};
                writeAddr16 = {writeAddr[12:0], 1'b0};
                writeAddr15 = {writeAddr[12:0], 1'b0};
                writeAddr14 = {writeAddr[12:0], 1'b0};
                writeAddr13 = {writeAddr[12:0], 1'b0};
                writeAddr12 = {writeAddr[12:0], 1'b0};
                writeAddr11 = {writeAddr[12:0], 1'b0};
                writeAddr10 = {writeAddr[12:0], 1'b0};
                writeAddr9 = {writeAddr[12:0], 1'b0};
                writeAddr8 = {writeAddr[12:0], 1'b0};
                writeAddr7 = {writeAddr[12:0], 1'b0};
                writeAddr6 = {writeAddr[10:0], 3'b0};
                writeAddr5 = {writeAddr[10:0], 3'b0};
                writeAddr4 = {writeAddr[10:0], 3'b0};
                writeAddr3 = {writeAddr[10:0], 3'b0};
                writeAddr2 = {writeAddr[9:0], 4'b0};
                writeAddr1 = {writeAddr[9:0], 4'b0};

                readAddr22  = {readAddr[12:0],  1'b0};
                readAddr21  = {readAddr[12:0],  1'b0};
                readAddr20  = {readAddr[12:0],  1'b0};
                readAddr19  = {readAddr[12:0],  1'b0};
                readAddr18  = {readAddr[12:0],  1'b0};
                readAddr17  = {readAddr[12:0],  1'b0};
                readAddr16  = {readAddr[12:0],  1'b0};
                readAddr15  = {readAddr[12:0],  1'b0};
                readAddr14  = {readAddr[12:0],  1'b0};
                readAddr13  = {readAddr[12:0],  1'b0};
                readAddr12  = {readAddr[12:0],  1'b0};
                readAddr11  = {readAddr[12:0],  1'b0};
                readAddr10  = {readAddr[12:0],  1'b0};
                readAddr9  = {readAddr[12:0],  1'b0};
                readAddr8  = {readAddr[12:0],  1'b0};
                readAddr7  = {readAddr[12:0],  1'b0};
                readAddr6  = {readAddr[10:0],  3'b0};
                readAddr5  = {readAddr[10:0],  3'b0};
                readAddr4  = {readAddr[10:0],  3'b0};
                readAddr3  = {readAddr[10:0],  3'b0};
                readAddr2  = {readAddr[9:0],  4'b0};
                readAddr1  = {readAddr[9:0],  4'b0};

                writeData22 = {16'b0, writeData[31:30]};
                writeData21 = {16'b0, writeData[29:28]};
                writeData20 = {16'b0, writeData[27:26]};
                writeData19 = {16'b0, writeData[25:24]};
                writeData18 = {16'b0, writeData[23:22]};
                writeData17 = {16'b0, writeData[21:20]};
                writeData16 = {16'b0, writeData[19:18]};
                writeData15 = {16'b0, writeData[17:16]};
                writeData14 = {16'b0, writeData[15:14]};
                writeData13 = {16'b0, writeData[13:12]};
                writeData12 = {16'b0, writeData[11:10]};
                writeData11 = {16'b0, writeData[9:8]};
                writeData10 = {16'b0, writeData[7:6]};
                writeData9 = {16'b0, writeData[5:4]};
                writeData8 = {16'b0, writeData[3:2]};
                writeData7 = {16'b0, writeData[1:0]};
                writeData6 = {10'b0, writeData[31:24]};
                writeData5 = {10'b0, writeData[23:16]};
                writeData4 = {10'b0, writeData[15:8]};
                writeData3 = {10'b0, writeData[7:0]};
                writeData2 = {1'b0, writeData[31:24], 1'b0, writeData[23:16]};
                writeData1 = {1'b0, writeData[15:8], 1'b0, writeData[7:0]};

                case (writeAddr[13:9])
                    5'b00000, 5'b00001, 5'b00010, 5'b00011,
                    5'b00100, 5'b00101, 5'b00110, 5'b00111,
                    5'b01000, 5'b01001, 5'b01010, 5'b01011,
                    5'b01100, 5'b01101, 5'b01110, 5'b01111 : begin
                        wen_a22 = {1'b0, wen};
                        wen_a21 = {1'b0, wen};
                        wen_a20 = {1'b0, wen};
                        wen_a19 = {1'b0, wen};
                        wen_a18 = {1'b0, wen};
                        wen_a17 = {1'b0, wen};
                        wen_a16 = {1'b0, wen};
                        wen_a15 = {1'b0, wen};
                        wen_a14 = {1'b0, wen};
                        wen_a13 = {1'b0, wen};
                        wen_a12 = {1'b0, wen};
                        wen_a11 = {1'b0, wen};
                        wen_a10 = {1'b0, wen};
                        wen_a9 = {1'b0, wen};
                        wen_a8 = {1'b0, wen};
                        wen_a7 = {1'b0, wen};
                        wen_a6 = {1'b0, 1'b0};
                        wen_a5 = {1'b0, 1'b0};
                        wen_a4 = {1'b0, 1'b0};
                        wen_a3 = {1'b0, 1'b0};
                        wen_a2 = {1'b0, 1'b0};
                        wen_a1 = {1'b0, 1'b0};
                    end
                    5'b10000, 5'b10001, 5'b10010, 5'b10011 : begin
                        wen_a22 = {1'b0, 1'b0};
                        wen_a21 = {1'b0, 1'b0};
                        wen_a20 = {1'b0, 1'b0};
                        wen_a19 = {1'b0, 1'b0};
                        wen_a18 = {1'b0, 1'b0};
                        wen_a17 = {1'b0, 1'b0};
                        wen_a16 = {1'b0, 1'b0};
                        wen_a15 = {1'b0, 1'b0};
                        wen_a14 = {1'b0, 1'b0};
                        wen_a13 = {1'b0, 1'b0};
                        wen_a12 = {1'b0, 1'b0};
                        wen_a11 = {1'b0, 1'b0};
                        wen_a10 = {1'b0, 1'b0};
                        wen_a9 = {1'b0, 1'b0};
                        wen_a8 = {1'b0, 1'b0};
                        wen_a7 = {1'b0, 1'b0};
                        wen_a6 = {1'b0, wen};
                        wen_a5 = {1'b0, wen};
                        wen_a4 = {1'b0, wen};
                        wen_a3 = {1'b0, wen};
                        wen_a2 = {1'b0, 1'b0};
                        wen_a1 = {1'b0, 1'b0};
                    end
                    5'b10100, 5'b10101 : begin
                        wen_a22 = {1'b0, 1'b0};
                        wen_a21 = {1'b0, 1'b0};
                        wen_a20 = {1'b0, 1'b0};
                        wen_a19 = {1'b0, 1'b0};
                        wen_a18 = {1'b0, 1'b0};
                        wen_a17 = {1'b0, 1'b0};
                        wen_a16 = {1'b0, 1'b0};
                        wen_a15 = {1'b0, 1'b0};
                        wen_a14 = {1'b0, 1'b0};
                        wen_a13 = {1'b0, 1'b0};
                        wen_a12 = {1'b0, 1'b0};
                        wen_a11 = {1'b0, 1'b0};
                        wen_a10 = {1'b0, 1'b0};
                        wen_a9 = {1'b0, 1'b0};
                        wen_a8 = {1'b0, 1'b0};
                        wen_a7 = {1'b0, 1'b0};
                        wen_a6 = {1'b0, 1'b0};
                        wen_a5 = {1'b0, 1'b0};
                        wen_a4 = {1'b0, 1'b0};
                        wen_a3 = {1'b0, 1'b0};
                        wen_a2 = {wen, wen};
                        wen_a1 = {wen, wen};
                    end
                    default : begin
                        wen_a22 = {1'b0, 1'b0};
                        wen_a21 = {1'b0, 1'b0};
                        wen_a20 = {1'b0, 1'b0};
                        wen_a19 = {1'b0, 1'b0};
                        wen_a18 = {1'b0, 1'b0};
                        wen_a17 = {1'b0, 1'b0};
                        wen_a16 = {1'b0, 1'b0};
                        wen_a15 = {1'b0, 1'b0};
                        wen_a14 = {1'b0, 1'b0};
                        wen_a13 = {1'b0, 1'b0};
                        wen_a12 = {1'b0, 1'b0};
                        wen_a11 = {1'b0, 1'b0};
                        wen_a10 = {1'b0, 1'b0};
                        wen_a9 = {1'b0, 1'b0};
                        wen_a8 = {1'b0, 1'b0};
                        wen_a7 = {1'b0, 1'b0};
                        wen_a6 = {1'b0, 1'b0};
                        wen_a5 = {1'b0, 1'b0};
                        wen_a4 = {1'b0, 1'b0};
                        wen_a3 = {1'b0, 1'b0};
                        wen_a2 = {1'b0, 1'b0};
                        wen_a1 = {1'b0, 1'b0};
                    end
                endcase
                case (ckRdAddr[13:9])
                    5'b00000, 5'b00001, 5'b00010, 5'b00011,
                    5'b00100, 5'b00101, 5'b00110, 5'b00111,
                    5'b01000, 5'b01001, 5'b01010, 5'b01011,
                    5'b01100, 5'b01101, 5'b01110, 5'b01111 : begin
                        readData = {
                                        readData22[1:0],
                                        readData21[1:0],
                                        readData20[1:0],
                                        readData19[1:0],
                                        readData18[1:0],
                                        readData17[1:0],
                                        readData16[1:0],
                                        readData15[1:0],
                                        readData14[1:0],
                                        readData13[1:0],
                                        readData12[1:0],
                                        readData11[1:0],
                                        readData10[1:0],
                                        readData9[1:0],
                                        readData8[1:0],
                                        readData7[1:0]
                        };
                    end
                    5'b10000, 5'b10001, 5'b10010, 5'b10011 : begin
                        readData = {readData6[7:0],readData5[7:0],readData4[7:0],readData3[7:0]};
                    end
                    5'b10100, 5'b10101 : begin
                        readData = {readData2[16:9],readData2[7:0],readData1[16:9],readData1[7:0]};
                    end
                    default : begin
                        readData = 32'b0;
                    end
                endcase
            end
            11776: begin
                width22 = 3'b001;
                width21 = 3'b001;
                width20 = 3'b001;
                width19 = 3'b001;
                width18 = 3'b001;
                width17 = 3'b001;
                width16 = 3'b001;
                width15 = 3'b001;
                width14 = 3'b001;
                width13 = 3'b001;
                width12 = 3'b001;
                width11 = 3'b001;
                width10 = 3'b001;
                width9 = 3'b001;
                width8 = 3'b001;
                width7 = 3'b001;
                width6 = 3'b011;
                width5 = 3'b011;
                width4 = 3'b011;
                width3 = 3'b011;
                width2 = 3'b100;
                width1 = 3'b100;
                width0 = 3'b101;

                writeAddr22 = {writeAddr[12:0], 1'b0};
                writeAddr21 = {writeAddr[12:0], 1'b0};
                writeAddr20 = {writeAddr[12:0], 1'b0};
                writeAddr19 = {writeAddr[12:0], 1'b0};
                writeAddr18 = {writeAddr[12:0], 1'b0};
                writeAddr17 = {writeAddr[12:0], 1'b0};
                writeAddr16 = {writeAddr[12:0], 1'b0};
                writeAddr15 = {writeAddr[12:0], 1'b0};
                writeAddr14 = {writeAddr[12:0], 1'b0};
                writeAddr13 = {writeAddr[12:0], 1'b0};
                writeAddr12 = {writeAddr[12:0], 1'b0};
                writeAddr11 = {writeAddr[12:0], 1'b0};
                writeAddr10 = {writeAddr[12:0], 1'b0};
                writeAddr9 = {writeAddr[12:0], 1'b0};
                writeAddr8 = {writeAddr[12:0], 1'b0};
                writeAddr7 = {writeAddr[12:0], 1'b0};
                writeAddr6 = {writeAddr[10:0], 3'b0};
                writeAddr5 = {writeAddr[10:0], 3'b0};
                writeAddr4 = {writeAddr[10:0], 3'b0};
                writeAddr3 = {writeAddr[10:0], 3'b0};
                writeAddr2 = {writeAddr[9:0], 4'b0};
                writeAddr1 = {writeAddr[9:0], 4'b0};
                writeAddr0 = {writeAddr[8:0], 5'b0};

                readAddr22  = {readAddr[12:0],  1'b0};
                readAddr21  = {readAddr[12:0],  1'b0};
                readAddr20  = {readAddr[12:0],  1'b0};
                readAddr19  = {readAddr[12:0],  1'b0};
                readAddr18  = {readAddr[12:0],  1'b0};
                readAddr17  = {readAddr[12:0],  1'b0};
                readAddr16  = {readAddr[12:0],  1'b0};
                readAddr15  = {readAddr[12:0],  1'b0};
                readAddr14  = {readAddr[12:0],  1'b0};
                readAddr13  = {readAddr[12:0],  1'b0};
                readAddr12  = {readAddr[12:0],  1'b0};
                readAddr11  = {readAddr[12:0],  1'b0};
                readAddr10  = {readAddr[12:0],  1'b0};
                readAddr9  = {readAddr[12:0],  1'b0};
                readAddr8  = {readAddr[12:0],  1'b0};
                readAddr7  = {readAddr[12:0],  1'b0};
                readAddr6  = {readAddr[10:0],  3'b0};
                readAddr5  = {readAddr[10:0],  3'b0};
                readAddr4  = {readAddr[10:0],  3'b0};
                readAddr3  = {readAddr[10:0],  3'b0};
                readAddr2  = {readAddr[9:0],  4'b0};
                readAddr1  = {readAddr[9:0],  4'b0};
                readAddr0  = {readAddr[8:0],  5'b0};

                writeData22 = {16'b0, writeData[31:30]};
                writeData21 = {16'b0, writeData[29:28]};
                writeData20 = {16'b0, writeData[27:26]};
                writeData19 = {16'b0, writeData[25:24]};
                writeData18 = {16'b0, writeData[23:22]};
                writeData17 = {16'b0, writeData[21:20]};
                writeData16 = {16'b0, writeData[19:18]};
                writeData15 = {16'b0, writeData[17:16]};
                writeData14 = {16'b0, writeData[15:14]};
                writeData13 = {16'b0, writeData[13:12]};
                writeData12 = {16'b0, writeData[11:10]};
                writeData11 = {16'b0, writeData[9:8]};
                writeData10 = {16'b0, writeData[7:6]};
                writeData9 = {16'b0, writeData[5:4]};
                writeData8 = {16'b0, writeData[3:2]};
                writeData7 = {16'b0, writeData[1:0]};
                writeData6 = {10'b0, writeData[31:24]};
                writeData5 = {10'b0, writeData[23:16]};
                writeData4 = {10'b0, writeData[15:8]};
                writeData3 = {10'b0, writeData[7:0]};
                writeData2 = {1'b0, writeData[31:24], 1'b0, writeData[23:16]};
                writeData1 = {1'b0, writeData[15:8], 1'b0, writeData[7:0]};
                writeData0 = {1'b0, writeData[31:24], 1'b0, writeData[23:16], 1'b0, writeData[15:8], 1'b0, writeData[7:0]};

                case (writeAddr[13:9])
                    5'b00000, 5'b00001, 5'b00010, 5'b00011,
                    5'b00100, 5'b00101, 5'b00110, 5'b00111,
                    5'b01000, 5'b01001, 5'b01010, 5'b01011,
                    5'b01100, 5'b01101, 5'b01110, 5'b01111 : begin
                        wen_a22 = {1'b0, wen};
                        wen_a21 = {1'b0, wen};
                        wen_a20 = {1'b0, wen};
                        wen_a19 = {1'b0, wen};
                        wen_a18 = {1'b0, wen};
                        wen_a17 = {1'b0, wen};
                        wen_a16 = {1'b0, wen};
                        wen_a15 = {1'b0, wen};
                        wen_a14 = {1'b0, wen};
                        wen_a13 = {1'b0, wen};
                        wen_a12 = {1'b0, wen};
                        wen_a11 = {1'b0, wen};
                        wen_a10 = {1'b0, wen};
                        wen_a9 = {1'b0, wen};
                        wen_a8 = {1'b0, wen};
                        wen_a7 = {1'b0, wen};
                        wen_a6 = {1'b0, 1'b0};
                        wen_a5 = {1'b0, 1'b0};
                        wen_a4 = {1'b0, 1'b0};
                        wen_a3 = {1'b0, 1'b0};
                        wen_a2 = {1'b0, 1'b0};
                        wen_a1 = {1'b0, 1'b0};
                        wen_a0 = {1'b0, 1'b0};
                        wen_b0 = {1'b0, 1'b0};
                    end
                    5'b10000, 5'b10001, 5'b10010, 5'b10011 : begin
                        wen_a22 = {1'b0, 1'b0};
                        wen_a21 = {1'b0, 1'b0};
                        wen_a20 = {1'b0, 1'b0};
                        wen_a19 = {1'b0, 1'b0};
                        wen_a18 = {1'b0, 1'b0};
                        wen_a17 = {1'b0, 1'b0};
                        wen_a16 = {1'b0, 1'b0};
                        wen_a15 = {1'b0, 1'b0};
                        wen_a14 = {1'b0, 1'b0};
                        wen_a13 = {1'b0, 1'b0};
                        wen_a12 = {1'b0, 1'b0};
                        wen_a11 = {1'b0, 1'b0};
                        wen_a10 = {1'b0, 1'b0};
                        wen_a9 = {1'b0, 1'b0};
                        wen_a8 = {1'b0, 1'b0};
                        wen_a7 = {1'b0, 1'b0};
                        wen_a6 = {1'b0, wen};
                        wen_a5 = {1'b0, wen};
                        wen_a4 = {1'b0, wen};
                        wen_a3 = {1'b0, wen};
                        wen_a2 = {1'b0, 1'b0};
                        wen_a1 = {1'b0, 1'b0};
                        wen_a0 = {1'b0, 1'b0};
                        wen_b0 = {1'b0, 1'b0};
                    end
                    5'b10100, 5'b10101 : begin
                        wen_a22 = {1'b0, 1'b0};
                        wen_a21 = {1'b0, 1'b0};
                        wen_a20 = {1'b0, 1'b0};
                        wen_a19 = {1'b0, 1'b0};
                        wen_a18 = {1'b0, 1'b0};
                        wen_a17 = {1'b0, 1'b0};
                        wen_a16 = {1'b0, 1'b0};
                        wen_a15 = {1'b0, 1'b0};
                        wen_a14 = {1'b0, 1'b0};
                        wen_a13 = {1'b0, 1'b0};
                        wen_a12 = {1'b0, 1'b0};
                        wen_a11 = {1'b0, 1'b0};
                        wen_a10 = {1'b0, 1'b0};
                        wen_a9 = {1'b0, 1'b0};
                        wen_a8 = {1'b0, 1'b0};
                        wen_a7 = {1'b0, 1'b0};
                        wen_a6 = {1'b0, 1'b0};
                        wen_a5 = {1'b0, 1'b0};
                        wen_a4 = {1'b0, 1'b0};
                        wen_a3 = {1'b0, 1'b0};
                        wen_a2 = {wen, wen};
                        wen_a1 = {wen, wen};
                        wen_a0 = {1'b0, 1'b0};
                        wen_b0 = {1'b0, 1'b0};
                    end
                    5'b10110 : begin
                        wen_a22 = {1'b0, 1'b0};
                        wen_a21 = {1'b0, 1'b0};
                        wen_a20 = {1'b0, 1'b0};
                        wen_a19 = {1'b0, 1'b0};
                        wen_a18 = {1'b0, 1'b0};
                        wen_a17 = {1'b0, 1'b0};
                        wen_a16 = {1'b0, 1'b0};
                        wen_a15 = {1'b0, 1'b0};
                        wen_a14 = {1'b0, 1'b0};
                        wen_a13 = {1'b0, 1'b0};
                        wen_a12 = {1'b0, 1'b0};
                        wen_a11 = {1'b0, 1'b0};
                        wen_a10 = {1'b0, 1'b0};
                        wen_a9 = {1'b0, 1'b0};
                        wen_a8 = {1'b0, 1'b0};
                        wen_a7 = {1'b0, 1'b0};
                        wen_a6 = {1'b0, 1'b0};
                        wen_a5 = {1'b0, 1'b0};
                        wen_a4 = {1'b0, 1'b0};
                        wen_a3 = {1'b0, 1'b0};
                        wen_a2 = {1'b0, 1'b0};
                        wen_a1 = {1'b0, 1'b0};
                        wen_a0 = {wen, wen};
                        wen_b0 = {wen, wen};
                    end
                    default : begin
                        wen_a22 = {1'b0, 1'b0};
                        wen_a21 = {1'b0, 1'b0};
                        wen_a20 = {1'b0, 1'b0};
                        wen_a19 = {1'b0, 1'b0};
                        wen_a18 = {1'b0, 1'b0};
                        wen_a17 = {1'b0, 1'b0};
                        wen_a16 = {1'b0, 1'b0};
                        wen_a15 = {1'b0, 1'b0};
                        wen_a14 = {1'b0, 1'b0};
                        wen_a13 = {1'b0, 1'b0};
                        wen_a12 = {1'b0, 1'b0};
                        wen_a11 = {1'b0, 1'b0};
                        wen_a10 = {1'b0, 1'b0};
                        wen_a9 = {1'b0, 1'b0};
                        wen_a8 = {1'b0, 1'b0};
                        wen_a7 = {1'b0, 1'b0};
                        wen_a6 = {1'b0, 1'b0};
                        wen_a5 = {1'b0, 1'b0};
                        wen_a4 = {1'b0, 1'b0};
                        wen_a3 = {1'b0, 1'b0};
                        wen_a2 = {1'b0, 1'b0};
                        wen_a1 = {1'b0, 1'b0};
                        wen_a0 = {1'b0, 1'b0};
                        wen_b0 = {1'b0, 1'b0};
                    end
                endcase
                case (ckRdAddr[13:9])
                    5'b00000, 5'b00001, 5'b00010, 5'b00011,
                    5'b00100, 5'b00101, 5'b00110, 5'b00111,
                    5'b01000, 5'b01001, 5'b01010, 5'b01011,
                    5'b01100, 5'b01101, 5'b01110, 5'b01111 : begin
                        readData = {
                                        readData22[1:0],
                                        readData21[1:0],
                                        readData20[1:0],
                                        readData19[1:0],
                                        readData18[1:0],
                                        readData17[1:0],
                                        readData16[1:0],
                                        readData15[1:0],
                                        readData14[1:0],
                                        readData13[1:0],
                                        readData12[1:0],
                                        readData11[1:0],
                                        readData10[1:0],
                                        readData9[1:0],
                                        readData8[1:0],
                                        readData7[1:0]
                        };
                    end
                    5'b10000, 5'b10001, 5'b10010, 5'b10011 : begin
                        readData = {readData6[7:0],readData5[7:0],readData4[7:0],readData3[7:0]};
                    end
                    5'b10100, 5'b10101 : begin
                        readData = {readData2[16:9],readData2[7:0],readData1[16:9],readData1[7:0]};
                    end
                    5'b10110 : begin
                        readData = {readData0[34:27],readData0[25:18],readData0[16:9],readData0[7:0]};
                    end
                    default : begin
                        readData = 32'b0;
                    end
                endcase
            end
            12288: begin
                width24 = 3'b001;
                width23 = 3'b001;
                width22 = 3'b001;
                width21 = 3'b001;
                width20 = 3'b001;
                width19 = 3'b001;
                width18 = 3'b001;
                width17 = 3'b001;
                width16 = 3'b001;
                width15 = 3'b001;
                width14 = 3'b001;
                width13 = 3'b001;
                width12 = 3'b001;
                width11 = 3'b001;
                width10 = 3'b001;
                width9 = 3'b001;
                width8 = 3'b010;
                width7 = 3'b010;
                width6 = 3'b010;
                width5 = 3'b010;
                width4 = 3'b010;
                width3 = 3'b010;
                width2 = 3'b010;
                width1 = 3'b010;

                writeAddr24 = {writeAddr[12:0], 1'b0};
                writeAddr23 = {writeAddr[12:0], 1'b0};
                writeAddr22 = {writeAddr[12:0], 1'b0};
                writeAddr21 = {writeAddr[12:0], 1'b0};
                writeAddr20 = {writeAddr[12:0], 1'b0};
                writeAddr19 = {writeAddr[12:0], 1'b0};
                writeAddr18 = {writeAddr[12:0], 1'b0};
                writeAddr17 = {writeAddr[12:0], 1'b0};
                writeAddr16 = {writeAddr[12:0], 1'b0};
                writeAddr15 = {writeAddr[12:0], 1'b0};
                writeAddr14 = {writeAddr[12:0], 1'b0};
                writeAddr13 = {writeAddr[12:0], 1'b0};
                writeAddr12 = {writeAddr[12:0], 1'b0};
                writeAddr11 = {writeAddr[12:0], 1'b0};
                writeAddr10 = {writeAddr[12:0], 1'b0};
                writeAddr9 = {writeAddr[12:0], 1'b0};
                writeAddr8 = {writeAddr[11:0], 2'b0};
                writeAddr7 = {writeAddr[11:0], 2'b0};
                writeAddr6 = {writeAddr[11:0], 2'b0};
                writeAddr5 = {writeAddr[11:0], 2'b0};
                writeAddr4 = {writeAddr[11:0], 2'b0};
                writeAddr3 = {writeAddr[11:0], 2'b0};
                writeAddr2 = {writeAddr[11:0], 2'b0};
                writeAddr1 = {writeAddr[11:0], 2'b0};

                readAddr24  = {readAddr[12:0],  1'b0};
                readAddr23  = {readAddr[12:0],  1'b0};
                readAddr22  = {readAddr[12:0],  1'b0};
                readAddr21  = {readAddr[12:0],  1'b0};
                readAddr20  = {readAddr[12:0],  1'b0};
                readAddr19  = {readAddr[12:0],  1'b0};
                readAddr18  = {readAddr[12:0],  1'b0};
                readAddr17  = {readAddr[12:0],  1'b0};
                readAddr16  = {readAddr[12:0],  1'b0};
                readAddr15  = {readAddr[12:0],  1'b0};
                readAddr14  = {readAddr[12:0],  1'b0};
                readAddr13  = {readAddr[12:0],  1'b0};
                readAddr12  = {readAddr[12:0],  1'b0};
                readAddr11  = {readAddr[12:0],  1'b0};
                readAddr10  = {readAddr[12:0],  1'b0};
                readAddr9  = {readAddr[12:0],  1'b0};
                readAddr8  = {readAddr[11:0],  2'b0};
                readAddr7  = {readAddr[11:0],  2'b0};
                readAddr6  = {readAddr[11:0],  2'b0};
                readAddr5  = {readAddr[11:0],  2'b0};
                readAddr4  = {readAddr[11:0],  2'b0};
                readAddr3  = {readAddr[11:0],  2'b0};
                readAddr2  = {readAddr[11:0],  2'b0};
                readAddr1  = {readAddr[11:0],  2'b0};

                writeData24 = {16'b0, writeData[31:30]};
                writeData23 = {16'b0, writeData[29:28]};
                writeData22 = {16'b0, writeData[27:26]};
                writeData21 = {16'b0, writeData[25:24]};
                writeData20 = {16'b0, writeData[23:22]};
                writeData19 = {16'b0, writeData[21:20]};
                writeData18 = {16'b0, writeData[19:18]};
                writeData17 = {16'b0, writeData[17:16]};
                writeData16 = {16'b0, writeData[15:14]};
                writeData15 = {16'b0, writeData[13:12]};
                writeData14 = {16'b0, writeData[11:10]};
                writeData13 = {16'b0, writeData[9:8]};
                writeData12 = {16'b0, writeData[7:6]};
                writeData11 = {16'b0, writeData[5:4]};
                writeData10 = {16'b0, writeData[3:2]};
                writeData9 = {16'b0, writeData[1:0]};
                writeData8 = {14'b0, writeData[31:28]};
                writeData7 = {14'b0, writeData[27:24]};
                writeData6 = {14'b0, writeData[23:20]};
                writeData5 = {14'b0, writeData[19:16]};
                writeData4 = {14'b0, writeData[15:12]};
                writeData3 = {14'b0, writeData[11:8]};
                writeData2 = {14'b0, writeData[7:4]};
                writeData1 = {14'b0, writeData[3:0]};

                case (writeAddr[13:9])
                    5'b00000, 5'b00001, 5'b00010, 5'b00011,
                    5'b00100, 5'b00101, 5'b00110, 5'b00111,
                    5'b01000, 5'b01001, 5'b01010, 5'b01011,
                    5'b01100, 5'b01101, 5'b01110, 5'b01111 : begin
                        wen_a24 = {1'b0, wen};
                        wen_a23 = {1'b0, wen};
                        wen_a22 = {1'b0, wen};
                        wen_a21 = {1'b0, wen};
                        wen_a20 = {1'b0, wen};
                        wen_a19 = {1'b0, wen};
                        wen_a18 = {1'b0, wen};
                        wen_a17 = {1'b0, wen};
                        wen_a16 = {1'b0, wen};
                        wen_a15 = {1'b0, wen};
                        wen_a14 = {1'b0, wen};
                        wen_a13 = {1'b0, wen};
                        wen_a12 = {1'b0, wen};
                        wen_a11 = {1'b0, wen};
                        wen_a10 = {1'b0, wen};
                        wen_a9 = {1'b0, wen};
                        wen_a8 = {1'b0, 1'b0};
                        wen_a7 = {1'b0, 1'b0};
                        wen_a6 = {1'b0, 1'b0};
                        wen_a5 = {1'b0, 1'b0};
                        wen_a4 = {1'b0, 1'b0};
                        wen_a3 = {1'b0, 1'b0};
                        wen_a2 = {1'b0, 1'b0};
                        wen_a1 = {1'b0, 1'b0};
                    end
                    5'b10000, 5'b10001, 5'b10010, 5'b10011,
                    5'b10100, 5'b10101, 5'b10110, 5'b10111 : begin
                        wen_a24 = {1'b0, 1'b0};
                        wen_a23 = {1'b0, 1'b0};
                        wen_a22 = {1'b0, 1'b0};
                        wen_a21 = {1'b0, 1'b0};
                        wen_a20 = {1'b0, 1'b0};
                        wen_a19 = {1'b0, 1'b0};
                        wen_a18 = {1'b0, 1'b0};
                        wen_a17 = {1'b0, 1'b0};
                        wen_a16 = {1'b0, 1'b0};
                        wen_a15 = {1'b0, 1'b0};
                        wen_a14 = {1'b0, 1'b0};
                        wen_a13 = {1'b0, 1'b0};
                        wen_a12 = {1'b0, 1'b0};
                        wen_a11 = {1'b0, 1'b0};
                        wen_a10 = {1'b0, 1'b0};
                        wen_a9 = {1'b0, 1'b0};
                        wen_a8 = {1'b0, wen};
                        wen_a7 = {1'b0, wen};
                        wen_a6 = {1'b0, wen};
                        wen_a5 = {1'b0, wen};
                        wen_a4 = {1'b0, wen};
                        wen_a3 = {1'b0, wen};
                        wen_a2 = {1'b0, wen};
                        wen_a1 = {1'b0, wen};
                    end
                    default : begin
                        wen_a24 = {1'b0, 1'b0};
                        wen_a23 = {1'b0, 1'b0};
                        wen_a22 = {1'b0, 1'b0};
                        wen_a21 = {1'b0, 1'b0};
                        wen_a20 = {1'b0, 1'b0};
                        wen_a19 = {1'b0, 1'b0};
                        wen_a18 = {1'b0, 1'b0};
                        wen_a17 = {1'b0, 1'b0};
                        wen_a16 = {1'b0, 1'b0};
                        wen_a15 = {1'b0, 1'b0};
                        wen_a14 = {1'b0, 1'b0};
                        wen_a13 = {1'b0, 1'b0};
                        wen_a12 = {1'b0, 1'b0};
                        wen_a11 = {1'b0, 1'b0};
                        wen_a10 = {1'b0, 1'b0};
                        wen_a9 = {1'b0, 1'b0};
                        wen_a8 = {1'b0, 1'b0};
                        wen_a7 = {1'b0, 1'b0};
                        wen_a6 = {1'b0, 1'b0};
                        wen_a5 = {1'b0, 1'b0};
                        wen_a4 = {1'b0, 1'b0};
                        wen_a3 = {1'b0, 1'b0};
                        wen_a2 = {1'b0, 1'b0};
                        wen_a1 = {1'b0, 1'b0};
                    end
                endcase
                case (ckRdAddr[13:9])
                    5'b00000, 5'b00001, 5'b00010, 5'b00011,
                    5'b00100, 5'b00101, 5'b00110, 5'b00111,
                    5'b01000, 5'b01001, 5'b01010, 5'b01011,
                    5'b01100, 5'b01101, 5'b01110, 5'b01111 : begin
                        readData = {
                                        readData24[1:0],
                                        readData23[1:0],
                                        readData22[1:0],
                                        readData21[1:0],
                                        readData20[1:0],
                                        readData19[1:0],
                                        readData18[1:0],
                                        readData17[1:0],
                                        readData16[1:0],
                                        readData15[1:0],
                                        readData14[1:0],
                                        readData13[1:0],
                                        readData12[1:0],
                                        readData11[1:0],
                                        readData10[1:0],
                                        readData9[1:0]
                        };
                    end
                    5'b10000, 5'b10001, 5'b10010, 5'b10011,
                    5'b10100, 5'b10101, 5'b10110, 5'b10111 : begin
                        readData = {
                                        readData8[3:0],
                                        readData7[3:0],
                                        readData6[3:0],
                                        readData5[3:0],
                                        readData4[3:0],
                                        readData3[3:0],
                                        readData2[3:0],
                                        readData1[3:0]
                        };
                    end
                    default : begin
                        readData = 32'b0;
                    end
                endcase
            end
            12800: begin
                width24 = 3'b001;
                width23 = 3'b001;
                width22 = 3'b001;
                width21 = 3'b001;
                width20 = 3'b001;
                width19 = 3'b001;
                width18 = 3'b001;
                width17 = 3'b001;
                width16 = 3'b001;
                width15 = 3'b001;
                width14 = 3'b001;
                width13 = 3'b001;
                width12 = 3'b001;
                width11 = 3'b001;
                width10 = 3'b001;
                width9 = 3'b001;
                width8 = 3'b010;
                width7 = 3'b010;
                width6 = 3'b010;
                width5 = 3'b010;
                width4 = 3'b010;
                width3 = 3'b010;
                width2 = 3'b010;
                width1 = 3'b010;
                width0 = 3'b101;

                writeAddr24 = {writeAddr[12:0], 1'b0};
                writeAddr23 = {writeAddr[12:0], 1'b0};
                writeAddr22 = {writeAddr[12:0], 1'b0};
                writeAddr21 = {writeAddr[12:0], 1'b0};
                writeAddr20 = {writeAddr[12:0], 1'b0};
                writeAddr19 = {writeAddr[12:0], 1'b0};
                writeAddr18 = {writeAddr[12:0], 1'b0};
                writeAddr17 = {writeAddr[12:0], 1'b0};
                writeAddr16 = {writeAddr[12:0], 1'b0};
                writeAddr15 = {writeAddr[12:0], 1'b0};
                writeAddr14 = {writeAddr[12:0], 1'b0};
                writeAddr13 = {writeAddr[12:0], 1'b0};
                writeAddr12 = {writeAddr[12:0], 1'b0};
                writeAddr11 = {writeAddr[12:0], 1'b0};
                writeAddr10 = {writeAddr[12:0], 1'b0};
                writeAddr9 = {writeAddr[12:0], 1'b0};
                writeAddr8 = {writeAddr[11:0], 2'b0};
                writeAddr7 = {writeAddr[11:0], 2'b0};
                writeAddr6 = {writeAddr[11:0], 2'b0};
                writeAddr5 = {writeAddr[11:0], 2'b0};
                writeAddr4 = {writeAddr[11:0], 2'b0};
                writeAddr3 = {writeAddr[11:0], 2'b0};
                writeAddr2 = {writeAddr[11:0], 2'b0};
                writeAddr1 = {writeAddr[11:0], 2'b0};
                writeAddr0 = {writeAddr[8:0], 5'b0};

                readAddr24  = {readAddr[12:0],  1'b0};
                readAddr23  = {readAddr[12:0],  1'b0};
                readAddr22  = {readAddr[12:0],  1'b0};
                readAddr21  = {readAddr[12:0],  1'b0};
                readAddr20  = {readAddr[12:0],  1'b0};
                readAddr19  = {readAddr[12:0],  1'b0};
                readAddr18  = {readAddr[12:0],  1'b0};
                readAddr17  = {readAddr[12:0],  1'b0};
                readAddr16  = {readAddr[12:0],  1'b0};
                readAddr15  = {readAddr[12:0],  1'b0};
                readAddr14  = {readAddr[12:0],  1'b0};
                readAddr13  = {readAddr[12:0],  1'b0};
                readAddr12  = {readAddr[12:0],  1'b0};
                readAddr11  = {readAddr[12:0],  1'b0};
                readAddr10  = {readAddr[12:0],  1'b0};
                readAddr9  = {readAddr[12:0],  1'b0};
                readAddr8  = {readAddr[11:0],  2'b0};
                readAddr7  = {readAddr[11:0],  2'b0};
                readAddr6  = {readAddr[11:0],  2'b0};
                readAddr5  = {readAddr[11:0],  2'b0};
                readAddr4  = {readAddr[11:0],  2'b0};
                readAddr3  = {readAddr[11:0],  2'b0};
                readAddr2  = {readAddr[11:0],  2'b0};
                readAddr1  = {readAddr[11:0],  2'b0};
                readAddr0  = {readAddr[8:0],  5'b0};

                writeData24 = {16'b0, writeData[31:30]};
                writeData23 = {16'b0, writeData[29:28]};
                writeData22 = {16'b0, writeData[27:26]};
                writeData21 = {16'b0, writeData[25:24]};
                writeData20 = {16'b0, writeData[23:22]};
                writeData19 = {16'b0, writeData[21:20]};
                writeData18 = {16'b0, writeData[19:18]};
                writeData17 = {16'b0, writeData[17:16]};
                writeData16 = {16'b0, writeData[15:14]};
                writeData15 = {16'b0, writeData[13:12]};
                writeData14 = {16'b0, writeData[11:10]};
                writeData13 = {16'b0, writeData[9:8]};
                writeData12 = {16'b0, writeData[7:6]};
                writeData11 = {16'b0, writeData[5:4]};
                writeData10 = {16'b0, writeData[3:2]};
                writeData9 = {16'b0, writeData[1:0]};
                writeData8 = {14'b0, writeData[31:28]};
                writeData7 = {14'b0, writeData[27:24]};
                writeData6 = {14'b0, writeData[23:20]};
                writeData5 = {14'b0, writeData[19:16]};
                writeData4 = {14'b0, writeData[15:12]};
                writeData3 = {14'b0, writeData[11:8]};
                writeData2 = {14'b0, writeData[7:4]};
                writeData1 = {14'b0, writeData[3:0]};
                writeData0 = {1'b0, writeData[31:24], 1'b0, writeData[23:16], 1'b0, writeData[15:8], 1'b0, writeData[7:0]};

                case (writeAddr[13:9])
                    5'b00000, 5'b00001, 5'b00010, 5'b00011,
                    5'b00100, 5'b00101, 5'b00110, 5'b00111,
                    5'b01000, 5'b01001, 5'b01010, 5'b01011,
                    5'b01100, 5'b01101, 5'b01110, 5'b01111 : begin
                        wen_a24 = {1'b0, wen};
                        wen_a23 = {1'b0, wen};
                        wen_a22 = {1'b0, wen};
                        wen_a21 = {1'b0, wen};
                        wen_a20 = {1'b0, wen};
                        wen_a19 = {1'b0, wen};
                        wen_a18 = {1'b0, wen};
                        wen_a17 = {1'b0, wen};
                        wen_a16 = {1'b0, wen};
                        wen_a15 = {1'b0, wen};
                        wen_a14 = {1'b0, wen};
                        wen_a13 = {1'b0, wen};
                        wen_a12 = {1'b0, wen};
                        wen_a11 = {1'b0, wen};
                        wen_a10 = {1'b0, wen};
                        wen_a9 = {1'b0, wen};
                        wen_a8 = {1'b0, 1'b0};
                        wen_a7 = {1'b0, 1'b0};
                        wen_a6 = {1'b0, 1'b0};
                        wen_a5 = {1'b0, 1'b0};
                        wen_a4 = {1'b0, 1'b0};
                        wen_a3 = {1'b0, 1'b0};
                        wen_a2 = {1'b0, 1'b0};
                        wen_a1 = {1'b0, 1'b0};
                        wen_a0 = {1'b0, 1'b0};
                        wen_b0 = {1'b0, 1'b0};
                    end
                    5'b10000, 5'b10001, 5'b10010, 5'b10011,
                    5'b10100, 5'b10101, 5'b10110, 5'b10111 : begin
                        wen_a24 = {1'b0, 1'b0};
                        wen_a23 = {1'b0, 1'b0};
                        wen_a22 = {1'b0, 1'b0};
                        wen_a21 = {1'b0, 1'b0};
                        wen_a20 = {1'b0, 1'b0};
                        wen_a19 = {1'b0, 1'b0};
                        wen_a18 = {1'b0, 1'b0};
                        wen_a17 = {1'b0, 1'b0};
                        wen_a16 = {1'b0, 1'b0};
                        wen_a15 = {1'b0, 1'b0};
                        wen_a14 = {1'b0, 1'b0};
                        wen_a13 = {1'b0, 1'b0};
                        wen_a12 = {1'b0, 1'b0};
                        wen_a11 = {1'b0, 1'b0};
                        wen_a10 = {1'b0, 1'b0};
                        wen_a9 = {1'b0, 1'b0};
                        wen_a8 = {1'b0, wen};
                        wen_a7 = {1'b0, wen};
                        wen_a6 = {1'b0, wen};
                        wen_a5 = {1'b0, wen};
                        wen_a4 = {1'b0, wen};
                        wen_a3 = {1'b0, wen};
                        wen_a2 = {1'b0, wen};
                        wen_a1 = {1'b0, wen};
                        wen_a0 = {1'b0, 1'b0};
                        wen_b0 = {1'b0, 1'b0};
                    end
                    5'b11000 : begin
                        wen_a24 = {1'b0, 1'b0};
                        wen_a23 = {1'b0, 1'b0};
                        wen_a22 = {1'b0, 1'b0};
                        wen_a21 = {1'b0, 1'b0};
                        wen_a20 = {1'b0, 1'b0};
                        wen_a19 = {1'b0, 1'b0};
                        wen_a18 = {1'b0, 1'b0};
                        wen_a17 = {1'b0, 1'b0};
                        wen_a16 = {1'b0, 1'b0};
                        wen_a15 = {1'b0, 1'b0};
                        wen_a14 = {1'b0, 1'b0};
                        wen_a13 = {1'b0, 1'b0};
                        wen_a12 = {1'b0, 1'b0};
                        wen_a11 = {1'b0, 1'b0};
                        wen_a10 = {1'b0, 1'b0};
                        wen_a9 = {1'b0, 1'b0};
                        wen_a8 = {1'b0, 1'b0};
                        wen_a7 = {1'b0, 1'b0};
                        wen_a6 = {1'b0, 1'b0};
                        wen_a5 = {1'b0, 1'b0};
                        wen_a4 = {1'b0, 1'b0};
                        wen_a3 = {1'b0, 1'b0};
                        wen_a2 = {1'b0, 1'b0};
                        wen_a1 = {1'b0, 1'b0};
                        wen_a0 = {wen, wen};
                        wen_b0 = {wen, wen};
                    end
                    default : begin
                        wen_a24 = {1'b0, 1'b0};
                        wen_a23 = {1'b0, 1'b0};
                        wen_a22 = {1'b0, 1'b0};
                        wen_a21 = {1'b0, 1'b0};
                        wen_a20 = {1'b0, 1'b0};
                        wen_a19 = {1'b0, 1'b0};
                        wen_a18 = {1'b0, 1'b0};
                        wen_a17 = {1'b0, 1'b0};
                        wen_a16 = {1'b0, 1'b0};
                        wen_a15 = {1'b0, 1'b0};
                        wen_a14 = {1'b0, 1'b0};
                        wen_a13 = {1'b0, 1'b0};
                        wen_a12 = {1'b0, 1'b0};
                        wen_a11 = {1'b0, 1'b0};
                        wen_a10 = {1'b0, 1'b0};
                        wen_a9 = {1'b0, 1'b0};
                        wen_a8 = {1'b0, 1'b0};
                        wen_a7 = {1'b0, 1'b0};
                        wen_a6 = {1'b0, 1'b0};
                        wen_a5 = {1'b0, 1'b0};
                        wen_a4 = {1'b0, 1'b0};
                        wen_a3 = {1'b0, 1'b0};
                        wen_a2 = {1'b0, 1'b0};
                        wen_a1 = {1'b0, 1'b0};
                        wen_a0 = {1'b0, 1'b0};
                        wen_b0 = {1'b0, 1'b0};
                    end
                endcase
                case (ckRdAddr[13:9])
                    5'b00000, 5'b00001, 5'b00010, 5'b00011,
                    5'b00100, 5'b00101, 5'b00110, 5'b00111,
                    5'b01000, 5'b01001, 5'b01010, 5'b01011,
                    5'b01100, 5'b01101, 5'b01110, 5'b01111 : begin
                        readData = {
                                        readData24[1:0],
                                        readData23[1:0],
                                        readData22[1:0],
                                        readData21[1:0],
                                        readData20[1:0],
                                        readData19[1:0],
                                        readData18[1:0],
                                        readData17[1:0],
                                        readData16[1:0],
                                        readData15[1:0],
                                        readData14[1:0],
                                        readData13[1:0],
                                        readData12[1:0],
                                        readData11[1:0],
                                        readData10[1:0],
                                        readData9[1:0]
                        };
                    end
                    5'b10000, 5'b10001, 5'b10010, 5'b10011,
                    5'b10100, 5'b10101, 5'b10110, 5'b10111 : begin
                        readData = {
                                        readData8[3:0],
                                        readData7[3:0],
                                        readData6[3:0],
                                        readData5[3:0],
                                        readData4[3:0],
                                        readData3[3:0],
                                        readData2[3:0],
                                        readData1[3:0]
                        };
                    end
                    5'b11000 : begin
                        readData = {readData0[34:27],readData0[25:18],readData0[16:9],readData0[7:0]};
                    end
                    default : begin
                        readData = 32'b0;
                    end
                endcase
            end
            13312: begin
                width26 = 3'b001;
                width25 = 3'b001;
                width24 = 3'b001;
                width23 = 3'b001;
                width22 = 3'b001;
                width21 = 3'b001;
                width20 = 3'b001;
                width19 = 3'b001;
                width18 = 3'b001;
                width17 = 3'b001;
                width16 = 3'b001;
                width15 = 3'b001;
                width14 = 3'b001;
                width13 = 3'b001;
                width12 = 3'b001;
                width11 = 3'b001;
                width10 = 3'b010;
                width9 = 3'b010;
                width8 = 3'b010;
                width7 = 3'b010;
                width6 = 3'b010;
                width5 = 3'b010;
                width4 = 3'b010;
                width3 = 3'b010;
                width2 = 3'b100;
                width1 = 3'b100;

                writeAddr26 = {writeAddr[12:0], 1'b0};
                writeAddr25 = {writeAddr[12:0], 1'b0};
                writeAddr24 = {writeAddr[12:0], 1'b0};
                writeAddr23 = {writeAddr[12:0], 1'b0};
                writeAddr22 = {writeAddr[12:0], 1'b0};
                writeAddr21 = {writeAddr[12:0], 1'b0};
                writeAddr20 = {writeAddr[12:0], 1'b0};
                writeAddr19 = {writeAddr[12:0], 1'b0};
                writeAddr18 = {writeAddr[12:0], 1'b0};
                writeAddr17 = {writeAddr[12:0], 1'b0};
                writeAddr16 = {writeAddr[12:0], 1'b0};
                writeAddr15 = {writeAddr[12:0], 1'b0};
                writeAddr14 = {writeAddr[12:0], 1'b0};
                writeAddr13 = {writeAddr[12:0], 1'b0};
                writeAddr12 = {writeAddr[12:0], 1'b0};
                writeAddr11 = {writeAddr[12:0], 1'b0};
                writeAddr10 = {writeAddr[11:0], 2'b0};
                writeAddr9 = {writeAddr[11:0], 2'b0};
                writeAddr8 = {writeAddr[11:0], 2'b0};
                writeAddr7 = {writeAddr[11:0], 2'b0};
                writeAddr6 = {writeAddr[11:0], 2'b0};
                writeAddr5 = {writeAddr[11:0], 2'b0};
                writeAddr4 = {writeAddr[11:0], 2'b0};
                writeAddr3 = {writeAddr[11:0], 2'b0};
                writeAddr2 = {writeAddr[9:0], 4'b0};
                writeAddr1 = {writeAddr[9:0], 4'b0};

                readAddr26  = {readAddr[12:0],  1'b0};
                readAddr25  = {readAddr[12:0],  1'b0};
                readAddr24  = {readAddr[12:0],  1'b0};
                readAddr23  = {readAddr[12:0],  1'b0};
                readAddr22  = {readAddr[12:0],  1'b0};
                readAddr21  = {readAddr[12:0],  1'b0};
                readAddr20  = {readAddr[12:0],  1'b0};
                readAddr19  = {readAddr[12:0],  1'b0};
                readAddr18  = {readAddr[12:0],  1'b0};
                readAddr17  = {readAddr[12:0],  1'b0};
                readAddr16  = {readAddr[12:0],  1'b0};
                readAddr15  = {readAddr[12:0],  1'b0};
                readAddr14  = {readAddr[12:0],  1'b0};
                readAddr13  = {readAddr[12:0],  1'b0};
                readAddr12  = {readAddr[12:0],  1'b0};
                readAddr11  = {readAddr[12:0],  1'b0};
                readAddr10  = {readAddr[11:0],  2'b0};
                readAddr9  = {readAddr[11:0],  2'b0};
                readAddr8  = {readAddr[11:0],  2'b0};
                readAddr7  = {readAddr[11:0],  2'b0};
                readAddr6  = {readAddr[11:0],  2'b0};
                readAddr5  = {readAddr[11:0],  2'b0};
                readAddr4  = {readAddr[11:0],  2'b0};
                readAddr3  = {readAddr[11:0],  2'b0};
                readAddr2  = {readAddr[9:0],  4'b0};
                readAddr1  = {readAddr[9:0],  4'b0};

                writeData26 = {16'b0, writeData[31:30]};
                writeData25 = {16'b0, writeData[29:28]};
                writeData24 = {16'b0, writeData[27:26]};
                writeData23 = {16'b0, writeData[25:24]};
                writeData22 = {16'b0, writeData[23:22]};
                writeData21 = {16'b0, writeData[21:20]};
                writeData20 = {16'b0, writeData[19:18]};
                writeData19 = {16'b0, writeData[17:16]};
                writeData18 = {16'b0, writeData[15:14]};
                writeData17 = {16'b0, writeData[13:12]};
                writeData16 = {16'b0, writeData[11:10]};
                writeData15 = {16'b0, writeData[9:8]};
                writeData14 = {16'b0, writeData[7:6]};
                writeData13 = {16'b0, writeData[5:4]};
                writeData12 = {16'b0, writeData[3:2]};
                writeData11 = {16'b0, writeData[1:0]};
                writeData10 = {14'b0, writeData[31:28]};
                writeData9 = {14'b0, writeData[27:24]};
                writeData8 = {14'b0, writeData[23:20]};
                writeData7 = {14'b0, writeData[19:16]};
                writeData6 = {14'b0, writeData[15:12]};
                writeData5 = {14'b0, writeData[11:8]};
                writeData4 = {14'b0, writeData[7:4]};
                writeData3 = {14'b0, writeData[3:0]};
                writeData2 = {1'b0, writeData[31:24], 1'b0, writeData[23:16]};
                writeData1 = {1'b0, writeData[15:8], 1'b0, writeData[7:0]};

                case (writeAddr[13:9])
                    5'b00000, 5'b00001, 5'b00010, 5'b00011,
                    5'b00100, 5'b00101, 5'b00110, 5'b00111,
                    5'b01000, 5'b01001, 5'b01010, 5'b01011,
                    5'b01100, 5'b01101, 5'b01110, 5'b01111 : begin
                        wen_a26 = {1'b0, wen};
                        wen_a25 = {1'b0, wen};
                        wen_a24 = {1'b0, wen};
                        wen_a23 = {1'b0, wen};
                        wen_a22 = {1'b0, wen};
                        wen_a21 = {1'b0, wen};
                        wen_a20 = {1'b0, wen};
                        wen_a19 = {1'b0, wen};
                        wen_a18 = {1'b0, wen};
                        wen_a17 = {1'b0, wen};
                        wen_a16 = {1'b0, wen};
                        wen_a15 = {1'b0, wen};
                        wen_a14 = {1'b0, wen};
                        wen_a13 = {1'b0, wen};
                        wen_a12 = {1'b0, wen};
                        wen_a11 = {1'b0, wen};
                        wen_a10 = {1'b0, 1'b0};
                        wen_a9 = {1'b0, 1'b0};
                        wen_a8 = {1'b0, 1'b0};
                        wen_a7 = {1'b0, 1'b0};
                        wen_a6 = {1'b0, 1'b0};
                        wen_a5 = {1'b0, 1'b0};
                        wen_a4 = {1'b0, 1'b0};
                        wen_a3 = {1'b0, 1'b0};
                        wen_a2 = {1'b0, 1'b0};
                        wen_a1 = {1'b0, 1'b0};
                    end
                    5'b10000, 5'b10001, 5'b10010, 5'b10011,
                    5'b10100, 5'b10101, 5'b10110, 5'b10111 : begin
                        wen_a26 = {1'b0, 1'b0};
                        wen_a25 = {1'b0, 1'b0};
                        wen_a24 = {1'b0, 1'b0};
                        wen_a23 = {1'b0, 1'b0};
                        wen_a22 = {1'b0, 1'b0};
                        wen_a21 = {1'b0, 1'b0};
                        wen_a20 = {1'b0, 1'b0};
                        wen_a19 = {1'b0, 1'b0};
                        wen_a18 = {1'b0, 1'b0};
                        wen_a17 = {1'b0, 1'b0};
                        wen_a16 = {1'b0, 1'b0};
                        wen_a15 = {1'b0, 1'b0};
                        wen_a14 = {1'b0, 1'b0};
                        wen_a13 = {1'b0, 1'b0};
                        wen_a12 = {1'b0, 1'b0};
                        wen_a11 = {1'b0, 1'b0};
                        wen_a10 = {1'b0, wen};
                        wen_a9 = {1'b0, wen};
                        wen_a8 = {1'b0, wen};
                        wen_a7 = {1'b0, wen};
                        wen_a6 = {1'b0, wen};
                        wen_a5 = {1'b0, wen};
                        wen_a4 = {1'b0, wen};
                        wen_a3 = {1'b0, wen};
                        wen_a2 = {1'b0, 1'b0};
                        wen_a1 = {1'b0, 1'b0};
                    end
                    5'b11000, 5'b11001 : begin
                        wen_a26 = {1'b0, 1'b0};
                        wen_a25 = {1'b0, 1'b0};
                        wen_a24 = {1'b0, 1'b0};
                        wen_a23 = {1'b0, 1'b0};
                        wen_a22 = {1'b0, 1'b0};
                        wen_a21 = {1'b0, 1'b0};
                        wen_a20 = {1'b0, 1'b0};
                        wen_a19 = {1'b0, 1'b0};
                        wen_a18 = {1'b0, 1'b0};
                        wen_a17 = {1'b0, 1'b0};
                        wen_a16 = {1'b0, 1'b0};
                        wen_a15 = {1'b0, 1'b0};
                        wen_a14 = {1'b0, 1'b0};
                        wen_a13 = {1'b0, 1'b0};
                        wen_a12 = {1'b0, 1'b0};
                        wen_a11 = {1'b0, 1'b0};
                        wen_a10 = {1'b0, 1'b0};
                        wen_a9 = {1'b0, 1'b0};
                        wen_a8 = {1'b0, 1'b0};
                        wen_a7 = {1'b0, 1'b0};
                        wen_a6 = {1'b0, 1'b0};
                        wen_a5 = {1'b0, 1'b0};
                        wen_a4 = {1'b0, 1'b0};
                        wen_a3 = {1'b0, 1'b0};
                        wen_a2 = {wen, wen};
                        wen_a1 = {wen, wen};
                    end
                    default : begin
                        wen_a26 = {1'b0, 1'b0};
                        wen_a25 = {1'b0, 1'b0};
                        wen_a24 = {1'b0, 1'b0};
                        wen_a23 = {1'b0, 1'b0};
                        wen_a22 = {1'b0, 1'b0};
                        wen_a21 = {1'b0, 1'b0};
                        wen_a20 = {1'b0, 1'b0};
                        wen_a19 = {1'b0, 1'b0};
                        wen_a18 = {1'b0, 1'b0};
                        wen_a17 = {1'b0, 1'b0};
                        wen_a16 = {1'b0, 1'b0};
                        wen_a15 = {1'b0, 1'b0};
                        wen_a14 = {1'b0, 1'b0};
                        wen_a13 = {1'b0, 1'b0};
                        wen_a12 = {1'b0, 1'b0};
                        wen_a11 = {1'b0, 1'b0};
                        wen_a10 = {1'b0, 1'b0};
                        wen_a9 = {1'b0, 1'b0};
                        wen_a8 = {1'b0, 1'b0};
                        wen_a7 = {1'b0, 1'b0};
                        wen_a6 = {1'b0, 1'b0};
                        wen_a5 = {1'b0, 1'b0};
                        wen_a4 = {1'b0, 1'b0};
                        wen_a3 = {1'b0, 1'b0};
                        wen_a2 = {1'b0, 1'b0};
                        wen_a1 = {1'b0, 1'b0};
                    end
                endcase
                case (ckRdAddr[13:9])
                    5'b00000, 5'b00001, 5'b00010, 5'b00011,
                    5'b00100, 5'b00101, 5'b00110, 5'b00111,
                    5'b01000, 5'b01001, 5'b01010, 5'b01011,
                    5'b01100, 5'b01101, 5'b01110, 5'b01111 : begin
                        readData = {
                                        readData26[1:0],
                                        readData25[1:0],
                                        readData24[1:0],
                                        readData23[1:0],
                                        readData22[1:0],
                                        readData21[1:0],
                                        readData20[1:0],
                                        readData19[1:0],
                                        readData18[1:0],
                                        readData17[1:0],
                                        readData16[1:0],
                                        readData15[1:0],
                                        readData14[1:0],
                                        readData13[1:0],
                                        readData12[1:0],
                                        readData11[1:0]
                        };
                    end
                    5'b10000, 5'b10001, 5'b10010, 5'b10011,
                    5'b10100, 5'b10101, 5'b10110, 5'b10111 : begin
                        readData = {
                                        readData10[3:0],
                                        readData9[3:0],
                                        readData8[3:0],
                                        readData7[3:0],
                                        readData6[3:0],
                                        readData5[3:0],
                                        readData4[3:0],
                                        readData3[3:0]
                        };
                    end
                    5'b11000, 5'b11001 : begin
                        readData = {readData2[16:9],readData2[7:0],readData1[16:9],readData1[7:0]};
                    end
                    default : begin
                        readData = 32'b0;
                    end
                endcase
            end
            13824: begin
                width26 = 3'b001;
                width25 = 3'b001;
                width24 = 3'b001;
                width23 = 3'b001;
                width22 = 3'b001;
                width21 = 3'b001;
                width20 = 3'b001;
                width19 = 3'b001;
                width18 = 3'b001;
                width17 = 3'b001;
                width16 = 3'b001;
                width15 = 3'b001;
                width14 = 3'b001;
                width13 = 3'b001;
                width12 = 3'b001;
                width11 = 3'b001;
                width10 = 3'b010;
                width9 = 3'b010;
                width8 = 3'b010;
                width7 = 3'b010;
                width6 = 3'b010;
                width5 = 3'b010;
                width4 = 3'b010;
                width3 = 3'b010;
                width2 = 3'b100;
                width1 = 3'b100;
                width0 = 3'b101;

                writeAddr26 = {writeAddr[12:0], 1'b0};
                writeAddr25 = {writeAddr[12:0], 1'b0};
                writeAddr24 = {writeAddr[12:0], 1'b0};
                writeAddr23 = {writeAddr[12:0], 1'b0};
                writeAddr22 = {writeAddr[12:0], 1'b0};
                writeAddr21 = {writeAddr[12:0], 1'b0};
                writeAddr20 = {writeAddr[12:0], 1'b0};
                writeAddr19 = {writeAddr[12:0], 1'b0};
                writeAddr18 = {writeAddr[12:0], 1'b0};
                writeAddr17 = {writeAddr[12:0], 1'b0};
                writeAddr16 = {writeAddr[12:0], 1'b0};
                writeAddr15 = {writeAddr[12:0], 1'b0};
                writeAddr14 = {writeAddr[12:0], 1'b0};
                writeAddr13 = {writeAddr[12:0], 1'b0};
                writeAddr12 = {writeAddr[12:0], 1'b0};
                writeAddr11 = {writeAddr[12:0], 1'b0};
                writeAddr10 = {writeAddr[11:0], 2'b0};
                writeAddr9 = {writeAddr[11:0], 2'b0};
                writeAddr8 = {writeAddr[11:0], 2'b0};
                writeAddr7 = {writeAddr[11:0], 2'b0};
                writeAddr6 = {writeAddr[11:0], 2'b0};
                writeAddr5 = {writeAddr[11:0], 2'b0};
                writeAddr4 = {writeAddr[11:0], 2'b0};
                writeAddr3 = {writeAddr[11:0], 2'b0};
                writeAddr2 = {writeAddr[9:0], 4'b0};
                writeAddr1 = {writeAddr[9:0], 4'b0};
                writeAddr0 = {writeAddr[8:0], 5'b0};

                readAddr26  = {readAddr[12:0],  1'b0};
                readAddr25  = {readAddr[12:0],  1'b0};
                readAddr24  = {readAddr[12:0],  1'b0};
                readAddr23  = {readAddr[12:0],  1'b0};
                readAddr22  = {readAddr[12:0],  1'b0};
                readAddr21  = {readAddr[12:0],  1'b0};
                readAddr20  = {readAddr[12:0],  1'b0};
                readAddr19  = {readAddr[12:0],  1'b0};
                readAddr18  = {readAddr[12:0],  1'b0};
                readAddr17  = {readAddr[12:0],  1'b0};
                readAddr16  = {readAddr[12:0],  1'b0};
                readAddr15  = {readAddr[12:0],  1'b0};
                readAddr14  = {readAddr[12:0],  1'b0};
                readAddr13  = {readAddr[12:0],  1'b0};
                readAddr12  = {readAddr[12:0],  1'b0};
                readAddr11  = {readAddr[12:0],  1'b0};
                readAddr10  = {readAddr[11:0],  2'b0};
                readAddr9  = {readAddr[11:0],  2'b0};
                readAddr8  = {readAddr[11:0],  2'b0};
                readAddr7  = {readAddr[11:0],  2'b0};
                readAddr6  = {readAddr[11:0],  2'b0};
                readAddr5  = {readAddr[11:0],  2'b0};
                readAddr4  = {readAddr[11:0],  2'b0};
                readAddr3  = {readAddr[11:0],  2'b0};
                readAddr2  = {readAddr[9:0],  4'b0};
                readAddr1  = {readAddr[9:0],  4'b0};
                readAddr0  = {readAddr[8:0],  5'b0};

                writeData26 = {16'b0, writeData[31:30]};
                writeData25 = {16'b0, writeData[29:28]};
                writeData24 = {16'b0, writeData[27:26]};
                writeData23 = {16'b0, writeData[25:24]};
                writeData22 = {16'b0, writeData[23:22]};
                writeData21 = {16'b0, writeData[21:20]};
                writeData20 = {16'b0, writeData[19:18]};
                writeData19 = {16'b0, writeData[17:16]};
                writeData18 = {16'b0, writeData[15:14]};
                writeData17 = {16'b0, writeData[13:12]};
                writeData16 = {16'b0, writeData[11:10]};
                writeData15 = {16'b0, writeData[9:8]};
                writeData14 = {16'b0, writeData[7:6]};
                writeData13 = {16'b0, writeData[5:4]};
                writeData12 = {16'b0, writeData[3:2]};
                writeData11 = {16'b0, writeData[1:0]};
                writeData10 = {14'b0, writeData[31:28]};
                writeData9 = {14'b0, writeData[27:24]};
                writeData8 = {14'b0, writeData[23:20]};
                writeData7 = {14'b0, writeData[19:16]};
                writeData6 = {14'b0, writeData[15:12]};
                writeData5 = {14'b0, writeData[11:8]};
                writeData4 = {14'b0, writeData[7:4]};
                writeData3 = {14'b0, writeData[3:0]};
                writeData2 = {1'b0, writeData[31:24], 1'b0, writeData[23:16]};
                writeData1 = {1'b0, writeData[15:8], 1'b0, writeData[7:0]};
                writeData0 = {1'b0, writeData[31:24], 1'b0, writeData[23:16], 1'b0, writeData[15:8], 1'b0, writeData[7:0]};

                case (writeAddr[13:9])
                    5'b00000, 5'b00001, 5'b00010, 5'b00011,
                    5'b00100, 5'b00101, 5'b00110, 5'b00111,
                    5'b01000, 5'b01001, 5'b01010, 5'b01011,
                    5'b01100, 5'b01101, 5'b01110, 5'b01111 : begin
                        wen_a26 = {1'b0, wen};
                        wen_a25 = {1'b0, wen};
                        wen_a24 = {1'b0, wen};
                        wen_a23 = {1'b0, wen};
                        wen_a22 = {1'b0, wen};
                        wen_a21 = {1'b0, wen};
                        wen_a20 = {1'b0, wen};
                        wen_a19 = {1'b0, wen};
                        wen_a18 = {1'b0, wen};
                        wen_a17 = {1'b0, wen};
                        wen_a16 = {1'b0, wen};
                        wen_a15 = {1'b0, wen};
                        wen_a14 = {1'b0, wen};
                        wen_a13 = {1'b0, wen};
                        wen_a12 = {1'b0, wen};
                        wen_a11 = {1'b0, wen};
                        wen_a10 = {1'b0, 1'b0};
                        wen_a9 = {1'b0, 1'b0};
                        wen_a8 = {1'b0, 1'b0};
                        wen_a7 = {1'b0, 1'b0};
                        wen_a6 = {1'b0, 1'b0};
                        wen_a5 = {1'b0, 1'b0};
                        wen_a4 = {1'b0, 1'b0};
                        wen_a3 = {1'b0, 1'b0};
                        wen_a2 = {1'b0, 1'b0};
                        wen_a1 = {1'b0, 1'b0};
                        wen_a0 = {1'b0, 1'b0};
                        wen_b0 = {1'b0, 1'b0};
                    end
                    5'b10000, 5'b10001, 5'b10010, 5'b10011,
                    5'b10100, 5'b10101, 5'b10110, 5'b10111 : begin
                        wen_a26 = {1'b0, 1'b0};
                        wen_a25 = {1'b0, 1'b0};
                        wen_a24 = {1'b0, 1'b0};
                        wen_a23 = {1'b0, 1'b0};
                        wen_a22 = {1'b0, 1'b0};
                        wen_a21 = {1'b0, 1'b0};
                        wen_a20 = {1'b0, 1'b0};
                        wen_a19 = {1'b0, 1'b0};
                        wen_a18 = {1'b0, 1'b0};
                        wen_a17 = {1'b0, 1'b0};
                        wen_a16 = {1'b0, 1'b0};
                        wen_a15 = {1'b0, 1'b0};
                        wen_a14 = {1'b0, 1'b0};
                        wen_a13 = {1'b0, 1'b0};
                        wen_a12 = {1'b0, 1'b0};
                        wen_a11 = {1'b0, 1'b0};
                        wen_a10 = {1'b0, wen};
                        wen_a9 = {1'b0, wen};
                        wen_a8 = {1'b0, wen};
                        wen_a7 = {1'b0, wen};
                        wen_a6 = {1'b0, wen};
                        wen_a5 = {1'b0, wen};
                        wen_a4 = {1'b0, wen};
                        wen_a3 = {1'b0, wen};
                        wen_a2 = {1'b0, 1'b0};
                        wen_a1 = {1'b0, 1'b0};
                        wen_a0 = {1'b0, 1'b0};
                        wen_b0 = {1'b0, 1'b0};
                    end
                    5'b11000, 5'b11001 : begin
                        wen_a26 = {1'b0, 1'b0};
                        wen_a25 = {1'b0, 1'b0};
                        wen_a24 = {1'b0, 1'b0};
                        wen_a23 = {1'b0, 1'b0};
                        wen_a22 = {1'b0, 1'b0};
                        wen_a21 = {1'b0, 1'b0};
                        wen_a20 = {1'b0, 1'b0};
                        wen_a19 = {1'b0, 1'b0};
                        wen_a18 = {1'b0, 1'b0};
                        wen_a17 = {1'b0, 1'b0};
                        wen_a16 = {1'b0, 1'b0};
                        wen_a15 = {1'b0, 1'b0};
                        wen_a14 = {1'b0, 1'b0};
                        wen_a13 = {1'b0, 1'b0};
                        wen_a12 = {1'b0, 1'b0};
                        wen_a11 = {1'b0, 1'b0};
                        wen_a10 = {1'b0, 1'b0};
                        wen_a9 = {1'b0, 1'b0};
                        wen_a8 = {1'b0, 1'b0};
                        wen_a7 = {1'b0, 1'b0};
                        wen_a6 = {1'b0, 1'b0};
                        wen_a5 = {1'b0, 1'b0};
                        wen_a4 = {1'b0, 1'b0};
                        wen_a3 = {1'b0, 1'b0};
                        wen_a2 = {wen, wen};
                        wen_a1 = {wen, wen};
                        wen_a0 = {1'b0, 1'b0};
                        wen_b0 = {1'b0, 1'b0};
                    end
                    5'b11010 : begin
                        wen_a26 = {1'b0, 1'b0};
                        wen_a25 = {1'b0, 1'b0};
                        wen_a24 = {1'b0, 1'b0};
                        wen_a23 = {1'b0, 1'b0};
                        wen_a22 = {1'b0, 1'b0};
                        wen_a21 = {1'b0, 1'b0};
                        wen_a20 = {1'b0, 1'b0};
                        wen_a19 = {1'b0, 1'b0};
                        wen_a18 = {1'b0, 1'b0};
                        wen_a17 = {1'b0, 1'b0};
                        wen_a16 = {1'b0, 1'b0};
                        wen_a15 = {1'b0, 1'b0};
                        wen_a14 = {1'b0, 1'b0};
                        wen_a13 = {1'b0, 1'b0};
                        wen_a12 = {1'b0, 1'b0};
                        wen_a11 = {1'b0, 1'b0};
                        wen_a10 = {1'b0, 1'b0};
                        wen_a9 = {1'b0, 1'b0};
                        wen_a8 = {1'b0, 1'b0};
                        wen_a7 = {1'b0, 1'b0};
                        wen_a6 = {1'b0, 1'b0};
                        wen_a5 = {1'b0, 1'b0};
                        wen_a4 = {1'b0, 1'b0};
                        wen_a3 = {1'b0, 1'b0};
                        wen_a2 = {1'b0, 1'b0};
                        wen_a1 = {1'b0, 1'b0};
                        wen_a0 = {wen, wen};
                        wen_b0 = {wen, wen};
                    end
                    default : begin
                        wen_a26 = {1'b0, 1'b0};
                        wen_a25 = {1'b0, 1'b0};
                        wen_a24 = {1'b0, 1'b0};
                        wen_a23 = {1'b0, 1'b0};
                        wen_a22 = {1'b0, 1'b0};
                        wen_a21 = {1'b0, 1'b0};
                        wen_a20 = {1'b0, 1'b0};
                        wen_a19 = {1'b0, 1'b0};
                        wen_a18 = {1'b0, 1'b0};
                        wen_a17 = {1'b0, 1'b0};
                        wen_a16 = {1'b0, 1'b0};
                        wen_a15 = {1'b0, 1'b0};
                        wen_a14 = {1'b0, 1'b0};
                        wen_a13 = {1'b0, 1'b0};
                        wen_a12 = {1'b0, 1'b0};
                        wen_a11 = {1'b0, 1'b0};
                        wen_a10 = {1'b0, 1'b0};
                        wen_a9 = {1'b0, 1'b0};
                        wen_a8 = {1'b0, 1'b0};
                        wen_a7 = {1'b0, 1'b0};
                        wen_a6 = {1'b0, 1'b0};
                        wen_a5 = {1'b0, 1'b0};
                        wen_a4 = {1'b0, 1'b0};
                        wen_a3 = {1'b0, 1'b0};
                        wen_a2 = {1'b0, 1'b0};
                        wen_a1 = {1'b0, 1'b0};
                        wen_a0 = {1'b0, 1'b0};
                        wen_b0 = {1'b0, 1'b0};
                    end
                endcase
                case (ckRdAddr[13:9])
                    5'b00000, 5'b00001, 5'b00010, 5'b00011,
                    5'b00100, 5'b00101, 5'b00110, 5'b00111,
                    5'b01000, 5'b01001, 5'b01010, 5'b01011,
                    5'b01100, 5'b01101, 5'b01110, 5'b01111 : begin
                        readData = {
                                        readData26[1:0],
                                        readData25[1:0],
                                        readData24[1:0],
                                        readData23[1:0],
                                        readData22[1:0],
                                        readData21[1:0],
                                        readData20[1:0],
                                        readData19[1:0],
                                        readData18[1:0],
                                        readData17[1:0],
                                        readData16[1:0],
                                        readData15[1:0],
                                        readData14[1:0],
                                        readData13[1:0],
                                        readData12[1:0],
                                        readData11[1:0]
                        };
                    end
                    5'b10000, 5'b10001, 5'b10010, 5'b10011,
                    5'b10100, 5'b10101, 5'b10110, 5'b10111 : begin
                        readData = {
                                        readData10[3:0],
                                        readData9[3:0],
                                        readData8[3:0],
                                        readData7[3:0],
                                        readData6[3:0],
                                        readData5[3:0],
                                        readData4[3:0],
                                        readData3[3:0]
                        };
                    end
                    5'b11000, 5'b11001 : begin
                        readData = {readData2[16:9],readData2[7:0],readData1[16:9],readData1[7:0]};
                    end
                    5'b11010 : begin
                        readData = {readData0[34:27],readData0[25:18],readData0[16:9],readData0[7:0]};
                    end
                    default : begin
                        readData = 32'b0;
                    end
                endcase
            end
            14336: begin
                width28 = 3'b001;
                width27 = 3'b001;
                width26 = 3'b001;
                width25 = 3'b001;
                width24 = 3'b001;
                width23 = 3'b001;
                width22 = 3'b001;
                width21 = 3'b001;
                width20 = 3'b001;
                width19 = 3'b001;
                width18 = 3'b001;
                width17 = 3'b001;
                width16 = 3'b001;
                width15 = 3'b001;
                width14 = 3'b001;
                width13 = 3'b001;
                width12 = 3'b010;
                width11 = 3'b010;
                width10 = 3'b010;
                width9 = 3'b010;
                width8 = 3'b010;
                width7 = 3'b010;
                width6 = 3'b010;
                width5 = 3'b010;
                width4 = 3'b011;
                width3 = 3'b011;
                width2 = 3'b011;
                width1 = 3'b011;

                writeAddr28 = {writeAddr[12:0], 1'b0};
                writeAddr27 = {writeAddr[12:0], 1'b0};
                writeAddr26 = {writeAddr[12:0], 1'b0};
                writeAddr25 = {writeAddr[12:0], 1'b0};
                writeAddr24 = {writeAddr[12:0], 1'b0};
                writeAddr23 = {writeAddr[12:0], 1'b0};
                writeAddr22 = {writeAddr[12:0], 1'b0};
                writeAddr21 = {writeAddr[12:0], 1'b0};
                writeAddr20 = {writeAddr[12:0], 1'b0};
                writeAddr19 = {writeAddr[12:0], 1'b0};
                writeAddr18 = {writeAddr[12:0], 1'b0};
                writeAddr17 = {writeAddr[12:0], 1'b0};
                writeAddr16 = {writeAddr[12:0], 1'b0};
                writeAddr15 = {writeAddr[12:0], 1'b0};
                writeAddr14 = {writeAddr[12:0], 1'b0};
                writeAddr13 = {writeAddr[12:0], 1'b0};
                writeAddr12 = {writeAddr[11:0], 2'b0};
                writeAddr11 = {writeAddr[11:0], 2'b0};
                writeAddr10 = {writeAddr[11:0], 2'b0};
                writeAddr9 = {writeAddr[11:0], 2'b0};
                writeAddr8 = {writeAddr[11:0], 2'b0};
                writeAddr7 = {writeAddr[11:0], 2'b0};
                writeAddr6 = {writeAddr[11:0], 2'b0};
                writeAddr5 = {writeAddr[11:0], 2'b0};
                writeAddr4 = {writeAddr[10:0], 3'b0};
                writeAddr3 = {writeAddr[10:0], 3'b0};
                writeAddr2 = {writeAddr[10:0], 3'b0};
                writeAddr1 = {writeAddr[10:0], 3'b0};

                readAddr28  = {readAddr[12:0],  1'b0};
                readAddr27  = {readAddr[12:0],  1'b0};
                readAddr26  = {readAddr[12:0],  1'b0};
                readAddr25  = {readAddr[12:0],  1'b0};
                readAddr24  = {readAddr[12:0],  1'b0};
                readAddr23  = {readAddr[12:0],  1'b0};
                readAddr22  = {readAddr[12:0],  1'b0};
                readAddr21  = {readAddr[12:0],  1'b0};
                readAddr20  = {readAddr[12:0],  1'b0};
                readAddr19  = {readAddr[12:0],  1'b0};
                readAddr18  = {readAddr[12:0],  1'b0};
                readAddr17  = {readAddr[12:0],  1'b0};
                readAddr16  = {readAddr[12:0],  1'b0};
                readAddr15  = {readAddr[12:0],  1'b0};
                readAddr14  = {readAddr[12:0],  1'b0};
                readAddr13  = {readAddr[12:0],  1'b0};
                readAddr12  = {readAddr[11:0],  2'b0};
                readAddr11  = {readAddr[11:0],  2'b0};
                readAddr10  = {readAddr[11:0],  2'b0};
                readAddr9  = {readAddr[11:0],  2'b0};
                readAddr8  = {readAddr[11:0],  2'b0};
                readAddr7  = {readAddr[11:0],  2'b0};
                readAddr6  = {readAddr[11:0],  2'b0};
                readAddr5  = {readAddr[11:0],  2'b0};
                readAddr4  = {readAddr[10:0],  3'b0};
                readAddr3  = {readAddr[10:0],  3'b0};
                readAddr2  = {readAddr[10:0],  3'b0};
                readAddr1  = {readAddr[10:0],  3'b0};

                writeData28 = {16'b0, writeData[31:30]};
                writeData27 = {16'b0, writeData[29:28]};
                writeData26 = {16'b0, writeData[27:26]};
                writeData25 = {16'b0, writeData[25:24]};
                writeData24 = {16'b0, writeData[23:22]};
                writeData23 = {16'b0, writeData[21:20]};
                writeData22 = {16'b0, writeData[19:18]};
                writeData21 = {16'b0, writeData[17:16]};
                writeData20 = {16'b0, writeData[15:14]};
                writeData19 = {16'b0, writeData[13:12]};
                writeData18 = {16'b0, writeData[11:10]};
                writeData17 = {16'b0, writeData[9:8]};
                writeData16 = {16'b0, writeData[7:6]};
                writeData15 = {16'b0, writeData[5:4]};
                writeData14 = {16'b0, writeData[3:2]};
                writeData13 = {16'b0, writeData[1:0]};
                writeData12 = {14'b0, writeData[31:28]};
                writeData11 = {14'b0, writeData[27:24]};
                writeData10 = {14'b0, writeData[23:20]};
                writeData9 = {14'b0, writeData[19:16]};
                writeData8 = {14'b0, writeData[15:12]};
                writeData7 = {14'b0, writeData[11:8]};
                writeData6 = {14'b0, writeData[7:4]};
                writeData5 = {14'b0, writeData[3:0]};
                writeData4 = {10'b0, writeData[31:24]};
                writeData3 = {10'b0, writeData[23:16]};
                writeData2 = {10'b0, writeData[15:8]};
                writeData1 = {10'b0, writeData[7:0]};

                case (writeAddr[13:9])
                    5'b00000, 5'b00001, 5'b00010, 5'b00011,
                    5'b00100, 5'b00101, 5'b00110, 5'b00111,
                    5'b01000, 5'b01001, 5'b01010, 5'b01011,
                    5'b01100, 5'b01101, 5'b01110, 5'b01111 : begin
                        wen_a28 = {1'b0, wen};
                        wen_a27 = {1'b0, wen};
                        wen_a26 = {1'b0, wen};
                        wen_a25 = {1'b0, wen};
                        wen_a24 = {1'b0, wen};
                        wen_a23 = {1'b0, wen};
                        wen_a22 = {1'b0, wen};
                        wen_a21 = {1'b0, wen};
                        wen_a20 = {1'b0, wen};
                        wen_a19 = {1'b0, wen};
                        wen_a18 = {1'b0, wen};
                        wen_a17 = {1'b0, wen};
                        wen_a16 = {1'b0, wen};
                        wen_a15 = {1'b0, wen};
                        wen_a14 = {1'b0, wen};
                        wen_a13 = {1'b0, wen};
                        wen_a12 = {1'b0, 1'b0};
                        wen_a11 = {1'b0, 1'b0};
                        wen_a10 = {1'b0, 1'b0};
                        wen_a9 = {1'b0, 1'b0};
                        wen_a8 = {1'b0, 1'b0};
                        wen_a7 = {1'b0, 1'b0};
                        wen_a6 = {1'b0, 1'b0};
                        wen_a5 = {1'b0, 1'b0};
                        wen_a4 = {1'b0, 1'b0};
                        wen_a3 = {1'b0, 1'b0};
                        wen_a2 = {1'b0, 1'b0};
                        wen_a1 = {1'b0, 1'b0};
                    end
                    5'b10000, 5'b10001, 5'b10010, 5'b10011,
                    5'b10100, 5'b10101, 5'b10110, 5'b10111 : begin
                        wen_a28 = {1'b0, 1'b0};
                        wen_a27 = {1'b0, 1'b0};
                        wen_a26 = {1'b0, 1'b0};
                        wen_a25 = {1'b0, 1'b0};
                        wen_a24 = {1'b0, 1'b0};
                        wen_a23 = {1'b0, 1'b0};
                        wen_a22 = {1'b0, 1'b0};
                        wen_a21 = {1'b0, 1'b0};
                        wen_a20 = {1'b0, 1'b0};
                        wen_a19 = {1'b0, 1'b0};
                        wen_a18 = {1'b0, 1'b0};
                        wen_a17 = {1'b0, 1'b0};
                        wen_a16 = {1'b0, 1'b0};
                        wen_a15 = {1'b0, 1'b0};
                        wen_a14 = {1'b0, 1'b0};
                        wen_a13 = {1'b0, 1'b0};
                        wen_a12 = {1'b0, wen};
                        wen_a11 = {1'b0, wen};
                        wen_a10 = {1'b0, wen};
                        wen_a9 = {1'b0, wen};
                        wen_a8 = {1'b0, wen};
                        wen_a7 = {1'b0, wen};
                        wen_a6 = {1'b0, wen};
                        wen_a5 = {1'b0, wen};
                        wen_a4 = {1'b0, 1'b0};
                        wen_a3 = {1'b0, 1'b0};
                        wen_a2 = {1'b0, 1'b0};
                        wen_a1 = {1'b0, 1'b0};
                    end
                    5'b11000, 5'b11001, 5'b11010, 5'b11011 : begin
                        wen_a28 = {1'b0, 1'b0};
                        wen_a27 = {1'b0, 1'b0};
                        wen_a26 = {1'b0, 1'b0};
                        wen_a25 = {1'b0, 1'b0};
                        wen_a24 = {1'b0, 1'b0};
                        wen_a23 = {1'b0, 1'b0};
                        wen_a22 = {1'b0, 1'b0};
                        wen_a21 = {1'b0, 1'b0};
                        wen_a20 = {1'b0, 1'b0};
                        wen_a19 = {1'b0, 1'b0};
                        wen_a18 = {1'b0, 1'b0};
                        wen_a17 = {1'b0, 1'b0};
                        wen_a16 = {1'b0, 1'b0};
                        wen_a15 = {1'b0, 1'b0};
                        wen_a14 = {1'b0, 1'b0};
                        wen_a13 = {1'b0, 1'b0};
                        wen_a12 = {1'b0, 1'b0};
                        wen_a11 = {1'b0, 1'b0};
                        wen_a10 = {1'b0, 1'b0};
                        wen_a9 = {1'b0, 1'b0};
                        wen_a8 = {1'b0, 1'b0};
                        wen_a7 = {1'b0, 1'b0};
                        wen_a6 = {1'b0, 1'b0};
                        wen_a5 = {1'b0, 1'b0};
                        wen_a4 = {1'b0, wen};
                        wen_a3 = {1'b0, wen};
                        wen_a2 = {1'b0, wen};
                        wen_a1 = {1'b0, wen};
                    end
                    default : begin
                        wen_a28 = {1'b0, 1'b0};
                        wen_a27 = {1'b0, 1'b0};
                        wen_a26 = {1'b0, 1'b0};
                        wen_a25 = {1'b0, 1'b0};
                        wen_a24 = {1'b0, 1'b0};
                        wen_a23 = {1'b0, 1'b0};
                        wen_a22 = {1'b0, 1'b0};
                        wen_a21 = {1'b0, 1'b0};
                        wen_a20 = {1'b0, 1'b0};
                        wen_a19 = {1'b0, 1'b0};
                        wen_a18 = {1'b0, 1'b0};
                        wen_a17 = {1'b0, 1'b0};
                        wen_a16 = {1'b0, 1'b0};
                        wen_a15 = {1'b0, 1'b0};
                        wen_a14 = {1'b0, 1'b0};
                        wen_a13 = {1'b0, 1'b0};
                        wen_a12 = {1'b0, 1'b0};
                        wen_a11 = {1'b0, 1'b0};
                        wen_a10 = {1'b0, 1'b0};
                        wen_a9 = {1'b0, 1'b0};
                        wen_a8 = {1'b0, 1'b0};
                        wen_a7 = {1'b0, 1'b0};
                        wen_a6 = {1'b0, 1'b0};
                        wen_a5 = {1'b0, 1'b0};
                        wen_a4 = {1'b0, 1'b0};
                        wen_a3 = {1'b0, 1'b0};
                        wen_a2 = {1'b0, 1'b0};
                        wen_a1 = {1'b0, 1'b0};
                    end
                endcase
                case (ckRdAddr[13:9])
                    5'b00000, 5'b00001, 5'b00010, 5'b00011,
                    5'b00100, 5'b00101, 5'b00110, 5'b00111,
                    5'b01000, 5'b01001, 5'b01010, 5'b01011,
                    5'b01100, 5'b01101, 5'b01110, 5'b01111 : begin
                        readData = {
                                        readData28[1:0],
                                        readData27[1:0],
                                        readData26[1:0],
                                        readData25[1:0],
                                        readData24[1:0],
                                        readData23[1:0],
                                        readData22[1:0],
                                        readData21[1:0],
                                        readData20[1:0],
                                        readData19[1:0],
                                        readData18[1:0],
                                        readData17[1:0],
                                        readData16[1:0],
                                        readData15[1:0],
                                        readData14[1:0],
                                        readData13[1:0]
                        };
                    end
                    5'b10000, 5'b10001, 5'b10010, 5'b10011,
                    5'b10100, 5'b10101, 5'b10110, 5'b10111 : begin
                        readData = {
                                        readData12[3:0],
                                        readData11[3:0],
                                        readData10[3:0],
                                        readData9[3:0],
                                        readData8[3:0],
                                        readData7[3:0],
                                        readData6[3:0],
                                        readData5[3:0]
                        };
                    end
                    5'b11000, 5'b11001, 5'b11010, 5'b11011 : begin
                        readData = {readData4[7:0],readData3[7:0],readData2[7:0],readData1[7:0]};
                    end
                    default : begin
                        readData = 32'b0;
                    end
                endcase
            end
            14848: begin
                width28 = 3'b001;
                width27 = 3'b001;
                width26 = 3'b001;
                width25 = 3'b001;
                width24 = 3'b001;
                width23 = 3'b001;
                width22 = 3'b001;
                width21 = 3'b001;
                width20 = 3'b001;
                width19 = 3'b001;
                width18 = 3'b001;
                width17 = 3'b001;
                width16 = 3'b001;
                width15 = 3'b001;
                width14 = 3'b001;
                width13 = 3'b001;
                width12 = 3'b010;
                width11 = 3'b010;
                width10 = 3'b010;
                width9 = 3'b010;
                width8 = 3'b010;
                width7 = 3'b010;
                width6 = 3'b010;
                width5 = 3'b010;
                width4 = 3'b011;
                width3 = 3'b011;
                width2 = 3'b011;
                width1 = 3'b011;
                width0 = 3'b101;

                writeAddr28 = {writeAddr[12:0], 1'b0};
                writeAddr27 = {writeAddr[12:0], 1'b0};
                writeAddr26 = {writeAddr[12:0], 1'b0};
                writeAddr25 = {writeAddr[12:0], 1'b0};
                writeAddr24 = {writeAddr[12:0], 1'b0};
                writeAddr23 = {writeAddr[12:0], 1'b0};
                writeAddr22 = {writeAddr[12:0], 1'b0};
                writeAddr21 = {writeAddr[12:0], 1'b0};
                writeAddr20 = {writeAddr[12:0], 1'b0};
                writeAddr19 = {writeAddr[12:0], 1'b0};
                writeAddr18 = {writeAddr[12:0], 1'b0};
                writeAddr17 = {writeAddr[12:0], 1'b0};
                writeAddr16 = {writeAddr[12:0], 1'b0};
                writeAddr15 = {writeAddr[12:0], 1'b0};
                writeAddr14 = {writeAddr[12:0], 1'b0};
                writeAddr13 = {writeAddr[12:0], 1'b0};
                writeAddr12 = {writeAddr[11:0], 2'b0};
                writeAddr11 = {writeAddr[11:0], 2'b0};
                writeAddr10 = {writeAddr[11:0], 2'b0};
                writeAddr9 = {writeAddr[11:0], 2'b0};
                writeAddr8 = {writeAddr[11:0], 2'b0};
                writeAddr7 = {writeAddr[11:0], 2'b0};
                writeAddr6 = {writeAddr[11:0], 2'b0};
                writeAddr5 = {writeAddr[11:0], 2'b0};
                writeAddr4 = {writeAddr[10:0], 3'b0};
                writeAddr3 = {writeAddr[10:0], 3'b0};
                writeAddr2 = {writeAddr[10:0], 3'b0};
                writeAddr1 = {writeAddr[10:0], 3'b0};
                writeAddr0 = {writeAddr[8:0], 5'b0};

                readAddr28  = {readAddr[12:0],  1'b0};
                readAddr27  = {readAddr[12:0],  1'b0};
                readAddr26  = {readAddr[12:0],  1'b0};
                readAddr25  = {readAddr[12:0],  1'b0};
                readAddr24  = {readAddr[12:0],  1'b0};
                readAddr23  = {readAddr[12:0],  1'b0};
                readAddr22  = {readAddr[12:0],  1'b0};
                readAddr21  = {readAddr[12:0],  1'b0};
                readAddr20  = {readAddr[12:0],  1'b0};
                readAddr19  = {readAddr[12:0],  1'b0};
                readAddr18  = {readAddr[12:0],  1'b0};
                readAddr17  = {readAddr[12:0],  1'b0};
                readAddr16  = {readAddr[12:0],  1'b0};
                readAddr15  = {readAddr[12:0],  1'b0};
                readAddr14  = {readAddr[12:0],  1'b0};
                readAddr13  = {readAddr[12:0],  1'b0};
                readAddr12  = {readAddr[11:0],  2'b0};
                readAddr11  = {readAddr[11:0],  2'b0};
                readAddr10  = {readAddr[11:0],  2'b0};
                readAddr9  = {readAddr[11:0],  2'b0};
                readAddr8  = {readAddr[11:0],  2'b0};
                readAddr7  = {readAddr[11:0],  2'b0};
                readAddr6  = {readAddr[11:0],  2'b0};
                readAddr5  = {readAddr[11:0],  2'b0};
                readAddr4  = {readAddr[10:0],  3'b0};
                readAddr3  = {readAddr[10:0],  3'b0};
                readAddr2  = {readAddr[10:0],  3'b0};
                readAddr1  = {readAddr[10:0],  3'b0};
                readAddr0  = {readAddr[8:0],  5'b0};

                writeData28 = {16'b0, writeData[31:30]};
                writeData27 = {16'b0, writeData[29:28]};
                writeData26 = {16'b0, writeData[27:26]};
                writeData25 = {16'b0, writeData[25:24]};
                writeData24 = {16'b0, writeData[23:22]};
                writeData23 = {16'b0, writeData[21:20]};
                writeData22 = {16'b0, writeData[19:18]};
                writeData21 = {16'b0, writeData[17:16]};
                writeData20 = {16'b0, writeData[15:14]};
                writeData19 = {16'b0, writeData[13:12]};
                writeData18 = {16'b0, writeData[11:10]};
                writeData17 = {16'b0, writeData[9:8]};
                writeData16 = {16'b0, writeData[7:6]};
                writeData15 = {16'b0, writeData[5:4]};
                writeData14 = {16'b0, writeData[3:2]};
                writeData13 = {16'b0, writeData[1:0]};
                writeData12 = {14'b0, writeData[31:28]};
                writeData11 = {14'b0, writeData[27:24]};
                writeData10 = {14'b0, writeData[23:20]};
                writeData9 = {14'b0, writeData[19:16]};
                writeData8 = {14'b0, writeData[15:12]};
                writeData7 = {14'b0, writeData[11:8]};
                writeData6 = {14'b0, writeData[7:4]};
                writeData5 = {14'b0, writeData[3:0]};
                writeData4 = {10'b0, writeData[31:24]};
                writeData3 = {10'b0, writeData[23:16]};
                writeData2 = {10'b0, writeData[15:8]};
                writeData1 = {10'b0, writeData[7:0]};
                writeData0 = {1'b0, writeData[31:24], 1'b0, writeData[23:16], 1'b0, writeData[15:8], 1'b0, writeData[7:0]};

                case (writeAddr[13:9])
                    5'b00000, 5'b00001, 5'b00010, 5'b00011,
                    5'b00100, 5'b00101, 5'b00110, 5'b00111,
                    5'b01000, 5'b01001, 5'b01010, 5'b01011,
                    5'b01100, 5'b01101, 5'b01110, 5'b01111 : begin
                        wen_a28 = {1'b0, wen};
                        wen_a27 = {1'b0, wen};
                        wen_a26 = {1'b0, wen};
                        wen_a25 = {1'b0, wen};
                        wen_a24 = {1'b0, wen};
                        wen_a23 = {1'b0, wen};
                        wen_a22 = {1'b0, wen};
                        wen_a21 = {1'b0, wen};
                        wen_a20 = {1'b0, wen};
                        wen_a19 = {1'b0, wen};
                        wen_a18 = {1'b0, wen};
                        wen_a17 = {1'b0, wen};
                        wen_a16 = {1'b0, wen};
                        wen_a15 = {1'b0, wen};
                        wen_a14 = {1'b0, wen};
                        wen_a13 = {1'b0, wen};
                        wen_a12 = {1'b0, 1'b0};
                        wen_a11 = {1'b0, 1'b0};
                        wen_a10 = {1'b0, 1'b0};
                        wen_a9 = {1'b0, 1'b0};
                        wen_a8 = {1'b0, 1'b0};
                        wen_a7 = {1'b0, 1'b0};
                        wen_a6 = {1'b0, 1'b0};
                        wen_a5 = {1'b0, 1'b0};
                        wen_a4 = {1'b0, 1'b0};
                        wen_a3 = {1'b0, 1'b0};
                        wen_a2 = {1'b0, 1'b0};
                        wen_a1 = {1'b0, 1'b0};
                        wen_a0 = {1'b0, 1'b0};
                        wen_b0 = {1'b0, 1'b0};
                    end
                    5'b10000, 5'b10001, 5'b10010, 5'b10011,
                    5'b10100, 5'b10101, 5'b10110, 5'b10111 : begin
                        wen_a28 = {1'b0, 1'b0};
                        wen_a27 = {1'b0, 1'b0};
                        wen_a26 = {1'b0, 1'b0};
                        wen_a25 = {1'b0, 1'b0};
                        wen_a24 = {1'b0, 1'b0};
                        wen_a23 = {1'b0, 1'b0};
                        wen_a22 = {1'b0, 1'b0};
                        wen_a21 = {1'b0, 1'b0};
                        wen_a20 = {1'b0, 1'b0};
                        wen_a19 = {1'b0, 1'b0};
                        wen_a18 = {1'b0, 1'b0};
                        wen_a17 = {1'b0, 1'b0};
                        wen_a16 = {1'b0, 1'b0};
                        wen_a15 = {1'b0, 1'b0};
                        wen_a14 = {1'b0, 1'b0};
                        wen_a13 = {1'b0, 1'b0};
                        wen_a12 = {1'b0, wen};
                        wen_a11 = {1'b0, wen};
                        wen_a10 = {1'b0, wen};
                        wen_a9 = {1'b0, wen};
                        wen_a8 = {1'b0, wen};
                        wen_a7 = {1'b0, wen};
                        wen_a6 = {1'b0, wen};
                        wen_a5 = {1'b0, wen};
                        wen_a4 = {1'b0, 1'b0};
                        wen_a3 = {1'b0, 1'b0};
                        wen_a2 = {1'b0, 1'b0};
                        wen_a1 = {1'b0, 1'b0};
                        wen_a0 = {1'b0, 1'b0};
                        wen_b0 = {1'b0, 1'b0};
                    end
                    5'b11000, 5'b11001, 5'b11010, 5'b11011 : begin
                        wen_a28 = {1'b0, 1'b0};
                        wen_a27 = {1'b0, 1'b0};
                        wen_a26 = {1'b0, 1'b0};
                        wen_a25 = {1'b0, 1'b0};
                        wen_a24 = {1'b0, 1'b0};
                        wen_a23 = {1'b0, 1'b0};
                        wen_a22 = {1'b0, 1'b0};
                        wen_a21 = {1'b0, 1'b0};
                        wen_a20 = {1'b0, 1'b0};
                        wen_a19 = {1'b0, 1'b0};
                        wen_a18 = {1'b0, 1'b0};
                        wen_a17 = {1'b0, 1'b0};
                        wen_a16 = {1'b0, 1'b0};
                        wen_a15 = {1'b0, 1'b0};
                        wen_a14 = {1'b0, 1'b0};
                        wen_a13 = {1'b0, 1'b0};
                        wen_a12 = {1'b0, 1'b0};
                        wen_a11 = {1'b0, 1'b0};
                        wen_a10 = {1'b0, 1'b0};
                        wen_a9 = {1'b0, 1'b0};
                        wen_a8 = {1'b0, 1'b0};
                        wen_a7 = {1'b0, 1'b0};
                        wen_a6 = {1'b0, 1'b0};
                        wen_a5 = {1'b0, 1'b0};
                        wen_a4 = {1'b0, wen};
                        wen_a3 = {1'b0, wen};
                        wen_a2 = {1'b0, wen};
                        wen_a1 = {1'b0, wen};
                        wen_a0 = {1'b0, 1'b0};
                        wen_b0 = {1'b0, 1'b0};
                    end
                    5'b11100 : begin
                        wen_a28 = {1'b0, 1'b0};
                        wen_a27 = {1'b0, 1'b0};
                        wen_a26 = {1'b0, 1'b0};
                        wen_a25 = {1'b0, 1'b0};
                        wen_a24 = {1'b0, 1'b0};
                        wen_a23 = {1'b0, 1'b0};
                        wen_a22 = {1'b0, 1'b0};
                        wen_a21 = {1'b0, 1'b0};
                        wen_a20 = {1'b0, 1'b0};
                        wen_a19 = {1'b0, 1'b0};
                        wen_a18 = {1'b0, 1'b0};
                        wen_a17 = {1'b0, 1'b0};
                        wen_a16 = {1'b0, 1'b0};
                        wen_a15 = {1'b0, 1'b0};
                        wen_a14 = {1'b0, 1'b0};
                        wen_a13 = {1'b0, 1'b0};
                        wen_a12 = {1'b0, 1'b0};
                        wen_a11 = {1'b0, 1'b0};
                        wen_a10 = {1'b0, 1'b0};
                        wen_a9 = {1'b0, 1'b0};
                        wen_a8 = {1'b0, 1'b0};
                        wen_a7 = {1'b0, 1'b0};
                        wen_a6 = {1'b0, 1'b0};
                        wen_a5 = {1'b0, 1'b0};
                        wen_a4 = {1'b0, 1'b0};
                        wen_a3 = {1'b0, 1'b0};
                        wen_a2 = {1'b0, 1'b0};
                        wen_a1 = {1'b0, 1'b0};
                        wen_a0 = {wen, wen};
                        wen_b0 = {wen, wen};
                    end
                    default : begin
                        wen_a28 = {1'b0, 1'b0};
                        wen_a27 = {1'b0, 1'b0};
                        wen_a26 = {1'b0, 1'b0};
                        wen_a25 = {1'b0, 1'b0};
                        wen_a24 = {1'b0, 1'b0};
                        wen_a23 = {1'b0, 1'b0};
                        wen_a22 = {1'b0, 1'b0};
                        wen_a21 = {1'b0, 1'b0};
                        wen_a20 = {1'b0, 1'b0};
                        wen_a19 = {1'b0, 1'b0};
                        wen_a18 = {1'b0, 1'b0};
                        wen_a17 = {1'b0, 1'b0};
                        wen_a16 = {1'b0, 1'b0};
                        wen_a15 = {1'b0, 1'b0};
                        wen_a14 = {1'b0, 1'b0};
                        wen_a13 = {1'b0, 1'b0};
                        wen_a12 = {1'b0, 1'b0};
                        wen_a11 = {1'b0, 1'b0};
                        wen_a10 = {1'b0, 1'b0};
                        wen_a9 = {1'b0, 1'b0};
                        wen_a8 = {1'b0, 1'b0};
                        wen_a7 = {1'b0, 1'b0};
                        wen_a6 = {1'b0, 1'b0};
                        wen_a5 = {1'b0, 1'b0};
                        wen_a4 = {1'b0, 1'b0};
                        wen_a3 = {1'b0, 1'b0};
                        wen_a2 = {1'b0, 1'b0};
                        wen_a1 = {1'b0, 1'b0};
                        wen_a0 = {1'b0, 1'b0};
                        wen_b0 = {1'b0, 1'b0};
                    end
                endcase
                case (ckRdAddr[13:9])
                    5'b00000, 5'b00001, 5'b00010, 5'b00011,
                    5'b00100, 5'b00101, 5'b00110, 5'b00111,
                    5'b01000, 5'b01001, 5'b01010, 5'b01011,
                    5'b01100, 5'b01101, 5'b01110, 5'b01111 : begin
                        readData = {
                                        readData28[1:0],
                                        readData27[1:0],
                                        readData26[1:0],
                                        readData25[1:0],
                                        readData24[1:0],
                                        readData23[1:0],
                                        readData22[1:0],
                                        readData21[1:0],
                                        readData20[1:0],
                                        readData19[1:0],
                                        readData18[1:0],
                                        readData17[1:0],
                                        readData16[1:0],
                                        readData15[1:0],
                                        readData14[1:0],
                                        readData13[1:0]
                        };
                    end
                    5'b10000, 5'b10001, 5'b10010, 5'b10011,
                    5'b10100, 5'b10101, 5'b10110, 5'b10111 : begin
                        readData = {
                                        readData12[3:0],
                                        readData11[3:0],
                                        readData10[3:0],
                                        readData9[3:0],
                                        readData8[3:0],
                                        readData7[3:0],
                                        readData6[3:0],
                                        readData5[3:0]
                        };
                    end
                    5'b11000, 5'b11001, 5'b11010, 5'b11011 : begin
                        readData = {readData4[7:0],readData3[7:0],readData2[7:0],readData1[7:0]};
                    end
                    5'b11100 : begin
                        readData = {readData0[34:27],readData0[25:18],readData0[16:9],readData0[7:0]};
                    end
                    default : begin
                        readData = 32'b0;
                    end
                endcase
            end
            15360: begin
                width30 = 3'b001;
                width29 = 3'b001;
                width28 = 3'b001;
                width27 = 3'b001;
                width26 = 3'b001;
                width25 = 3'b001;
                width24 = 3'b001;
                width23 = 3'b001;
                width22 = 3'b001;
                width21 = 3'b001;
                width20 = 3'b001;
                width19 = 3'b001;
                width18 = 3'b001;
                width17 = 3'b001;
                width16 = 3'b001;
                width15 = 3'b001;
                width14 = 3'b010;
                width13 = 3'b010;
                width12 = 3'b010;
                width11 = 3'b010;
                width10 = 3'b010;
                width9 = 3'b010;
                width8 = 3'b010;
                width7 = 3'b010;
                width6 = 3'b011;
                width5 = 3'b011;
                width4 = 3'b011;
                width3 = 3'b011;
                width2 = 3'b100;
                width1 = 3'b100;

                writeAddr30 = {writeAddr[12:0], 1'b0};
                writeAddr29 = {writeAddr[12:0], 1'b0};
                writeAddr28 = {writeAddr[12:0], 1'b0};
                writeAddr27 = {writeAddr[12:0], 1'b0};
                writeAddr26 = {writeAddr[12:0], 1'b0};
                writeAddr25 = {writeAddr[12:0], 1'b0};
                writeAddr24 = {writeAddr[12:0], 1'b0};
                writeAddr23 = {writeAddr[12:0], 1'b0};
                writeAddr22 = {writeAddr[12:0], 1'b0};
                writeAddr21 = {writeAddr[12:0], 1'b0};
                writeAddr20 = {writeAddr[12:0], 1'b0};
                writeAddr19 = {writeAddr[12:0], 1'b0};
                writeAddr18 = {writeAddr[12:0], 1'b0};
                writeAddr17 = {writeAddr[12:0], 1'b0};
                writeAddr16 = {writeAddr[12:0], 1'b0};
                writeAddr15 = {writeAddr[12:0], 1'b0};
                writeAddr14 = {writeAddr[11:0], 2'b0};
                writeAddr13 = {writeAddr[11:0], 2'b0};
                writeAddr12 = {writeAddr[11:0], 2'b0};
                writeAddr11 = {writeAddr[11:0], 2'b0};
                writeAddr10 = {writeAddr[11:0], 2'b0};
                writeAddr9 = {writeAddr[11:0], 2'b0};
                writeAddr8 = {writeAddr[11:0], 2'b0};
                writeAddr7 = {writeAddr[11:0], 2'b0};
                writeAddr6 = {writeAddr[10:0], 3'b0};
                writeAddr5 = {writeAddr[10:0], 3'b0};
                writeAddr4 = {writeAddr[10:0], 3'b0};
                writeAddr3 = {writeAddr[10:0], 3'b0};
                writeAddr2 = {writeAddr[9:0], 4'b0};
                writeAddr1 = {writeAddr[9:0], 4'b0};

                readAddr30  = {readAddr[12:0],  1'b0};
                readAddr29  = {readAddr[12:0],  1'b0};
                readAddr28  = {readAddr[12:0],  1'b0};
                readAddr27  = {readAddr[12:0],  1'b0};
                readAddr26  = {readAddr[12:0],  1'b0};
                readAddr25  = {readAddr[12:0],  1'b0};
                readAddr24  = {readAddr[12:0],  1'b0};
                readAddr23  = {readAddr[12:0],  1'b0};
                readAddr22  = {readAddr[12:0],  1'b0};
                readAddr21  = {readAddr[12:0],  1'b0};
                readAddr20  = {readAddr[12:0],  1'b0};
                readAddr19  = {readAddr[12:0],  1'b0};
                readAddr18  = {readAddr[12:0],  1'b0};
                readAddr17  = {readAddr[12:0],  1'b0};
                readAddr16  = {readAddr[12:0],  1'b0};
                readAddr15  = {readAddr[12:0],  1'b0};
                readAddr14  = {readAddr[11:0],  2'b0};
                readAddr13  = {readAddr[11:0],  2'b0};
                readAddr12  = {readAddr[11:0],  2'b0};
                readAddr11  = {readAddr[11:0],  2'b0};
                readAddr10  = {readAddr[11:0],  2'b0};
                readAddr9  = {readAddr[11:0],  2'b0};
                readAddr8  = {readAddr[11:0],  2'b0};
                readAddr7  = {readAddr[11:0],  2'b0};
                readAddr6  = {readAddr[10:0],  3'b0};
                readAddr5  = {readAddr[10:0],  3'b0};
                readAddr4  = {readAddr[10:0],  3'b0};
                readAddr3  = {readAddr[10:0],  3'b0};
                readAddr2  = {readAddr[9:0],  4'b0};
                readAddr1  = {readAddr[9:0],  4'b0};

                writeData30 = {16'b0, writeData[31:30]};
                writeData29 = {16'b0, writeData[29:28]};
                writeData28 = {16'b0, writeData[27:26]};
                writeData27 = {16'b0, writeData[25:24]};
                writeData26 = {16'b0, writeData[23:22]};
                writeData25 = {16'b0, writeData[21:20]};
                writeData24 = {16'b0, writeData[19:18]};
                writeData23 = {16'b0, writeData[17:16]};
                writeData22 = {16'b0, writeData[15:14]};
                writeData21 = {16'b0, writeData[13:12]};
                writeData20 = {16'b0, writeData[11:10]};
                writeData19 = {16'b0, writeData[9:8]};
                writeData18 = {16'b0, writeData[7:6]};
                writeData17 = {16'b0, writeData[5:4]};
                writeData16 = {16'b0, writeData[3:2]};
                writeData15 = {16'b0, writeData[1:0]};
                writeData14 = {14'b0, writeData[31:28]};
                writeData13 = {14'b0, writeData[27:24]};
                writeData12 = {14'b0, writeData[23:20]};
                writeData11 = {14'b0, writeData[19:16]};
                writeData10 = {14'b0, writeData[15:12]};
                writeData9 = {14'b0, writeData[11:8]};
                writeData8 = {14'b0, writeData[7:4]};
                writeData7 = {14'b0, writeData[3:0]};
                writeData6 = {10'b0, writeData[31:24]};
                writeData5 = {10'b0, writeData[23:16]};
                writeData4 = {10'b0, writeData[15:8]};
                writeData3 = {10'b0, writeData[7:0]};
                writeData2 = {1'b0, writeData[31:24], 1'b0, writeData[23:16]};
                writeData1 = {1'b0, writeData[15:8], 1'b0, writeData[7:0]};

                case (writeAddr[13:9])
                    5'b00000, 5'b00001, 5'b00010, 5'b00011,
                    5'b00100, 5'b00101, 5'b00110, 5'b00111,
                    5'b01000, 5'b01001, 5'b01010, 5'b01011,
                    5'b01100, 5'b01101, 5'b01110, 5'b01111 : begin
                        wen_a30 = {1'b0, wen};
                        wen_a29 = {1'b0, wen};
                        wen_a28 = {1'b0, wen};
                        wen_a27 = {1'b0, wen};
                        wen_a26 = {1'b0, wen};
                        wen_a25 = {1'b0, wen};
                        wen_a24 = {1'b0, wen};
                        wen_a23 = {1'b0, wen};
                        wen_a22 = {1'b0, wen};
                        wen_a21 = {1'b0, wen};
                        wen_a20 = {1'b0, wen};
                        wen_a19 = {1'b0, wen};
                        wen_a18 = {1'b0, wen};
                        wen_a17 = {1'b0, wen};
                        wen_a16 = {1'b0, wen};
                        wen_a15 = {1'b0, wen};
                        wen_a14 = {1'b0, 1'b0};
                        wen_a13 = {1'b0, 1'b0};
                        wen_a12 = {1'b0, 1'b0};
                        wen_a11 = {1'b0, 1'b0};
                        wen_a10 = {1'b0, 1'b0};
                        wen_a9 = {1'b0, 1'b0};
                        wen_a8 = {1'b0, 1'b0};
                        wen_a7 = {1'b0, 1'b0};
                        wen_a6 = {1'b0, 1'b0};
                        wen_a5 = {1'b0, 1'b0};
                        wen_a4 = {1'b0, 1'b0};
                        wen_a3 = {1'b0, 1'b0};
                        wen_a2 = {1'b0, 1'b0};
                        wen_a1 = {1'b0, 1'b0};
                    end
                    5'b10000, 5'b10001, 5'b10010, 5'b10011,
                    5'b10100, 5'b10101, 5'b10110, 5'b10111 : begin
                        wen_a30 = {1'b0, 1'b0};
                        wen_a29 = {1'b0, 1'b0};
                        wen_a28 = {1'b0, 1'b0};
                        wen_a27 = {1'b0, 1'b0};
                        wen_a26 = {1'b0, 1'b0};
                        wen_a25 = {1'b0, 1'b0};
                        wen_a24 = {1'b0, 1'b0};
                        wen_a23 = {1'b0, 1'b0};
                        wen_a22 = {1'b0, 1'b0};
                        wen_a21 = {1'b0, 1'b0};
                        wen_a20 = {1'b0, 1'b0};
                        wen_a19 = {1'b0, 1'b0};
                        wen_a18 = {1'b0, 1'b0};
                        wen_a17 = {1'b0, 1'b0};
                        wen_a16 = {1'b0, 1'b0};
                        wen_a15 = {1'b0, 1'b0};
                        wen_a14 = {1'b0, wen};
                        wen_a13 = {1'b0, wen};
                        wen_a12 = {1'b0, wen};
                        wen_a11 = {1'b0, wen};
                        wen_a10 = {1'b0, wen};
                        wen_a9 = {1'b0, wen};
                        wen_a8 = {1'b0, wen};
                        wen_a7 = {1'b0, wen};
                        wen_a6 = {1'b0, 1'b0};
                        wen_a5 = {1'b0, 1'b0};
                        wen_a4 = {1'b0, 1'b0};
                        wen_a3 = {1'b0, 1'b0};
                        wen_a2 = {1'b0, 1'b0};
                        wen_a1 = {1'b0, 1'b0};
                    end
                    5'b11000, 5'b11001, 5'b11010, 5'b11011 : begin
                        wen_a30 = {1'b0, 1'b0};
                        wen_a29 = {1'b0, 1'b0};
                        wen_a28 = {1'b0, 1'b0};
                        wen_a27 = {1'b0, 1'b0};
                        wen_a26 = {1'b0, 1'b0};
                        wen_a25 = {1'b0, 1'b0};
                        wen_a24 = {1'b0, 1'b0};
                        wen_a23 = {1'b0, 1'b0};
                        wen_a22 = {1'b0, 1'b0};
                        wen_a21 = {1'b0, 1'b0};
                        wen_a20 = {1'b0, 1'b0};
                        wen_a19 = {1'b0, 1'b0};
                        wen_a18 = {1'b0, 1'b0};
                        wen_a17 = {1'b0, 1'b0};
                        wen_a16 = {1'b0, 1'b0};
                        wen_a15 = {1'b0, 1'b0};
                        wen_a14 = {1'b0, 1'b0};
                        wen_a13 = {1'b0, 1'b0};
                        wen_a12 = {1'b0, 1'b0};
                        wen_a11 = {1'b0, 1'b0};
                        wen_a10 = {1'b0, 1'b0};
                        wen_a9 = {1'b0, 1'b0};
                        wen_a8 = {1'b0, 1'b0};
                        wen_a7 = {1'b0, 1'b0};
                        wen_a6 = {1'b0, wen};
                        wen_a5 = {1'b0, wen};
                        wen_a4 = {1'b0, wen};
                        wen_a3 = {1'b0, wen};
                        wen_a2 = {1'b0, 1'b0};
                        wen_a1 = {1'b0, 1'b0};
                    end
                    5'b11100, 5'b11101 : begin
                        wen_a30 = {1'b0, 1'b0};
                        wen_a29 = {1'b0, 1'b0};
                        wen_a28 = {1'b0, 1'b0};
                        wen_a27 = {1'b0, 1'b0};
                        wen_a26 = {1'b0, 1'b0};
                        wen_a25 = {1'b0, 1'b0};
                        wen_a24 = {1'b0, 1'b0};
                        wen_a23 = {1'b0, 1'b0};
                        wen_a22 = {1'b0, 1'b0};
                        wen_a21 = {1'b0, 1'b0};
                        wen_a20 = {1'b0, 1'b0};
                        wen_a19 = {1'b0, 1'b0};
                        wen_a18 = {1'b0, 1'b0};
                        wen_a17 = {1'b0, 1'b0};
                        wen_a16 = {1'b0, 1'b0};
                        wen_a15 = {1'b0, 1'b0};
                        wen_a14 = {1'b0, 1'b0};
                        wen_a13 = {1'b0, 1'b0};
                        wen_a12 = {1'b0, 1'b0};
                        wen_a11 = {1'b0, 1'b0};
                        wen_a10 = {1'b0, 1'b0};
                        wen_a9 = {1'b0, 1'b0};
                        wen_a8 = {1'b0, 1'b0};
                        wen_a7 = {1'b0, 1'b0};
                        wen_a6 = {1'b0, 1'b0};
                        wen_a5 = {1'b0, 1'b0};
                        wen_a4 = {1'b0, 1'b0};
                        wen_a3 = {1'b0, 1'b0};
                        wen_a2 = {wen, wen};
                        wen_a1 = {wen, wen};
                    end
                    default : begin
                        wen_a30 = {1'b0, 1'b0};
                        wen_a29 = {1'b0, 1'b0};
                        wen_a28 = {1'b0, 1'b0};
                        wen_a27 = {1'b0, 1'b0};
                        wen_a26 = {1'b0, 1'b0};
                        wen_a25 = {1'b0, 1'b0};
                        wen_a24 = {1'b0, 1'b0};
                        wen_a23 = {1'b0, 1'b0};
                        wen_a22 = {1'b0, 1'b0};
                        wen_a21 = {1'b0, 1'b0};
                        wen_a20 = {1'b0, 1'b0};
                        wen_a19 = {1'b0, 1'b0};
                        wen_a18 = {1'b0, 1'b0};
                        wen_a17 = {1'b0, 1'b0};
                        wen_a16 = {1'b0, 1'b0};
                        wen_a15 = {1'b0, 1'b0};
                        wen_a14 = {1'b0, 1'b0};
                        wen_a13 = {1'b0, 1'b0};
                        wen_a12 = {1'b0, 1'b0};
                        wen_a11 = {1'b0, 1'b0};
                        wen_a10 = {1'b0, 1'b0};
                        wen_a9 = {1'b0, 1'b0};
                        wen_a8 = {1'b0, 1'b0};
                        wen_a7 = {1'b0, 1'b0};
                        wen_a6 = {1'b0, 1'b0};
                        wen_a5 = {1'b0, 1'b0};
                        wen_a4 = {1'b0, 1'b0};
                        wen_a3 = {1'b0, 1'b0};
                        wen_a2 = {1'b0, 1'b0};
                        wen_a1 = {1'b0, 1'b0};
                    end
                endcase
                case (ckRdAddr[13:9])
                    5'b00000, 5'b00001, 5'b00010, 5'b00011,
                    5'b00100, 5'b00101, 5'b00110, 5'b00111,
                    5'b01000, 5'b01001, 5'b01010, 5'b01011,
                    5'b01100, 5'b01101, 5'b01110, 5'b01111 : begin
                        readData = {
                                        readData30[1:0],
                                        readData29[1:0],
                                        readData28[1:0],
                                        readData27[1:0],
                                        readData26[1:0],
                                        readData25[1:0],
                                        readData24[1:0],
                                        readData23[1:0],
                                        readData22[1:0],
                                        readData21[1:0],
                                        readData20[1:0],
                                        readData19[1:0],
                                        readData18[1:0],
                                        readData17[1:0],
                                        readData16[1:0],
                                        readData15[1:0]
                        };
                    end
                    5'b10000, 5'b10001, 5'b10010, 5'b10011,
                    5'b10100, 5'b10101, 5'b10110, 5'b10111 : begin
                        readData = {
                                        readData14[3:0],
                                        readData13[3:0],
                                        readData12[3:0],
                                        readData11[3:0],
                                        readData10[3:0],
                                        readData9[3:0],
                                        readData8[3:0],
                                        readData7[3:0]
                        };
                    end
                    5'b11000, 5'b11001, 5'b11010, 5'b11011 : begin
                        readData = {readData6[7:0],readData5[7:0],readData4[7:0],readData3[7:0]};
                    end
                    5'b11100, 5'b11101 : begin
                        readData = {readData2[16:9],readData2[7:0],readData1[16:9],readData1[7:0]};
                    end
                    default : begin
                        readData = 32'b0;
                    end
                endcase
            end
            15872: begin
                width30 = 3'b001;
                width29 = 3'b001;
                width28 = 3'b001;
                width27 = 3'b001;
                width26 = 3'b001;
                width25 = 3'b001;
                width24 = 3'b001;
                width23 = 3'b001;
                width22 = 3'b001;
                width21 = 3'b001;
                width20 = 3'b001;
                width19 = 3'b001;
                width18 = 3'b001;
                width17 = 3'b001;
                width16 = 3'b001;
                width15 = 3'b001;
                width14 = 3'b010;
                width13 = 3'b010;
                width12 = 3'b010;
                width11 = 3'b010;
                width10 = 3'b010;
                width9 = 3'b010;
                width8 = 3'b010;
                width7 = 3'b010;
                width6 = 3'b011;
                width5 = 3'b011;
                width4 = 3'b011;
                width3 = 3'b011;
                width2 = 3'b100;
                width1 = 3'b100;
                width0 = 3'b101;

                writeAddr30 = {writeAddr[12:0], 1'b0};
                writeAddr29 = {writeAddr[12:0], 1'b0};
                writeAddr28 = {writeAddr[12:0], 1'b0};
                writeAddr27 = {writeAddr[12:0], 1'b0};
                writeAddr26 = {writeAddr[12:0], 1'b0};
                writeAddr25 = {writeAddr[12:0], 1'b0};
                writeAddr24 = {writeAddr[12:0], 1'b0};
                writeAddr23 = {writeAddr[12:0], 1'b0};
                writeAddr22 = {writeAddr[12:0], 1'b0};
                writeAddr21 = {writeAddr[12:0], 1'b0};
                writeAddr20 = {writeAddr[12:0], 1'b0};
                writeAddr19 = {writeAddr[12:0], 1'b0};
                writeAddr18 = {writeAddr[12:0], 1'b0};
                writeAddr17 = {writeAddr[12:0], 1'b0};
                writeAddr16 = {writeAddr[12:0], 1'b0};
                writeAddr15 = {writeAddr[12:0], 1'b0};
                writeAddr14 = {writeAddr[11:0], 2'b0};
                writeAddr13 = {writeAddr[11:0], 2'b0};
                writeAddr12 = {writeAddr[11:0], 2'b0};
                writeAddr11 = {writeAddr[11:0], 2'b0};
                writeAddr10 = {writeAddr[11:0], 2'b0};
                writeAddr9 = {writeAddr[11:0], 2'b0};
                writeAddr8 = {writeAddr[11:0], 2'b0};
                writeAddr7 = {writeAddr[11:0], 2'b0};
                writeAddr6 = {writeAddr[10:0], 3'b0};
                writeAddr5 = {writeAddr[10:0], 3'b0};
                writeAddr4 = {writeAddr[10:0], 3'b0};
                writeAddr3 = {writeAddr[10:0], 3'b0};
                writeAddr2 = {writeAddr[9:0], 4'b0};
                writeAddr1 = {writeAddr[9:0], 4'b0};
                writeAddr0 = {writeAddr[8:0], 5'b0};

                readAddr30  = {readAddr[12:0],  1'b0};
                readAddr29  = {readAddr[12:0],  1'b0};
                readAddr28  = {readAddr[12:0],  1'b0};
                readAddr27  = {readAddr[12:0],  1'b0};
                readAddr26  = {readAddr[12:0],  1'b0};
                readAddr25  = {readAddr[12:0],  1'b0};
                readAddr24  = {readAddr[12:0],  1'b0};
                readAddr23  = {readAddr[12:0],  1'b0};
                readAddr22  = {readAddr[12:0],  1'b0};
                readAddr21  = {readAddr[12:0],  1'b0};
                readAddr20  = {readAddr[12:0],  1'b0};
                readAddr19  = {readAddr[12:0],  1'b0};
                readAddr18  = {readAddr[12:0],  1'b0};
                readAddr17  = {readAddr[12:0],  1'b0};
                readAddr16  = {readAddr[12:0],  1'b0};
                readAddr15  = {readAddr[12:0],  1'b0};
                readAddr14  = {readAddr[11:0],  2'b0};
                readAddr13  = {readAddr[11:0],  2'b0};
                readAddr12  = {readAddr[11:0],  2'b0};
                readAddr11  = {readAddr[11:0],  2'b0};
                readAddr10  = {readAddr[11:0],  2'b0};
                readAddr9  = {readAddr[11:0],  2'b0};
                readAddr8  = {readAddr[11:0],  2'b0};
                readAddr7  = {readAddr[11:0],  2'b0};
                readAddr6  = {readAddr[10:0],  3'b0};
                readAddr5  = {readAddr[10:0],  3'b0};
                readAddr4  = {readAddr[10:0],  3'b0};
                readAddr3  = {readAddr[10:0],  3'b0};
                readAddr2  = {readAddr[9:0],  4'b0};
                readAddr1  = {readAddr[9:0],  4'b0};
                readAddr0  = {readAddr[8:0],  5'b0};

                writeData30 = {16'b0, writeData[31:30]};
                writeData29 = {16'b0, writeData[29:28]};
                writeData28 = {16'b0, writeData[27:26]};
                writeData27 = {16'b0, writeData[25:24]};
                writeData26 = {16'b0, writeData[23:22]};
                writeData25 = {16'b0, writeData[21:20]};
                writeData24 = {16'b0, writeData[19:18]};
                writeData23 = {16'b0, writeData[17:16]};
                writeData22 = {16'b0, writeData[15:14]};
                writeData21 = {16'b0, writeData[13:12]};
                writeData20 = {16'b0, writeData[11:10]};
                writeData19 = {16'b0, writeData[9:8]};
                writeData18 = {16'b0, writeData[7:6]};
                writeData17 = {16'b0, writeData[5:4]};
                writeData16 = {16'b0, writeData[3:2]};
                writeData15 = {16'b0, writeData[1:0]};
                writeData14 = {14'b0, writeData[31:28]};
                writeData13 = {14'b0, writeData[27:24]};
                writeData12 = {14'b0, writeData[23:20]};
                writeData11 = {14'b0, writeData[19:16]};
                writeData10 = {14'b0, writeData[15:12]};
                writeData9 = {14'b0, writeData[11:8]};
                writeData8 = {14'b0, writeData[7:4]};
                writeData7 = {14'b0, writeData[3:0]};
                writeData6 = {10'b0, writeData[31:24]};
                writeData5 = {10'b0, writeData[23:16]};
                writeData4 = {10'b0, writeData[15:8]};
                writeData3 = {10'b0, writeData[7:0]};
                writeData2 = {1'b0, writeData[31:24], 1'b0, writeData[23:16]};
                writeData1 = {1'b0, writeData[15:8], 1'b0, writeData[7:0]};
                writeData0 = {1'b0, writeData[31:24], 1'b0, writeData[23:16], 1'b0, writeData[15:8], 1'b0, writeData[7:0]};

                case (writeAddr[13:9])
                    5'b00000, 5'b00001, 5'b00010, 5'b00011,
                    5'b00100, 5'b00101, 5'b00110, 5'b00111,
                    5'b01000, 5'b01001, 5'b01010, 5'b01011,
                    5'b01100, 5'b01101, 5'b01110, 5'b01111 : begin
                        wen_a30 = {1'b0, wen};
                        wen_a29 = {1'b0, wen};
                        wen_a28 = {1'b0, wen};
                        wen_a27 = {1'b0, wen};
                        wen_a26 = {1'b0, wen};
                        wen_a25 = {1'b0, wen};
                        wen_a24 = {1'b0, wen};
                        wen_a23 = {1'b0, wen};
                        wen_a22 = {1'b0, wen};
                        wen_a21 = {1'b0, wen};
                        wen_a20 = {1'b0, wen};
                        wen_a19 = {1'b0, wen};
                        wen_a18 = {1'b0, wen};
                        wen_a17 = {1'b0, wen};
                        wen_a16 = {1'b0, wen};
                        wen_a15 = {1'b0, wen};
                        wen_a14 = {1'b0, 1'b0};
                        wen_a13 = {1'b0, 1'b0};
                        wen_a12 = {1'b0, 1'b0};
                        wen_a11 = {1'b0, 1'b0};
                        wen_a10 = {1'b0, 1'b0};
                        wen_a9 = {1'b0, 1'b0};
                        wen_a8 = {1'b0, 1'b0};
                        wen_a7 = {1'b0, 1'b0};
                        wen_a6 = {1'b0, 1'b0};
                        wen_a5 = {1'b0, 1'b0};
                        wen_a4 = {1'b0, 1'b0};
                        wen_a3 = {1'b0, 1'b0};
                        wen_a2 = {1'b0, 1'b0};
                        wen_a1 = {1'b0, 1'b0};
                        wen_a0 = {1'b0, 1'b0};
                        wen_b0 = {1'b0, 1'b0};
                    end
                    5'b10000, 5'b10001, 5'b10010, 5'b10011,
                    5'b10100, 5'b10101, 5'b10110, 5'b10111 : begin
                        wen_a30 = {1'b0, 1'b0};
                        wen_a29 = {1'b0, 1'b0};
                        wen_a28 = {1'b0, 1'b0};
                        wen_a27 = {1'b0, 1'b0};
                        wen_a26 = {1'b0, 1'b0};
                        wen_a25 = {1'b0, 1'b0};
                        wen_a24 = {1'b0, 1'b0};
                        wen_a23 = {1'b0, 1'b0};
                        wen_a22 = {1'b0, 1'b0};
                        wen_a21 = {1'b0, 1'b0};
                        wen_a20 = {1'b0, 1'b0};
                        wen_a19 = {1'b0, 1'b0};
                        wen_a18 = {1'b0, 1'b0};
                        wen_a17 = {1'b0, 1'b0};
                        wen_a16 = {1'b0, 1'b0};
                        wen_a15 = {1'b0, 1'b0};
                        wen_a14 = {1'b0, wen};
                        wen_a13 = {1'b0, wen};
                        wen_a12 = {1'b0, wen};
                        wen_a11 = {1'b0, wen};
                        wen_a10 = {1'b0, wen};
                        wen_a9 = {1'b0, wen};
                        wen_a8 = {1'b0, wen};
                        wen_a7 = {1'b0, wen};
                        wen_a6 = {1'b0, 1'b0};
                        wen_a5 = {1'b0, 1'b0};
                        wen_a4 = {1'b0, 1'b0};
                        wen_a3 = {1'b0, 1'b0};
                        wen_a2 = {1'b0, 1'b0};
                        wen_a1 = {1'b0, 1'b0};
                        wen_a0 = {1'b0, 1'b0};
                        wen_b0 = {1'b0, 1'b0};
                    end
                    5'b11000, 5'b11001, 5'b11010, 5'b11011 : begin
                        wen_a30 = {1'b0, 1'b0};
                        wen_a29 = {1'b0, 1'b0};
                        wen_a28 = {1'b0, 1'b0};
                        wen_a27 = {1'b0, 1'b0};
                        wen_a26 = {1'b0, 1'b0};
                        wen_a25 = {1'b0, 1'b0};
                        wen_a24 = {1'b0, 1'b0};
                        wen_a23 = {1'b0, 1'b0};
                        wen_a22 = {1'b0, 1'b0};
                        wen_a21 = {1'b0, 1'b0};
                        wen_a20 = {1'b0, 1'b0};
                        wen_a19 = {1'b0, 1'b0};
                        wen_a18 = {1'b0, 1'b0};
                        wen_a17 = {1'b0, 1'b0};
                        wen_a16 = {1'b0, 1'b0};
                        wen_a15 = {1'b0, 1'b0};
                        wen_a14 = {1'b0, 1'b0};
                        wen_a13 = {1'b0, 1'b0};
                        wen_a12 = {1'b0, 1'b0};
                        wen_a11 = {1'b0, 1'b0};
                        wen_a10 = {1'b0, 1'b0};
                        wen_a9 = {1'b0, 1'b0};
                        wen_a8 = {1'b0, 1'b0};
                        wen_a7 = {1'b0, 1'b0};
                        wen_a6 = {1'b0, wen};
                        wen_a5 = {1'b0, wen};
                        wen_a4 = {1'b0, wen};
                        wen_a3 = {1'b0, wen};
                        wen_a2 = {1'b0, 1'b0};
                        wen_a1 = {1'b0, 1'b0};
                        wen_a0 = {1'b0, 1'b0};
                        wen_b0 = {1'b0, 1'b0};
                    end
                    5'b11100, 5'b11101 : begin
                        wen_a30 = {1'b0, 1'b0};
                        wen_a29 = {1'b0, 1'b0};
                        wen_a28 = {1'b0, 1'b0};
                        wen_a27 = {1'b0, 1'b0};
                        wen_a26 = {1'b0, 1'b0};
                        wen_a25 = {1'b0, 1'b0};
                        wen_a24 = {1'b0, 1'b0};
                        wen_a23 = {1'b0, 1'b0};
                        wen_a22 = {1'b0, 1'b0};
                        wen_a21 = {1'b0, 1'b0};
                        wen_a20 = {1'b0, 1'b0};
                        wen_a19 = {1'b0, 1'b0};
                        wen_a18 = {1'b0, 1'b0};
                        wen_a17 = {1'b0, 1'b0};
                        wen_a16 = {1'b0, 1'b0};
                        wen_a15 = {1'b0, 1'b0};
                        wen_a14 = {1'b0, 1'b0};
                        wen_a13 = {1'b0, 1'b0};
                        wen_a12 = {1'b0, 1'b0};
                        wen_a11 = {1'b0, 1'b0};
                        wen_a10 = {1'b0, 1'b0};
                        wen_a9 = {1'b0, 1'b0};
                        wen_a8 = {1'b0, 1'b0};
                        wen_a7 = {1'b0, 1'b0};
                        wen_a6 = {1'b0, 1'b0};
                        wen_a5 = {1'b0, 1'b0};
                        wen_a4 = {1'b0, 1'b0};
                        wen_a3 = {1'b0, 1'b0};
                        wen_a2 = {wen, wen};
                        wen_a1 = {wen, wen};
                        wen_a0 = {1'b0, 1'b0};
                        wen_b0 = {1'b0, 1'b0};
                    end
                    5'b11110 : begin
                        wen_a30 = {1'b0, 1'b0};
                        wen_a29 = {1'b0, 1'b0};
                        wen_a28 = {1'b0, 1'b0};
                        wen_a27 = {1'b0, 1'b0};
                        wen_a26 = {1'b0, 1'b0};
                        wen_a25 = {1'b0, 1'b0};
                        wen_a24 = {1'b0, 1'b0};
                        wen_a23 = {1'b0, 1'b0};
                        wen_a22 = {1'b0, 1'b0};
                        wen_a21 = {1'b0, 1'b0};
                        wen_a20 = {1'b0, 1'b0};
                        wen_a19 = {1'b0, 1'b0};
                        wen_a18 = {1'b0, 1'b0};
                        wen_a17 = {1'b0, 1'b0};
                        wen_a16 = {1'b0, 1'b0};
                        wen_a15 = {1'b0, 1'b0};
                        wen_a14 = {1'b0, 1'b0};
                        wen_a13 = {1'b0, 1'b0};
                        wen_a12 = {1'b0, 1'b0};
                        wen_a11 = {1'b0, 1'b0};
                        wen_a10 = {1'b0, 1'b0};
                        wen_a9 = {1'b0, 1'b0};
                        wen_a8 = {1'b0, 1'b0};
                        wen_a7 = {1'b0, 1'b0};
                        wen_a6 = {1'b0, 1'b0};
                        wen_a5 = {1'b0, 1'b0};
                        wen_a4 = {1'b0, 1'b0};
                        wen_a3 = {1'b0, 1'b0};
                        wen_a2 = {1'b0, 1'b0};
                        wen_a1 = {1'b0, 1'b0};
                        wen_a0 = {wen, wen};
                        wen_b0 = {wen, wen};
                    end
                    default : begin
                        wen_a30 = {1'b0, 1'b0};
                        wen_a29 = {1'b0, 1'b0};
                        wen_a28 = {1'b0, 1'b0};
                        wen_a27 = {1'b0, 1'b0};
                        wen_a26 = {1'b0, 1'b0};
                        wen_a25 = {1'b0, 1'b0};
                        wen_a24 = {1'b0, 1'b0};
                        wen_a23 = {1'b0, 1'b0};
                        wen_a22 = {1'b0, 1'b0};
                        wen_a21 = {1'b0, 1'b0};
                        wen_a20 = {1'b0, 1'b0};
                        wen_a19 = {1'b0, 1'b0};
                        wen_a18 = {1'b0, 1'b0};
                        wen_a17 = {1'b0, 1'b0};
                        wen_a16 = {1'b0, 1'b0};
                        wen_a15 = {1'b0, 1'b0};
                        wen_a14 = {1'b0, 1'b0};
                        wen_a13 = {1'b0, 1'b0};
                        wen_a12 = {1'b0, 1'b0};
                        wen_a11 = {1'b0, 1'b0};
                        wen_a10 = {1'b0, 1'b0};
                        wen_a9 = {1'b0, 1'b0};
                        wen_a8 = {1'b0, 1'b0};
                        wen_a7 = {1'b0, 1'b0};
                        wen_a6 = {1'b0, 1'b0};
                        wen_a5 = {1'b0, 1'b0};
                        wen_a4 = {1'b0, 1'b0};
                        wen_a3 = {1'b0, 1'b0};
                        wen_a2 = {1'b0, 1'b0};
                        wen_a1 = {1'b0, 1'b0};
                        wen_a0 = {1'b0, 1'b0};
                        wen_b0 = {1'b0, 1'b0};
                    end
                endcase
                case (ckRdAddr[13:9])
                    5'b00000, 5'b00001, 5'b00010, 5'b00011,
                    5'b00100, 5'b00101, 5'b00110, 5'b00111,
                    5'b01000, 5'b01001, 5'b01010, 5'b01011,
                    5'b01100, 5'b01101, 5'b01110, 5'b01111 : begin
                        readData = {
                                        readData30[1:0],
                                        readData29[1:0],
                                        readData28[1:0],
                                        readData27[1:0],
                                        readData26[1:0],
                                        readData25[1:0],
                                        readData24[1:0],
                                        readData23[1:0],
                                        readData22[1:0],
                                        readData21[1:0],
                                        readData20[1:0],
                                        readData19[1:0],
                                        readData18[1:0],
                                        readData17[1:0],
                                        readData16[1:0],
                                        readData15[1:0]
                        };
                    end
                    5'b10000, 5'b10001, 5'b10010, 5'b10011,
                    5'b10100, 5'b10101, 5'b10110, 5'b10111 : begin
                        readData = {
                                        readData14[3:0],
                                        readData13[3:0],
                                        readData12[3:0],
                                        readData11[3:0],
                                        readData10[3:0],
                                        readData9[3:0],
                                        readData8[3:0],
                                        readData7[3:0]
                        };
                    end
                    5'b11000, 5'b11001, 5'b11010, 5'b11011 : begin
                        readData = {readData6[7:0],readData5[7:0],readData4[7:0],readData3[7:0]};
                    end
                    5'b11100, 5'b11101 : begin
                        readData = {readData2[16:9],readData2[7:0],readData1[16:9],readData1[7:0]};
                    end
                    5'b11110 : begin
                        readData = {readData0[34:27],readData0[25:18],readData0[16:9],readData0[7:0]};
                    end
                    default : begin
                        readData = 32'b0;
                    end
                endcase
            end
            16384: begin
                width32 = 3'b000;
                width31 = 3'b000;
                width30 = 3'b000;
                width29 = 3'b000;
                width28 = 3'b000;
                width27 = 3'b000;
                width26 = 3'b000;
                width25 = 3'b000;
                width24 = 3'b000;
                width23 = 3'b000;
                width22 = 3'b000;
                width21 = 3'b000;
                width20 = 3'b000;
                width19 = 3'b000;
                width18 = 3'b000;
                width17 = 3'b000;
                width16 = 3'b000;
                width15 = 3'b000;
                width14 = 3'b000;
                width13 = 3'b000;
                width12 = 3'b000;
                width11 = 3'b000;
                width10 = 3'b000;
                width9 = 3'b000;
                width8 = 3'b000;
                width7 = 3'b000;
                width6 = 3'b000;
                width5 = 3'b000;
                width4 = 3'b000;
                width3 = 3'b000;
                width2 = 3'b000;
                width1 = 3'b000;

                writeAddr32 = {writeAddr[13:0]};
                writeAddr31 = {writeAddr[13:0]};
                writeAddr30 = {writeAddr[13:0]};
                writeAddr29 = {writeAddr[13:0]};
                writeAddr28 = {writeAddr[13:0]};
                writeAddr27 = {writeAddr[13:0]};
                writeAddr26 = {writeAddr[13:0]};
                writeAddr25 = {writeAddr[13:0]};
                writeAddr24 = {writeAddr[13:0]};
                writeAddr23 = {writeAddr[13:0]};
                writeAddr22 = {writeAddr[13:0]};
                writeAddr21 = {writeAddr[13:0]};
                writeAddr20 = {writeAddr[13:0]};
                writeAddr19 = {writeAddr[13:0]};
                writeAddr18 = {writeAddr[13:0]};
                writeAddr17 = {writeAddr[13:0]};
                writeAddr16 = {writeAddr[13:0]};
                writeAddr15 = {writeAddr[13:0]};
                writeAddr14 = {writeAddr[13:0]};
                writeAddr13 = {writeAddr[13:0]};
                writeAddr12 = {writeAddr[13:0]};
                writeAddr11 = {writeAddr[13:0]};
                writeAddr10 = {writeAddr[13:0]};
                writeAddr9 = {writeAddr[13:0]};
                writeAddr8 = {writeAddr[13:0]};
                writeAddr7 = {writeAddr[13:0]};
                writeAddr6 = {writeAddr[13:0]};
                writeAddr5 = {writeAddr[13:0]};
                writeAddr4 = {writeAddr[13:0]};
                writeAddr3 = {writeAddr[13:0]};
                writeAddr2 = {writeAddr[13:0]};
                writeAddr1 = {writeAddr[13:0]};

                readAddr32 = {writeAddr[13:0]};
                readAddr31 = {writeAddr[13:0]};
                readAddr30 = {writeAddr[13:0]};
                readAddr29 = {writeAddr[13:0]};
                readAddr28 = {writeAddr[13:0]};
                readAddr27 = {writeAddr[13:0]};
                readAddr26 = {writeAddr[13:0]};
                readAddr25 = {writeAddr[13:0]};
                readAddr24 = {writeAddr[13:0]};
                readAddr23 = {writeAddr[13:0]};
                readAddr22 = {writeAddr[13:0]};
                readAddr21 = {writeAddr[13:0]};
                readAddr20 = {writeAddr[13:0]};
                readAddr19 = {writeAddr[13:0]};
                readAddr18 = {writeAddr[13:0]};
                readAddr17 = {writeAddr[13:0]};
                readAddr16 = {writeAddr[13:0]};
                readAddr15 = {writeAddr[13:0]};
                readAddr14 = {writeAddr[13:0]};
                readAddr13 = {writeAddr[13:0]};
                readAddr12 = {writeAddr[13:0]};
                readAddr11 = {writeAddr[13:0]};
                readAddr10 = {writeAddr[13:0]};
                readAddr9 = {writeAddr[13:0]};
                readAddr8 = {writeAddr[13:0]};
                readAddr7 = {writeAddr[13:0]};
                readAddr6 = {writeAddr[13:0]};
                readAddr5 = {writeAddr[13:0]};
                readAddr4 = {writeAddr[13:0]};
                readAddr3 = {writeAddr[13:0]};
                readAddr2 = {writeAddr[13:0]};
                readAddr1 = {writeAddr[13:0]};

                writeData32 = {17'b0, writeData[31]};
                writeData31 = {17'b0, writeData[30]};
                writeData30 = {17'b0, writeData[29]};
                writeData29 = {17'b0, writeData[28]};
                writeData28 = {17'b0, writeData[27]};
                writeData27 = {17'b0, writeData[26]};
                writeData26 = {17'b0, writeData[25]};
                writeData25 = {17'b0, writeData[24]};
                writeData24 = {17'b0, writeData[23]};
                writeData23 = {17'b0, writeData[22]};
                writeData22 = {17'b0, writeData[21]};
                writeData21 = {17'b0, writeData[20]};
                writeData20 = {17'b0, writeData[19]};
                writeData19 = {17'b0, writeData[18]};
                writeData18 = {17'b0, writeData[17]};
                writeData17 = {17'b0, writeData[16]};
                writeData16 = {17'b0, writeData[15]};
                writeData15 = {17'b0, writeData[14]};
                writeData14 = {17'b0, writeData[13]};
                writeData13 = {17'b0, writeData[12]};
                writeData12 = {17'b0, writeData[11]};
                writeData11 = {17'b0, writeData[10]};
                writeData10 = {17'b0, writeData[9]};
                writeData9 = {17'b0, writeData[8]};
                writeData8 = {17'b0, writeData[7]};
                writeData7 = {17'b0, writeData[6]};
                writeData6 = {17'b0, writeData[5]};
                writeData5 = {17'b0, writeData[4]};
                writeData4 = {17'b0, writeData[3]};
                writeData3 = {17'b0, writeData[2]};
                writeData2 = {17'b0, writeData[1]};
                writeData1 = {17'b0, writeData[0]};

                wen_a32 = {1'b0, wen};
                wen_a31 = {1'b0, wen};
                wen_a30 = {1'b0, wen};
                wen_a29 = {1'b0, wen};
                wen_a28 = {1'b0, wen};
                wen_a27 = {1'b0, wen};
                wen_a26 = {1'b0, wen};
                wen_a25 = {1'b0, wen};
                wen_a24 = {1'b0, wen};
                wen_a23 = {1'b0, wen};
                wen_a22 = {1'b0, wen};
                wen_a21 = {1'b0, wen};
                wen_a20 = {1'b0, wen};
                wen_a19 = {1'b0, wen};
                wen_a18 = {1'b0, wen};
                wen_a17 = {1'b0, wen};
                wen_a16 = {1'b0, wen};
                wen_a15 = {1'b0, wen};
                wen_a14 = {1'b0, wen};
                wen_a13 = {1'b0, wen};
                wen_a12 = {1'b0, wen};
                wen_a11 = {1'b0, wen};
                wen_a10 = {1'b0, wen};
                wen_a9 = {1'b0, wen};
                wen_a8 = {1'b0, wen};
                wen_a7 = {1'b0, wen};
                wen_a6 = {1'b0, wen};
                wen_a5 = {1'b0, wen};
                wen_a4 = {1'b0, wen};
                wen_a3 = {1'b0, wen};
                wen_a2 = {1'b0, wen};
                wen_a1 = {1'b0, wen};

                readData = {
                                readData32[0],
                                readData31[0],
                                readData30[0],
                                readData29[0],
                                readData28[0],
                                readData27[0],
                                readData26[0],
                                readData25[0],
                                readData24[0],
                                readData23[0],
                                readData22[0],
                                readData21[0],
                                readData20[0],
                                readData19[0],
                                readData18[0],
                                readData17[0],
                                readData16[0],
                                readData15[0],
                                readData14[0],
                                readData13[0],
                                readData12[0],
                                readData11[0],
                                readData10[0],
                                readData9[0],
                                readData8[0],
                                readData7[0],
                                readData6[0],
                                readData5[0],
                                readData4[0],
                                readData3[0],
                                readData2[0],
                                readData1[0]
                };
            end
            16896: begin
                width32 = 3'b000;
                width31 = 3'b000;
                width30 = 3'b000;
                width29 = 3'b000;
                width28 = 3'b000;
                width27 = 3'b000;
                width26 = 3'b000;
                width25 = 3'b000;
                width24 = 3'b000;
                width23 = 3'b000;
                width22 = 3'b000;
                width21 = 3'b000;
                width20 = 3'b000;
                width19 = 3'b000;
                width18 = 3'b000;
                width17 = 3'b000;
                width16 = 3'b000;
                width15 = 3'b000;
                width14 = 3'b000;
                width13 = 3'b000;
                width12 = 3'b000;
                width11 = 3'b000;
                width10 = 3'b000;
                width9 = 3'b000;
                width8 = 3'b000;
                width7 = 3'b000;
                width6 = 3'b000;
                width5 = 3'b000;
                width4 = 3'b000;
                width3 = 3'b000;
                width2 = 3'b000;
                width1 = 3'b000;
                width0 = 3'b101;

                writeAddr32 = {writeAddr[13:0]};
                writeAddr31 = {writeAddr[13:0]};
                writeAddr30 = {writeAddr[13:0]};
                writeAddr29 = {writeAddr[13:0]};
                writeAddr28 = {writeAddr[13:0]};
                writeAddr27 = {writeAddr[13:0]};
                writeAddr26 = {writeAddr[13:0]};
                writeAddr25 = {writeAddr[13:0]};
                writeAddr24 = {writeAddr[13:0]};
                writeAddr23 = {writeAddr[13:0]};
                writeAddr22 = {writeAddr[13:0]};
                writeAddr21 = {writeAddr[13:0]};
                writeAddr20 = {writeAddr[13:0]};
                writeAddr19 = {writeAddr[13:0]};
                writeAddr18 = {writeAddr[13:0]};
                writeAddr17 = {writeAddr[13:0]};
                writeAddr16 = {writeAddr[13:0]};
                writeAddr15 = {writeAddr[13:0]};
                writeAddr14 = {writeAddr[13:0]};
                writeAddr13 = {writeAddr[13:0]};
                writeAddr12 = {writeAddr[13:0]};
                writeAddr11 = {writeAddr[13:0]};
                writeAddr10 = {writeAddr[13:0]};
                writeAddr9 = {writeAddr[13:0]};
                writeAddr8 = {writeAddr[13:0]};
                writeAddr7 = {writeAddr[13:0]};
                writeAddr6 = {writeAddr[13:0]};
                writeAddr5 = {writeAddr[13:0]};
                writeAddr4 = {writeAddr[13:0]};
                writeAddr3 = {writeAddr[13:0]};
                writeAddr2 = {writeAddr[13:0]};
                writeAddr1 = {writeAddr[13:0]};
                writeAddr0 = {writeAddr[8:0], 5'b0};

                readAddr32 = {writeAddr[13:0]};
                readAddr31 = {writeAddr[13:0]};
                readAddr30 = {writeAddr[13:0]};
                readAddr29 = {writeAddr[13:0]};
                readAddr28 = {writeAddr[13:0]};
                readAddr27 = {writeAddr[13:0]};
                readAddr26 = {writeAddr[13:0]};
                readAddr25 = {writeAddr[13:0]};
                readAddr24 = {writeAddr[13:0]};
                readAddr23 = {writeAddr[13:0]};
                readAddr22 = {writeAddr[13:0]};
                readAddr21 = {writeAddr[13:0]};
                readAddr20 = {writeAddr[13:0]};
                readAddr19 = {writeAddr[13:0]};
                readAddr18 = {writeAddr[13:0]};
                readAddr17 = {writeAddr[13:0]};
                readAddr16 = {writeAddr[13:0]};
                readAddr15 = {writeAddr[13:0]};
                readAddr14 = {writeAddr[13:0]};
                readAddr13 = {writeAddr[13:0]};
                readAddr12 = {writeAddr[13:0]};
                readAddr11 = {writeAddr[13:0]};
                readAddr10 = {writeAddr[13:0]};
                readAddr9 = {writeAddr[13:0]};
                readAddr8 = {writeAddr[13:0]};
                readAddr7 = {writeAddr[13:0]};
                readAddr6 = {writeAddr[13:0]};
                readAddr5 = {writeAddr[13:0]};
                readAddr4 = {writeAddr[13:0]};
                readAddr3 = {writeAddr[13:0]};
                readAddr2 = {writeAddr[13:0]};
                readAddr1 = {writeAddr[13:0]};
                readAddr0  = {readAddr[8:0],  5'b0};

                writeData32 = {17'b0, writeData[31]};
                writeData31 = {17'b0, writeData[30]};
                writeData30 = {17'b0, writeData[29]};
                writeData29 = {17'b0, writeData[28]};
                writeData28 = {17'b0, writeData[27]};
                writeData27 = {17'b0, writeData[26]};
                writeData26 = {17'b0, writeData[25]};
                writeData25 = {17'b0, writeData[24]};
                writeData24 = {17'b0, writeData[23]};
                writeData23 = {17'b0, writeData[22]};
                writeData22 = {17'b0, writeData[21]};
                writeData21 = {17'b0, writeData[20]};
                writeData20 = {17'b0, writeData[19]};
                writeData19 = {17'b0, writeData[18]};
                writeData18 = {17'b0, writeData[17]};
                writeData17 = {17'b0, writeData[16]};
                writeData16 = {17'b0, writeData[15]};
                writeData15 = {17'b0, writeData[14]};
                writeData14 = {17'b0, writeData[13]};
                writeData13 = {17'b0, writeData[12]};
                writeData12 = {17'b0, writeData[11]};
                writeData11 = {17'b0, writeData[10]};
                writeData10 = {17'b0, writeData[9]};
                writeData9 = {17'b0, writeData[8]};
                writeData8 = {17'b0, writeData[7]};
                writeData7 = {17'b0, writeData[6]};
                writeData6 = {17'b0, writeData[5]};
                writeData5 = {17'b0, writeData[4]};
                writeData4 = {17'b0, writeData[3]};
                writeData3 = {17'b0, writeData[2]};
                writeData2 = {17'b0, writeData[1]};
                writeData1 = {17'b0, writeData[0]};
                writeData0 = {1'b0, writeData[31:24], 1'b0, writeData[23:16], 1'b0, writeData[15:8], 1'b0, writeData[7:0]};

                case (writeAddr[14:9])
                    6'b000000, 6'b000001, 6'b000010, 6'b000011,
                    6'b000100, 6'b000101, 6'b000110, 6'b000111,
                    6'b001000, 6'b001001, 6'b001010, 6'b001011,
                    6'b001100, 6'b001101, 6'b001110, 6'b001111,
                    6'b010000, 6'b010001, 6'b010010, 6'b010011,
                    6'b010100, 6'b010101, 6'b010110, 6'b010111,
                    6'b011000, 6'b011001, 6'b011010, 6'b011011,
                    6'b011100, 6'b011101, 6'b011110, 6'b011111 : begin
                        wen_a32 = {1'b0, wen};
                        wen_a31 = {1'b0, wen};
                        wen_a30 = {1'b0, wen};
                        wen_a29 = {1'b0, wen};
                        wen_a28 = {1'b0, wen};
                        wen_a27 = {1'b0, wen};
                        wen_a26 = {1'b0, wen};
                        wen_a25 = {1'b0, wen};
                        wen_a24 = {1'b0, wen};
                        wen_a23 = {1'b0, wen};
                        wen_a22 = {1'b0, wen};
                        wen_a21 = {1'b0, wen};
                        wen_a20 = {1'b0, wen};
                        wen_a19 = {1'b0, wen};
                        wen_a18 = {1'b0, wen};
                        wen_a17 = {1'b0, wen};
                        wen_a16 = {1'b0, wen};
                        wen_a15 = {1'b0, wen};
                        wen_a14 = {1'b0, wen};
                        wen_a13 = {1'b0, wen};
                        wen_a12 = {1'b0, wen};
                        wen_a11 = {1'b0, wen};
                        wen_a10 = {1'b0, wen};
                        wen_a9 = {1'b0, wen};
                        wen_a8 = {1'b0, wen};
                        wen_a7 = {1'b0, wen};
                        wen_a6 = {1'b0, wen};
                        wen_a5 = {1'b0, wen};
                        wen_a4 = {1'b0, wen};
                        wen_a3 = {1'b0, wen};
                        wen_a2 = {1'b0, wen};
                        wen_a1 = {1'b0, wen};
                        wen_a0 = {1'b0, 1'b0};
                        wen_b0 = {1'b0, 1'b0};
                    end
                    6'b100000 : begin
                        wen_a32 = {1'b0, 1'b0};
                        wen_a31 = {1'b0, 1'b0};
                        wen_a30 = {1'b0, 1'b0};
                        wen_a29 = {1'b0, 1'b0};
                        wen_a28 = {1'b0, 1'b0};
                        wen_a27 = {1'b0, 1'b0};
                        wen_a26 = {1'b0, 1'b0};
                        wen_a25 = {1'b0, 1'b0};
                        wen_a24 = {1'b0, 1'b0};
                        wen_a23 = {1'b0, 1'b0};
                        wen_a22 = {1'b0, 1'b0};
                        wen_a21 = {1'b0, 1'b0};
                        wen_a20 = {1'b0, 1'b0};
                        wen_a19 = {1'b0, 1'b0};
                        wen_a18 = {1'b0, 1'b0};
                        wen_a17 = {1'b0, 1'b0};
                        wen_a16 = {1'b0, 1'b0};
                        wen_a15 = {1'b0, 1'b0};
                        wen_a14 = {1'b0, 1'b0};
                        wen_a13 = {1'b0, 1'b0};
                        wen_a12 = {1'b0, 1'b0};
                        wen_a11 = {1'b0, 1'b0};
                        wen_a10 = {1'b0, 1'b0};
                        wen_a9 = {1'b0, 1'b0};
                        wen_a8 = {1'b0, 1'b0};
                        wen_a7 = {1'b0, 1'b0};
                        wen_a6 = {1'b0, 1'b0};
                        wen_a5 = {1'b0, 1'b0};
                        wen_a4 = {1'b0, 1'b0};
                        wen_a3 = {1'b0, 1'b0};
                        wen_a2 = {1'b0, 1'b0};
                        wen_a1 = {1'b0, 1'b0};
                        wen_a0 = {wen, wen};
                        wen_b0 = {wen, wen};
                    end
                    default : begin
                        wen_a32 = {1'b0, 1'b0};
                        wen_a31 = {1'b0, 1'b0};
                        wen_a30 = {1'b0, 1'b0};
                        wen_a29 = {1'b0, 1'b0};
                        wen_a28 = {1'b0, 1'b0};
                        wen_a27 = {1'b0, 1'b0};
                        wen_a26 = {1'b0, 1'b0};
                        wen_a25 = {1'b0, 1'b0};
                        wen_a24 = {1'b0, 1'b0};
                        wen_a23 = {1'b0, 1'b0};
                        wen_a22 = {1'b0, 1'b0};
                        wen_a21 = {1'b0, 1'b0};
                        wen_a20 = {1'b0, 1'b0};
                        wen_a19 = {1'b0, 1'b0};
                        wen_a18 = {1'b0, 1'b0};
                        wen_a17 = {1'b0, 1'b0};
                        wen_a16 = {1'b0, 1'b0};
                        wen_a15 = {1'b0, 1'b0};
                        wen_a14 = {1'b0, 1'b0};
                        wen_a13 = {1'b0, 1'b0};
                        wen_a12 = {1'b0, 1'b0};
                        wen_a11 = {1'b0, 1'b0};
                        wen_a10 = {1'b0, 1'b0};
                        wen_a9 = {1'b0, 1'b0};
                        wen_a8 = {1'b0, 1'b0};
                        wen_a7 = {1'b0, 1'b0};
                        wen_a6 = {1'b0, 1'b0};
                        wen_a5 = {1'b0, 1'b0};
                        wen_a4 = {1'b0, 1'b0};
                        wen_a3 = {1'b0, 1'b0};
                        wen_a2 = {1'b0, 1'b0};
                        wen_a1 = {1'b0, 1'b0};
                        wen_a0 = {1'b0, 1'b0};
                        wen_b0 = {1'b0, 1'b0};
                    end
                endcase

                case (ckRdAddr[14:9])
                    6'b000000, 6'b000001, 6'b000010, 6'b000011,
                    6'b000100, 6'b000101, 6'b000110, 6'b000111,
                    6'b001000, 6'b001001, 6'b001010, 6'b001011,
                    6'b001100, 6'b001101, 6'b001110, 6'b001111,
                    6'b010000, 6'b010001, 6'b010010, 6'b010011,
                    6'b010100, 6'b010101, 6'b010110, 6'b010111,
                    6'b011000, 6'b011001, 6'b011010, 6'b011011,
                    6'b011100, 6'b011101, 6'b011110, 6'b011111 : begin
                        readData = {
                                        readData32[0],
                                        readData31[0],
                                        readData30[0],
                                        readData29[0],
                                        readData28[0],
                                        readData27[0],
                                        readData26[0],
                                        readData25[0],
                                        readData24[0],
                                        readData23[0],
                                        readData22[0],
                                        readData21[0],
                                        readData20[0],
                                        readData19[0],
                                        readData18[0],
                                        readData17[0],
                                        readData16[0],
                                        readData15[0],
                                        readData14[0],
                                        readData13[0],
                                        readData12[0],
                                        readData11[0],
                                        readData10[0],
                                        readData9[0],
                                        readData8[0],
                                        readData7[0],
                                        readData6[0],
                                        readData5[0],
                                        readData4[0],
                                        readData3[0],
                                        readData2[0],
                                        readData1[0]
                        };
                    end
                    6'b100000 : begin
                        readData = {readData0[34:27],readData0[25:18],readData0[16:9],readData0[7:0]};
                    end
                    default : begin
                        readData = 32'b0;
                    end
                endcase
            end
            17408: begin
                width34 = 3'b000;
                width33 = 3'b000;
                width32 = 3'b000;
                width31 = 3'b000;
                width30 = 3'b000;
                width29 = 3'b000;
                width28 = 3'b000;
                width27 = 3'b000;
                width26 = 3'b000;
                width25 = 3'b000;
                width24 = 3'b000;
                width23 = 3'b000;
                width22 = 3'b000;
                width21 = 3'b000;
                width20 = 3'b000;
                width19 = 3'b000;
                width18 = 3'b000;
                width17 = 3'b000;
                width16 = 3'b000;
                width15 = 3'b000;
                width14 = 3'b000;
                width13 = 3'b000;
                width12 = 3'b000;
                width11 = 3'b000;
                width10 = 3'b000;
                width9 = 3'b000;
                width8 = 3'b000;
                width7 = 3'b000;
                width6 = 3'b000;
                width5 = 3'b000;
                width4 = 3'b000;
                width3 = 3'b000;
                width2 = 3'b100;
                width1 = 3'b100;

                writeAddr34 = {writeAddr[13:0]};
                writeAddr33 = {writeAddr[13:0]};
                writeAddr32 = {writeAddr[13:0]};
                writeAddr31 = {writeAddr[13:0]};
                writeAddr30 = {writeAddr[13:0]};
                writeAddr29 = {writeAddr[13:0]};
                writeAddr28 = {writeAddr[13:0]};
                writeAddr27 = {writeAddr[13:0]};
                writeAddr26 = {writeAddr[13:0]};
                writeAddr25 = {writeAddr[13:0]};
                writeAddr24 = {writeAddr[13:0]};
                writeAddr23 = {writeAddr[13:0]};
                writeAddr22 = {writeAddr[13:0]};
                writeAddr21 = {writeAddr[13:0]};
                writeAddr20 = {writeAddr[13:0]};
                writeAddr19 = {writeAddr[13:0]};
                writeAddr18 = {writeAddr[13:0]};
                writeAddr17 = {writeAddr[13:0]};
                writeAddr16 = {writeAddr[13:0]};
                writeAddr15 = {writeAddr[13:0]};
                writeAddr14 = {writeAddr[13:0]};
                writeAddr13 = {writeAddr[13:0]};
                writeAddr12 = {writeAddr[13:0]};
                writeAddr11 = {writeAddr[13:0]};
                writeAddr10 = {writeAddr[13:0]};
                writeAddr9 = {writeAddr[13:0]};
                writeAddr8 = {writeAddr[13:0]};
                writeAddr7 = {writeAddr[13:0]};
                writeAddr6 = {writeAddr[13:0]};
                writeAddr5 = {writeAddr[13:0]};
                writeAddr4 = {writeAddr[13:0]};
                writeAddr3 = {writeAddr[13:0]};
                writeAddr2 = {writeAddr[9:0], 4'b0};
                writeAddr1 = {writeAddr[9:0], 4'b0};

                readAddr34 = {writeAddr[13:0]};
                readAddr33 = {writeAddr[13:0]};
                readAddr32 = {writeAddr[13:0]};
                readAddr31 = {writeAddr[13:0]};
                readAddr30 = {writeAddr[13:0]};
                readAddr29 = {writeAddr[13:0]};
                readAddr28 = {writeAddr[13:0]};
                readAddr27 = {writeAddr[13:0]};
                readAddr26 = {writeAddr[13:0]};
                readAddr25 = {writeAddr[13:0]};
                readAddr24 = {writeAddr[13:0]};
                readAddr23 = {writeAddr[13:0]};
                readAddr22 = {writeAddr[13:0]};
                readAddr21 = {writeAddr[13:0]};
                readAddr20 = {writeAddr[13:0]};
                readAddr19 = {writeAddr[13:0]};
                readAddr18 = {writeAddr[13:0]};
                readAddr17 = {writeAddr[13:0]};
                readAddr16 = {writeAddr[13:0]};
                readAddr15 = {writeAddr[13:0]};
                readAddr14 = {writeAddr[13:0]};
                readAddr13 = {writeAddr[13:0]};
                readAddr12 = {writeAddr[13:0]};
                readAddr11 = {writeAddr[13:0]};
                readAddr10 = {writeAddr[13:0]};
                readAddr9 = {writeAddr[13:0]};
                readAddr8 = {writeAddr[13:0]};
                readAddr7 = {writeAddr[13:0]};
                readAddr6 = {writeAddr[13:0]};
                readAddr5 = {writeAddr[13:0]};
                readAddr4 = {writeAddr[13:0]};
                readAddr3 = {writeAddr[13:0]};
                readAddr2  = {readAddr[9:0],  4'b0};
                readAddr1  = {readAddr[9:0],  4'b0};

                writeData34 = {17'b0, writeData[31]};
                writeData33 = {17'b0, writeData[30]};
                writeData32 = {17'b0, writeData[29]};
                writeData31 = {17'b0, writeData[28]};
                writeData30 = {17'b0, writeData[27]};
                writeData29 = {17'b0, writeData[26]};
                writeData28 = {17'b0, writeData[25]};
                writeData27 = {17'b0, writeData[24]};
                writeData26 = {17'b0, writeData[23]};
                writeData25 = {17'b0, writeData[22]};
                writeData24 = {17'b0, writeData[21]};
                writeData23 = {17'b0, writeData[20]};
                writeData22 = {17'b0, writeData[19]};
                writeData21 = {17'b0, writeData[18]};
                writeData20 = {17'b0, writeData[17]};
                writeData19 = {17'b0, writeData[16]};
                writeData18 = {17'b0, writeData[15]};
                writeData17 = {17'b0, writeData[14]};
                writeData16 = {17'b0, writeData[13]};
                writeData15 = {17'b0, writeData[12]};
                writeData14 = {17'b0, writeData[11]};
                writeData13 = {17'b0, writeData[10]};
                writeData12 = {17'b0, writeData[9]};
                writeData11 = {17'b0, writeData[8]};
                writeData10 = {17'b0, writeData[7]};
                writeData9 = {17'b0, writeData[6]};
                writeData8 = {17'b0, writeData[5]};
                writeData7 = {17'b0, writeData[4]};
                writeData6 = {17'b0, writeData[3]};
                writeData5 = {17'b0, writeData[2]};
                writeData4 = {17'b0, writeData[1]};
                writeData3 = {17'b0, writeData[0]};
                writeData2 = {1'b0, writeData[31:24], 1'b0, writeData[23:16]};
                writeData1 = {1'b0, writeData[15:8], 1'b0, writeData[7:0]};

                case (writeAddr[14:9])
                    6'b000000, 6'b000001, 6'b000010, 6'b000011,
                    6'b000100, 6'b000101, 6'b000110, 6'b000111,
                    6'b001000, 6'b001001, 6'b001010, 6'b001011,
                    6'b001100, 6'b001101, 6'b001110, 6'b001111,
                    6'b010000, 6'b010001, 6'b010010, 6'b010011,
                    6'b010100, 6'b010101, 6'b010110, 6'b010111,
                    6'b011000, 6'b011001, 6'b011010, 6'b011011,
                    6'b011100, 6'b011101, 6'b011110, 6'b011111 : begin
                        wen_a34 = {1'b0, wen};
                        wen_a33 = {1'b0, wen};
                        wen_a32 = {1'b0, wen};
                        wen_a31 = {1'b0, wen};
                        wen_a30 = {1'b0, wen};
                        wen_a29 = {1'b0, wen};
                        wen_a28 = {1'b0, wen};
                        wen_a27 = {1'b0, wen};
                        wen_a26 = {1'b0, wen};
                        wen_a25 = {1'b0, wen};
                        wen_a24 = {1'b0, wen};
                        wen_a23 = {1'b0, wen};
                        wen_a22 = {1'b0, wen};
                        wen_a21 = {1'b0, wen};
                        wen_a20 = {1'b0, wen};
                        wen_a19 = {1'b0, wen};
                        wen_a18 = {1'b0, wen};
                        wen_a17 = {1'b0, wen};
                        wen_a16 = {1'b0, wen};
                        wen_a15 = {1'b0, wen};
                        wen_a14 = {1'b0, wen};
                        wen_a13 = {1'b0, wen};
                        wen_a12 = {1'b0, wen};
                        wen_a11 = {1'b0, wen};
                        wen_a10 = {1'b0, wen};
                        wen_a9 = {1'b0, wen};
                        wen_a8 = {1'b0, wen};
                        wen_a7 = {1'b0, wen};
                        wen_a6 = {1'b0, wen};
                        wen_a5 = {1'b0, wen};
                        wen_a4 = {1'b0, wen};
                        wen_a3 = {1'b0, wen};
                        wen_a2 = {1'b0, 1'b0};
                        wen_a1 = {1'b0, 1'b0};
                    end
                    6'b100000, 6'b100001 : begin
                        wen_a34 = {1'b0, 1'b0};
                        wen_a33 = {1'b0, 1'b0};
                        wen_a32 = {1'b0, 1'b0};
                        wen_a31 = {1'b0, 1'b0};
                        wen_a30 = {1'b0, 1'b0};
                        wen_a29 = {1'b0, 1'b0};
                        wen_a28 = {1'b0, 1'b0};
                        wen_a27 = {1'b0, 1'b0};
                        wen_a26 = {1'b0, 1'b0};
                        wen_a25 = {1'b0, 1'b0};
                        wen_a24 = {1'b0, 1'b0};
                        wen_a23 = {1'b0, 1'b0};
                        wen_a22 = {1'b0, 1'b0};
                        wen_a21 = {1'b0, 1'b0};
                        wen_a20 = {1'b0, 1'b0};
                        wen_a19 = {1'b0, 1'b0};
                        wen_a18 = {1'b0, 1'b0};
                        wen_a17 = {1'b0, 1'b0};
                        wen_a16 = {1'b0, 1'b0};
                        wen_a15 = {1'b0, 1'b0};
                        wen_a14 = {1'b0, 1'b0};
                        wen_a13 = {1'b0, 1'b0};
                        wen_a12 = {1'b0, 1'b0};
                        wen_a11 = {1'b0, 1'b0};
                        wen_a10 = {1'b0, 1'b0};
                        wen_a9 = {1'b0, 1'b0};
                        wen_a8 = {1'b0, 1'b0};
                        wen_a7 = {1'b0, 1'b0};
                        wen_a6 = {1'b0, 1'b0};
                        wen_a5 = {1'b0, 1'b0};
                        wen_a4 = {1'b0, 1'b0};
                        wen_a3 = {1'b0, 1'b0};
                        wen_a2 = {wen, wen};
                        wen_a1 = {wen, wen};
                    end
                    default : begin
                        wen_a34 = {1'b0, 1'b0};
                        wen_a33 = {1'b0, 1'b0};
                        wen_a32 = {1'b0, 1'b0};
                        wen_a31 = {1'b0, 1'b0};
                        wen_a30 = {1'b0, 1'b0};
                        wen_a29 = {1'b0, 1'b0};
                        wen_a28 = {1'b0, 1'b0};
                        wen_a27 = {1'b0, 1'b0};
                        wen_a26 = {1'b0, 1'b0};
                        wen_a25 = {1'b0, 1'b0};
                        wen_a24 = {1'b0, 1'b0};
                        wen_a23 = {1'b0, 1'b0};
                        wen_a22 = {1'b0, 1'b0};
                        wen_a21 = {1'b0, 1'b0};
                        wen_a20 = {1'b0, 1'b0};
                        wen_a19 = {1'b0, 1'b0};
                        wen_a18 = {1'b0, 1'b0};
                        wen_a17 = {1'b0, 1'b0};
                        wen_a16 = {1'b0, 1'b0};
                        wen_a15 = {1'b0, 1'b0};
                        wen_a14 = {1'b0, 1'b0};
                        wen_a13 = {1'b0, 1'b0};
                        wen_a12 = {1'b0, 1'b0};
                        wen_a11 = {1'b0, 1'b0};
                        wen_a10 = {1'b0, 1'b0};
                        wen_a9 = {1'b0, 1'b0};
                        wen_a8 = {1'b0, 1'b0};
                        wen_a7 = {1'b0, 1'b0};
                        wen_a6 = {1'b0, 1'b0};
                        wen_a5 = {1'b0, 1'b0};
                        wen_a4 = {1'b0, 1'b0};
                        wen_a3 = {1'b0, 1'b0};
                        wen_a2 = {1'b0, 1'b0};
                        wen_a1 = {1'b0, 1'b0};
                    end
                endcase

                case (ckRdAddr[14:9])
                    6'b000000, 6'b000001, 6'b000010, 6'b000011,
                    6'b000100, 6'b000101, 6'b000110, 6'b000111,
                    6'b001000, 6'b001001, 6'b001010, 6'b001011,
                    6'b001100, 6'b001101, 6'b001110, 6'b001111,
                    6'b010000, 6'b010001, 6'b010010, 6'b010011,
                    6'b010100, 6'b010101, 6'b010110, 6'b010111,
                    6'b011000, 6'b011001, 6'b011010, 6'b011011,
                    6'b011100, 6'b011101, 6'b011110, 6'b011111 : begin
                        readData = {
                                        readData34[0],
                                        readData33[0],
                                        readData32[0],
                                        readData31[0],
                                        readData30[0],
                                        readData29[0],
                                        readData28[0],
                                        readData27[0],
                                        readData26[0],
                                        readData25[0],
                                        readData24[0],
                                        readData23[0],
                                        readData22[0],
                                        readData21[0],
                                        readData20[0],
                                        readData19[0],
                                        readData18[0],
                                        readData17[0],
                                        readData16[0],
                                        readData15[0],
                                        readData14[0],
                                        readData13[0],
                                        readData12[0],
                                        readData11[0],
                                        readData10[0],
                                        readData9[0],
                                        readData8[0],
                                        readData7[0],
                                        readData6[0],
                                        readData5[0],
                                        readData4[0],
                                        readData3[0]
                        };
                    end
                    6'b100000, 6'b100001 : begin
                        readData = {readData2[16:9],readData2[7:0],readData1[16:9],readData1[7:0]};
                    end
                    default : begin
                        readData = 32'b0;
                    end
                endcase
            end
            17920: begin
                width34 = 3'b000;
                width33 = 3'b000;
                width32 = 3'b000;
                width31 = 3'b000;
                width30 = 3'b000;
                width29 = 3'b000;
                width28 = 3'b000;
                width27 = 3'b000;
                width26 = 3'b000;
                width25 = 3'b000;
                width24 = 3'b000;
                width23 = 3'b000;
                width22 = 3'b000;
                width21 = 3'b000;
                width20 = 3'b000;
                width19 = 3'b000;
                width18 = 3'b000;
                width17 = 3'b000;
                width16 = 3'b000;
                width15 = 3'b000;
                width14 = 3'b000;
                width13 = 3'b000;
                width12 = 3'b000;
                width11 = 3'b000;
                width10 = 3'b000;
                width9 = 3'b000;
                width8 = 3'b000;
                width7 = 3'b000;
                width6 = 3'b000;
                width5 = 3'b000;
                width4 = 3'b000;
                width3 = 3'b000;
                width2 = 3'b100;
                width1 = 3'b100;
                width0 = 3'b101;

                writeAddr34 = {writeAddr[13:0]};
                writeAddr33 = {writeAddr[13:0]};
                writeAddr32 = {writeAddr[13:0]};
                writeAddr31 = {writeAddr[13:0]};
                writeAddr30 = {writeAddr[13:0]};
                writeAddr29 = {writeAddr[13:0]};
                writeAddr28 = {writeAddr[13:0]};
                writeAddr27 = {writeAddr[13:0]};
                writeAddr26 = {writeAddr[13:0]};
                writeAddr25 = {writeAddr[13:0]};
                writeAddr24 = {writeAddr[13:0]};
                writeAddr23 = {writeAddr[13:0]};
                writeAddr22 = {writeAddr[13:0]};
                writeAddr21 = {writeAddr[13:0]};
                writeAddr20 = {writeAddr[13:0]};
                writeAddr19 = {writeAddr[13:0]};
                writeAddr18 = {writeAddr[13:0]};
                writeAddr17 = {writeAddr[13:0]};
                writeAddr16 = {writeAddr[13:0]};
                writeAddr15 = {writeAddr[13:0]};
                writeAddr14 = {writeAddr[13:0]};
                writeAddr13 = {writeAddr[13:0]};
                writeAddr12 = {writeAddr[13:0]};
                writeAddr11 = {writeAddr[13:0]};
                writeAddr10 = {writeAddr[13:0]};
                writeAddr9 = {writeAddr[13:0]};
                writeAddr8 = {writeAddr[13:0]};
                writeAddr7 = {writeAddr[13:0]};
                writeAddr6 = {writeAddr[13:0]};
                writeAddr5 = {writeAddr[13:0]};
                writeAddr4 = {writeAddr[13:0]};
                writeAddr3 = {writeAddr[13:0]};
                writeAddr2 = {writeAddr[9:0], 4'b0};
                writeAddr1 = {writeAddr[9:0], 4'b0};
                writeAddr0 = {writeAddr[8:0], 5'b0};

                readAddr34 = {writeAddr[13:0]};
                readAddr33 = {writeAddr[13:0]};
                readAddr32 = {writeAddr[13:0]};
                readAddr31 = {writeAddr[13:0]};
                readAddr30 = {writeAddr[13:0]};
                readAddr29 = {writeAddr[13:0]};
                readAddr28 = {writeAddr[13:0]};
                readAddr27 = {writeAddr[13:0]};
                readAddr26 = {writeAddr[13:0]};
                readAddr25 = {writeAddr[13:0]};
                readAddr24 = {writeAddr[13:0]};
                readAddr23 = {writeAddr[13:0]};
                readAddr22 = {writeAddr[13:0]};
                readAddr21 = {writeAddr[13:0]};
                readAddr20 = {writeAddr[13:0]};
                readAddr19 = {writeAddr[13:0]};
                readAddr18 = {writeAddr[13:0]};
                readAddr17 = {writeAddr[13:0]};
                readAddr16 = {writeAddr[13:0]};
                readAddr15 = {writeAddr[13:0]};
                readAddr14 = {writeAddr[13:0]};
                readAddr13 = {writeAddr[13:0]};
                readAddr12 = {writeAddr[13:0]};
                readAddr11 = {writeAddr[13:0]};
                readAddr10 = {writeAddr[13:0]};
                readAddr9 = {writeAddr[13:0]};
                readAddr8 = {writeAddr[13:0]};
                readAddr7 = {writeAddr[13:0]};
                readAddr6 = {writeAddr[13:0]};
                readAddr5 = {writeAddr[13:0]};
                readAddr4 = {writeAddr[13:0]};
                readAddr3 = {writeAddr[13:0]};
                readAddr2  = {readAddr[9:0],  4'b0};
                readAddr1  = {readAddr[9:0],  4'b0};
                readAddr0  = {readAddr[8:0],  5'b0};

                writeData34 = {17'b0, writeData[31]};
                writeData33 = {17'b0, writeData[30]};
                writeData32 = {17'b0, writeData[29]};
                writeData31 = {17'b0, writeData[28]};
                writeData30 = {17'b0, writeData[27]};
                writeData29 = {17'b0, writeData[26]};
                writeData28 = {17'b0, writeData[25]};
                writeData27 = {17'b0, writeData[24]};
                writeData26 = {17'b0, writeData[23]};
                writeData25 = {17'b0, writeData[22]};
                writeData24 = {17'b0, writeData[21]};
                writeData23 = {17'b0, writeData[20]};
                writeData22 = {17'b0, writeData[19]};
                writeData21 = {17'b0, writeData[18]};
                writeData20 = {17'b0, writeData[17]};
                writeData19 = {17'b0, writeData[16]};
                writeData18 = {17'b0, writeData[15]};
                writeData17 = {17'b0, writeData[14]};
                writeData16 = {17'b0, writeData[13]};
                writeData15 = {17'b0, writeData[12]};
                writeData14 = {17'b0, writeData[11]};
                writeData13 = {17'b0, writeData[10]};
                writeData12 = {17'b0, writeData[9]};
                writeData11 = {17'b0, writeData[8]};
                writeData10 = {17'b0, writeData[7]};
                writeData9 = {17'b0, writeData[6]};
                writeData8 = {17'b0, writeData[5]};
                writeData7 = {17'b0, writeData[4]};
                writeData6 = {17'b0, writeData[3]};
                writeData5 = {17'b0, writeData[2]};
                writeData4 = {17'b0, writeData[1]};
                writeData3 = {17'b0, writeData[0]};
                writeData2 = {1'b0, writeData[31:24], 1'b0, writeData[23:16]};
                writeData1 = {1'b0, writeData[15:8], 1'b0, writeData[7:0]};
                writeData0 = {1'b0, writeData[31:24], 1'b0, writeData[23:16], 1'b0, writeData[15:8], 1'b0, writeData[7:0]};

                case (writeAddr[14:9])
                    6'b000000, 6'b000001, 6'b000010, 6'b000011,
                    6'b000100, 6'b000101, 6'b000110, 6'b000111,
                    6'b001000, 6'b001001, 6'b001010, 6'b001011,
                    6'b001100, 6'b001101, 6'b001110, 6'b001111,
                    6'b010000, 6'b010001, 6'b010010, 6'b010011,
                    6'b010100, 6'b010101, 6'b010110, 6'b010111,
                    6'b011000, 6'b011001, 6'b011010, 6'b011011,
                    6'b011100, 6'b011101, 6'b011110, 6'b011111 : begin
                        wen_a34 = {1'b0, wen};
                        wen_a33 = {1'b0, wen};
                        wen_a32 = {1'b0, wen};
                        wen_a31 = {1'b0, wen};
                        wen_a30 = {1'b0, wen};
                        wen_a29 = {1'b0, wen};
                        wen_a28 = {1'b0, wen};
                        wen_a27 = {1'b0, wen};
                        wen_a26 = {1'b0, wen};
                        wen_a25 = {1'b0, wen};
                        wen_a24 = {1'b0, wen};
                        wen_a23 = {1'b0, wen};
                        wen_a22 = {1'b0, wen};
                        wen_a21 = {1'b0, wen};
                        wen_a20 = {1'b0, wen};
                        wen_a19 = {1'b0, wen};
                        wen_a18 = {1'b0, wen};
                        wen_a17 = {1'b0, wen};
                        wen_a16 = {1'b0, wen};
                        wen_a15 = {1'b0, wen};
                        wen_a14 = {1'b0, wen};
                        wen_a13 = {1'b0, wen};
                        wen_a12 = {1'b0, wen};
                        wen_a11 = {1'b0, wen};
                        wen_a10 = {1'b0, wen};
                        wen_a9 = {1'b0, wen};
                        wen_a8 = {1'b0, wen};
                        wen_a7 = {1'b0, wen};
                        wen_a6 = {1'b0, wen};
                        wen_a5 = {1'b0, wen};
                        wen_a4 = {1'b0, wen};
                        wen_a3 = {1'b0, wen};
                        wen_a2 = {1'b0, 1'b0};
                        wen_a1 = {1'b0, 1'b0};
                        wen_a0 = {1'b0, 1'b0};
                        wen_b0 = {1'b0, 1'b0};
                    end
                    6'b100000, 6'b100001 : begin
                        wen_a34 = {1'b0, 1'b0};
                        wen_a33 = {1'b0, 1'b0};
                        wen_a32 = {1'b0, 1'b0};
                        wen_a31 = {1'b0, 1'b0};
                        wen_a30 = {1'b0, 1'b0};
                        wen_a29 = {1'b0, 1'b0};
                        wen_a28 = {1'b0, 1'b0};
                        wen_a27 = {1'b0, 1'b0};
                        wen_a26 = {1'b0, 1'b0};
                        wen_a25 = {1'b0, 1'b0};
                        wen_a24 = {1'b0, 1'b0};
                        wen_a23 = {1'b0, 1'b0};
                        wen_a22 = {1'b0, 1'b0};
                        wen_a21 = {1'b0, 1'b0};
                        wen_a20 = {1'b0, 1'b0};
                        wen_a19 = {1'b0, 1'b0};
                        wen_a18 = {1'b0, 1'b0};
                        wen_a17 = {1'b0, 1'b0};
                        wen_a16 = {1'b0, 1'b0};
                        wen_a15 = {1'b0, 1'b0};
                        wen_a14 = {1'b0, 1'b0};
                        wen_a13 = {1'b0, 1'b0};
                        wen_a12 = {1'b0, 1'b0};
                        wen_a11 = {1'b0, 1'b0};
                        wen_a10 = {1'b0, 1'b0};
                        wen_a9 = {1'b0, 1'b0};
                        wen_a8 = {1'b0, 1'b0};
                        wen_a7 = {1'b0, 1'b0};
                        wen_a6 = {1'b0, 1'b0};
                        wen_a5 = {1'b0, 1'b0};
                        wen_a4 = {1'b0, 1'b0};
                        wen_a3 = {1'b0, 1'b0};
                        wen_a2 = {wen, wen};
                        wen_a1 = {wen, wen};
                        wen_a0 = {1'b0, 1'b0};
                        wen_b0 = {1'b0, 1'b0};
                    end
                    6'b100010 : begin
                        wen_a34 = {1'b0, 1'b0};
                        wen_a33 = {1'b0, 1'b0};
                        wen_a32 = {1'b0, 1'b0};
                        wen_a31 = {1'b0, 1'b0};
                        wen_a30 = {1'b0, 1'b0};
                        wen_a29 = {1'b0, 1'b0};
                        wen_a28 = {1'b0, 1'b0};
                        wen_a27 = {1'b0, 1'b0};
                        wen_a26 = {1'b0, 1'b0};
                        wen_a25 = {1'b0, 1'b0};
                        wen_a24 = {1'b0, 1'b0};
                        wen_a23 = {1'b0, 1'b0};
                        wen_a22 = {1'b0, 1'b0};
                        wen_a21 = {1'b0, 1'b0};
                        wen_a20 = {1'b0, 1'b0};
                        wen_a19 = {1'b0, 1'b0};
                        wen_a18 = {1'b0, 1'b0};
                        wen_a17 = {1'b0, 1'b0};
                        wen_a16 = {1'b0, 1'b0};
                        wen_a15 = {1'b0, 1'b0};
                        wen_a14 = {1'b0, 1'b0};
                        wen_a13 = {1'b0, 1'b0};
                        wen_a12 = {1'b0, 1'b0};
                        wen_a11 = {1'b0, 1'b0};
                        wen_a10 = {1'b0, 1'b0};
                        wen_a9 = {1'b0, 1'b0};
                        wen_a8 = {1'b0, 1'b0};
                        wen_a7 = {1'b0, 1'b0};
                        wen_a6 = {1'b0, 1'b0};
                        wen_a5 = {1'b0, 1'b0};
                        wen_a4 = {1'b0, 1'b0};
                        wen_a3 = {1'b0, 1'b0};
                        wen_a2 = {1'b0, 1'b0};
                        wen_a1 = {1'b0, 1'b0};
                        wen_a0 = {wen, wen};
                        wen_b0 = {wen, wen};
                    end
                    default : begin
                        wen_a34 = {1'b0, 1'b0};
                        wen_a33 = {1'b0, 1'b0};
                        wen_a32 = {1'b0, 1'b0};
                        wen_a31 = {1'b0, 1'b0};
                        wen_a30 = {1'b0, 1'b0};
                        wen_a29 = {1'b0, 1'b0};
                        wen_a28 = {1'b0, 1'b0};
                        wen_a27 = {1'b0, 1'b0};
                        wen_a26 = {1'b0, 1'b0};
                        wen_a25 = {1'b0, 1'b0};
                        wen_a24 = {1'b0, 1'b0};
                        wen_a23 = {1'b0, 1'b0};
                        wen_a22 = {1'b0, 1'b0};
                        wen_a21 = {1'b0, 1'b0};
                        wen_a20 = {1'b0, 1'b0};
                        wen_a19 = {1'b0, 1'b0};
                        wen_a18 = {1'b0, 1'b0};
                        wen_a17 = {1'b0, 1'b0};
                        wen_a16 = {1'b0, 1'b0};
                        wen_a15 = {1'b0, 1'b0};
                        wen_a14 = {1'b0, 1'b0};
                        wen_a13 = {1'b0, 1'b0};
                        wen_a12 = {1'b0, 1'b0};
                        wen_a11 = {1'b0, 1'b0};
                        wen_a10 = {1'b0, 1'b0};
                        wen_a9 = {1'b0, 1'b0};
                        wen_a8 = {1'b0, 1'b0};
                        wen_a7 = {1'b0, 1'b0};
                        wen_a6 = {1'b0, 1'b0};
                        wen_a5 = {1'b0, 1'b0};
                        wen_a4 = {1'b0, 1'b0};
                        wen_a3 = {1'b0, 1'b0};
                        wen_a2 = {1'b0, 1'b0};
                        wen_a1 = {1'b0, 1'b0};
                        wen_a0 = {1'b0, 1'b0};
                        wen_b0 = {1'b0, 1'b0};
                    end
                endcase

                case (ckRdAddr[14:9])
                    6'b000000, 6'b000001, 6'b000010, 6'b000011,
                    6'b000100, 6'b000101, 6'b000110, 6'b000111,
                    6'b001000, 6'b001001, 6'b001010, 6'b001011,
                    6'b001100, 6'b001101, 6'b001110, 6'b001111,
                    6'b010000, 6'b010001, 6'b010010, 6'b010011,
                    6'b010100, 6'b010101, 6'b010110, 6'b010111,
                    6'b011000, 6'b011001, 6'b011010, 6'b011011,
                    6'b011100, 6'b011101, 6'b011110, 6'b011111 : begin
                        readData = {
                                        readData34[0],
                                        readData33[0],
                                        readData32[0],
                                        readData31[0],
                                        readData30[0],
                                        readData29[0],
                                        readData28[0],
                                        readData27[0],
                                        readData26[0],
                                        readData25[0],
                                        readData24[0],
                                        readData23[0],
                                        readData22[0],
                                        readData21[0],
                                        readData20[0],
                                        readData19[0],
                                        readData18[0],
                                        readData17[0],
                                        readData16[0],
                                        readData15[0],
                                        readData14[0],
                                        readData13[0],
                                        readData12[0],
                                        readData11[0],
                                        readData10[0],
                                        readData9[0],
                                        readData8[0],
                                        readData7[0],
                                        readData6[0],
                                        readData5[0],
                                        readData4[0],
                                        readData3[0]
                        };
                    end
                    6'b100000, 6'b100001 : begin
                        readData = {readData2[16:9],readData2[7:0],readData1[16:9],readData1[7:0]};
                    end
                    6'b100010 : begin
                        readData = {readData0[34:27],readData0[25:18],readData0[16:9],readData0[7:0]};
                    end
                    default : begin
                        readData = 32'b0;
                    end
                endcase
            end
            18432: begin
                width36 = 3'b000;
                width35 = 3'b000;
                width34 = 3'b000;
                width33 = 3'b000;
                width32 = 3'b000;
                width31 = 3'b000;
                width30 = 3'b000;
                width29 = 3'b000;
                width28 = 3'b000;
                width27 = 3'b000;
                width26 = 3'b000;
                width25 = 3'b000;
                width24 = 3'b000;
                width23 = 3'b000;
                width22 = 3'b000;
                width21 = 3'b000;
                width20 = 3'b000;
                width19 = 3'b000;
                width18 = 3'b000;
                width17 = 3'b000;
                width16 = 3'b000;
                width15 = 3'b000;
                width14 = 3'b000;
                width13 = 3'b000;
                width12 = 3'b000;
                width11 = 3'b000;
                width10 = 3'b000;
                width9 = 3'b000;
                width8 = 3'b000;
                width7 = 3'b000;
                width6 = 3'b000;
                width5 = 3'b000;
                width4 = 3'b011;
                width3 = 3'b011;
                width2 = 3'b011;
                width1 = 3'b011;

                writeAddr36 = {writeAddr[13:0]};
                writeAddr35 = {writeAddr[13:0]};
                writeAddr34 = {writeAddr[13:0]};
                writeAddr33 = {writeAddr[13:0]};
                writeAddr32 = {writeAddr[13:0]};
                writeAddr31 = {writeAddr[13:0]};
                writeAddr30 = {writeAddr[13:0]};
                writeAddr29 = {writeAddr[13:0]};
                writeAddr28 = {writeAddr[13:0]};
                writeAddr27 = {writeAddr[13:0]};
                writeAddr26 = {writeAddr[13:0]};
                writeAddr25 = {writeAddr[13:0]};
                writeAddr24 = {writeAddr[13:0]};
                writeAddr23 = {writeAddr[13:0]};
                writeAddr22 = {writeAddr[13:0]};
                writeAddr21 = {writeAddr[13:0]};
                writeAddr20 = {writeAddr[13:0]};
                writeAddr19 = {writeAddr[13:0]};
                writeAddr18 = {writeAddr[13:0]};
                writeAddr17 = {writeAddr[13:0]};
                writeAddr16 = {writeAddr[13:0]};
                writeAddr15 = {writeAddr[13:0]};
                writeAddr14 = {writeAddr[13:0]};
                writeAddr13 = {writeAddr[13:0]};
                writeAddr12 = {writeAddr[13:0]};
                writeAddr11 = {writeAddr[13:0]};
                writeAddr10 = {writeAddr[13:0]};
                writeAddr9 = {writeAddr[13:0]};
                writeAddr8 = {writeAddr[13:0]};
                writeAddr7 = {writeAddr[13:0]};
                writeAddr6 = {writeAddr[13:0]};
                writeAddr5 = {writeAddr[13:0]};
                writeAddr4 = {writeAddr[10:0], 3'b0};
                writeAddr3 = {writeAddr[10:0], 3'b0};
                writeAddr2 = {writeAddr[10:0], 3'b0};
                writeAddr1 = {writeAddr[10:0], 3'b0};

                readAddr36 = {writeAddr[13:0]};
                readAddr35 = {writeAddr[13:0]};
                readAddr34 = {writeAddr[13:0]};
                readAddr33 = {writeAddr[13:0]};
                readAddr32 = {writeAddr[13:0]};
                readAddr31 = {writeAddr[13:0]};
                readAddr30 = {writeAddr[13:0]};
                readAddr29 = {writeAddr[13:0]};
                readAddr28 = {writeAddr[13:0]};
                readAddr27 = {writeAddr[13:0]};
                readAddr26 = {writeAddr[13:0]};
                readAddr25 = {writeAddr[13:0]};
                readAddr24 = {writeAddr[13:0]};
                readAddr23 = {writeAddr[13:0]};
                readAddr22 = {writeAddr[13:0]};
                readAddr21 = {writeAddr[13:0]};
                readAddr20 = {writeAddr[13:0]};
                readAddr19 = {writeAddr[13:0]};
                readAddr18 = {writeAddr[13:0]};
                readAddr17 = {writeAddr[13:0]};
                readAddr16 = {writeAddr[13:0]};
                readAddr15 = {writeAddr[13:0]};
                readAddr14 = {writeAddr[13:0]};
                readAddr13 = {writeAddr[13:0]};
                readAddr12 = {writeAddr[13:0]};
                readAddr11 = {writeAddr[13:0]};
                readAddr10 = {writeAddr[13:0]};
                readAddr9 = {writeAddr[13:0]};
                readAddr8 = {writeAddr[13:0]};
                readAddr7 = {writeAddr[13:0]};
                readAddr6 = {writeAddr[13:0]};
                readAddr5 = {writeAddr[13:0]};
                readAddr4  = {readAddr[10:0],  3'b0};
                readAddr3  = {readAddr[10:0],  3'b0};
                readAddr2  = {readAddr[10:0],  3'b0};
                readAddr1  = {readAddr[10:0],  3'b0};

                writeData36 = {17'b0, writeData[31]};
                writeData35 = {17'b0, writeData[30]};
                writeData34 = {17'b0, writeData[29]};
                writeData33 = {17'b0, writeData[28]};
                writeData32 = {17'b0, writeData[27]};
                writeData31 = {17'b0, writeData[26]};
                writeData30 = {17'b0, writeData[25]};
                writeData29 = {17'b0, writeData[24]};
                writeData28 = {17'b0, writeData[23]};
                writeData27 = {17'b0, writeData[22]};
                writeData26 = {17'b0, writeData[21]};
                writeData25 = {17'b0, writeData[20]};
                writeData24 = {17'b0, writeData[19]};
                writeData23 = {17'b0, writeData[18]};
                writeData22 = {17'b0, writeData[17]};
                writeData21 = {17'b0, writeData[16]};
                writeData20 = {17'b0, writeData[15]};
                writeData19 = {17'b0, writeData[14]};
                writeData18 = {17'b0, writeData[13]};
                writeData17 = {17'b0, writeData[12]};
                writeData16 = {17'b0, writeData[11]};
                writeData15 = {17'b0, writeData[10]};
                writeData14 = {17'b0, writeData[9]};
                writeData13 = {17'b0, writeData[8]};
                writeData12 = {17'b0, writeData[7]};
                writeData11 = {17'b0, writeData[6]};
                writeData10 = {17'b0, writeData[5]};
                writeData9 = {17'b0, writeData[4]};
                writeData8 = {17'b0, writeData[3]};
                writeData7 = {17'b0, writeData[2]};
                writeData6 = {17'b0, writeData[1]};
                writeData5 = {17'b0, writeData[0]};
                writeData4 = {10'b0, writeData[31:24]};
                writeData3 = {10'b0, writeData[23:16]};
                writeData2 = {10'b0, writeData[15:8]};
                writeData1 = {10'b0, writeData[7:0]};

                case (writeAddr[14:9])
                    6'b000000, 6'b000001, 6'b000010, 6'b000011,
                    6'b000100, 6'b000101, 6'b000110, 6'b000111,
                    6'b001000, 6'b001001, 6'b001010, 6'b001011,
                    6'b001100, 6'b001101, 6'b001110, 6'b001111,
                    6'b010000, 6'b010001, 6'b010010, 6'b010011,
                    6'b010100, 6'b010101, 6'b010110, 6'b010111,
                    6'b011000, 6'b011001, 6'b011010, 6'b011011,
                    6'b011100, 6'b011101, 6'b011110, 6'b011111 : begin
                        wen_a36 = {1'b0, wen};
                        wen_a35 = {1'b0, wen};
                        wen_a34 = {1'b0, wen};
                        wen_a33 = {1'b0, wen};
                        wen_a32 = {1'b0, wen};
                        wen_a31 = {1'b0, wen};
                        wen_a30 = {1'b0, wen};
                        wen_a29 = {1'b0, wen};
                        wen_a28 = {1'b0, wen};
                        wen_a27 = {1'b0, wen};
                        wen_a26 = {1'b0, wen};
                        wen_a25 = {1'b0, wen};
                        wen_a24 = {1'b0, wen};
                        wen_a23 = {1'b0, wen};
                        wen_a22 = {1'b0, wen};
                        wen_a21 = {1'b0, wen};
                        wen_a20 = {1'b0, wen};
                        wen_a19 = {1'b0, wen};
                        wen_a18 = {1'b0, wen};
                        wen_a17 = {1'b0, wen};
                        wen_a16 = {1'b0, wen};
                        wen_a15 = {1'b0, wen};
                        wen_a14 = {1'b0, wen};
                        wen_a13 = {1'b0, wen};
                        wen_a12 = {1'b0, wen};
                        wen_a11 = {1'b0, wen};
                        wen_a10 = {1'b0, wen};
                        wen_a9 = {1'b0, wen};
                        wen_a8 = {1'b0, wen};
                        wen_a7 = {1'b0, wen};
                        wen_a6 = {1'b0, wen};
                        wen_a5 = {1'b0, wen};
                        wen_a4 = {1'b0, 1'b0};
                        wen_a3 = {1'b0, 1'b0};
                        wen_a2 = {1'b0, 1'b0};
                        wen_a1 = {1'b0, 1'b0};
                    end
                    6'b100000, 6'b100001, 6'b100010, 6'b100011 : begin
                        wen_a36 = {1'b0, 1'b0};
                        wen_a35 = {1'b0, 1'b0};
                        wen_a34 = {1'b0, 1'b0};
                        wen_a33 = {1'b0, 1'b0};
                        wen_a32 = {1'b0, 1'b0};
                        wen_a31 = {1'b0, 1'b0};
                        wen_a30 = {1'b0, 1'b0};
                        wen_a29 = {1'b0, 1'b0};
                        wen_a28 = {1'b0, 1'b0};
                        wen_a27 = {1'b0, 1'b0};
                        wen_a26 = {1'b0, 1'b0};
                        wen_a25 = {1'b0, 1'b0};
                        wen_a24 = {1'b0, 1'b0};
                        wen_a23 = {1'b0, 1'b0};
                        wen_a22 = {1'b0, 1'b0};
                        wen_a21 = {1'b0, 1'b0};
                        wen_a20 = {1'b0, 1'b0};
                        wen_a19 = {1'b0, 1'b0};
                        wen_a18 = {1'b0, 1'b0};
                        wen_a17 = {1'b0, 1'b0};
                        wen_a16 = {1'b0, 1'b0};
                        wen_a15 = {1'b0, 1'b0};
                        wen_a14 = {1'b0, 1'b0};
                        wen_a13 = {1'b0, 1'b0};
                        wen_a12 = {1'b0, 1'b0};
                        wen_a11 = {1'b0, 1'b0};
                        wen_a10 = {1'b0, 1'b0};
                        wen_a9 = {1'b0, 1'b0};
                        wen_a8 = {1'b0, 1'b0};
                        wen_a7 = {1'b0, 1'b0};
                        wen_a6 = {1'b0, 1'b0};
                        wen_a5 = {1'b0, 1'b0};
                        wen_a4 = {1'b0, wen};
                        wen_a3 = {1'b0, wen};
                        wen_a2 = {1'b0, wen};
                        wen_a1 = {1'b0, wen};
                    end
                    default : begin
                        wen_a36 = {1'b0, 1'b0};
                        wen_a35 = {1'b0, 1'b0};
                        wen_a34 = {1'b0, 1'b0};
                        wen_a33 = {1'b0, 1'b0};
                        wen_a32 = {1'b0, 1'b0};
                        wen_a31 = {1'b0, 1'b0};
                        wen_a30 = {1'b0, 1'b0};
                        wen_a29 = {1'b0, 1'b0};
                        wen_a28 = {1'b0, 1'b0};
                        wen_a27 = {1'b0, 1'b0};
                        wen_a26 = {1'b0, 1'b0};
                        wen_a25 = {1'b0, 1'b0};
                        wen_a24 = {1'b0, 1'b0};
                        wen_a23 = {1'b0, 1'b0};
                        wen_a22 = {1'b0, 1'b0};
                        wen_a21 = {1'b0, 1'b0};
                        wen_a20 = {1'b0, 1'b0};
                        wen_a19 = {1'b0, 1'b0};
                        wen_a18 = {1'b0, 1'b0};
                        wen_a17 = {1'b0, 1'b0};
                        wen_a16 = {1'b0, 1'b0};
                        wen_a15 = {1'b0, 1'b0};
                        wen_a14 = {1'b0, 1'b0};
                        wen_a13 = {1'b0, 1'b0};
                        wen_a12 = {1'b0, 1'b0};
                        wen_a11 = {1'b0, 1'b0};
                        wen_a10 = {1'b0, 1'b0};
                        wen_a9 = {1'b0, 1'b0};
                        wen_a8 = {1'b0, 1'b0};
                        wen_a7 = {1'b0, 1'b0};
                        wen_a6 = {1'b0, 1'b0};
                        wen_a5 = {1'b0, 1'b0};
                        wen_a4 = {1'b0, 1'b0};
                        wen_a3 = {1'b0, 1'b0};
                        wen_a2 = {1'b0, 1'b0};
                        wen_a1 = {1'b0, 1'b0};
                    end
                endcase

                case (ckRdAddr[14:9])
                    6'b000000, 6'b000001, 6'b000010, 6'b000011,
                    6'b000100, 6'b000101, 6'b000110, 6'b000111,
                    6'b001000, 6'b001001, 6'b001010, 6'b001011,
                    6'b001100, 6'b001101, 6'b001110, 6'b001111,
                    6'b010000, 6'b010001, 6'b010010, 6'b010011,
                    6'b010100, 6'b010101, 6'b010110, 6'b010111,
                    6'b011000, 6'b011001, 6'b011010, 6'b011011,
                    6'b011100, 6'b011101, 6'b011110, 6'b011111 : begin
                        readData = {
                                        readData36[0],
                                        readData35[0],
                                        readData34[0],
                                        readData33[0],
                                        readData32[0],
                                        readData31[0],
                                        readData30[0],
                                        readData29[0],
                                        readData28[0],
                                        readData27[0],
                                        readData26[0],
                                        readData25[0],
                                        readData24[0],
                                        readData23[0],
                                        readData22[0],
                                        readData21[0],
                                        readData20[0],
                                        readData19[0],
                                        readData18[0],
                                        readData17[0],
                                        readData16[0],
                                        readData15[0],
                                        readData14[0],
                                        readData13[0],
                                        readData12[0],
                                        readData11[0],
                                        readData10[0],
                                        readData9[0],
                                        readData8[0],
                                        readData7[0],
                                        readData6[0],
                                        readData5[0]
                        };
                    end
                    6'b100000, 6'b100001, 6'b100010, 6'b100011 : begin
                        readData = {readData4[7:0],readData3[7:0],readData2[7:0],readData1[7:0]};
                    end
                    default : begin
                        readData = 32'b0;
                    end
                endcase
            end
            18944: begin
                width36 = 3'b000;
                width35 = 3'b000;
                width34 = 3'b000;
                width33 = 3'b000;
                width32 = 3'b000;
                width31 = 3'b000;
                width30 = 3'b000;
                width29 = 3'b000;
                width28 = 3'b000;
                width27 = 3'b000;
                width26 = 3'b000;
                width25 = 3'b000;
                width24 = 3'b000;
                width23 = 3'b000;
                width22 = 3'b000;
                width21 = 3'b000;
                width20 = 3'b000;
                width19 = 3'b000;
                width18 = 3'b000;
                width17 = 3'b000;
                width16 = 3'b000;
                width15 = 3'b000;
                width14 = 3'b000;
                width13 = 3'b000;
                width12 = 3'b000;
                width11 = 3'b000;
                width10 = 3'b000;
                width9 = 3'b000;
                width8 = 3'b000;
                width7 = 3'b000;
                width6 = 3'b000;
                width5 = 3'b000;
                width4 = 3'b011;
                width3 = 3'b011;
                width2 = 3'b011;
                width1 = 3'b011;
                width0 = 3'b101;

                writeAddr36 = {writeAddr[13:0]};
                writeAddr35 = {writeAddr[13:0]};
                writeAddr34 = {writeAddr[13:0]};
                writeAddr33 = {writeAddr[13:0]};
                writeAddr32 = {writeAddr[13:0]};
                writeAddr31 = {writeAddr[13:0]};
                writeAddr30 = {writeAddr[13:0]};
                writeAddr29 = {writeAddr[13:0]};
                writeAddr28 = {writeAddr[13:0]};
                writeAddr27 = {writeAddr[13:0]};
                writeAddr26 = {writeAddr[13:0]};
                writeAddr25 = {writeAddr[13:0]};
                writeAddr24 = {writeAddr[13:0]};
                writeAddr23 = {writeAddr[13:0]};
                writeAddr22 = {writeAddr[13:0]};
                writeAddr21 = {writeAddr[13:0]};
                writeAddr20 = {writeAddr[13:0]};
                writeAddr19 = {writeAddr[13:0]};
                writeAddr18 = {writeAddr[13:0]};
                writeAddr17 = {writeAddr[13:0]};
                writeAddr16 = {writeAddr[13:0]};
                writeAddr15 = {writeAddr[13:0]};
                writeAddr14 = {writeAddr[13:0]};
                writeAddr13 = {writeAddr[13:0]};
                writeAddr12 = {writeAddr[13:0]};
                writeAddr11 = {writeAddr[13:0]};
                writeAddr10 = {writeAddr[13:0]};
                writeAddr9 = {writeAddr[13:0]};
                writeAddr8 = {writeAddr[13:0]};
                writeAddr7 = {writeAddr[13:0]};
                writeAddr6 = {writeAddr[13:0]};
                writeAddr5 = {writeAddr[13:0]};
                writeAddr4 = {writeAddr[10:0], 3'b0};
                writeAddr3 = {writeAddr[10:0], 3'b0};
                writeAddr2 = {writeAddr[10:0], 3'b0};
                writeAddr1 = {writeAddr[10:0], 3'b0};
                writeAddr0 = {writeAddr[8:0], 5'b0};

                readAddr36 = {writeAddr[13:0]};
                readAddr35 = {writeAddr[13:0]};
                readAddr34 = {writeAddr[13:0]};
                readAddr33 = {writeAddr[13:0]};
                readAddr32 = {writeAddr[13:0]};
                readAddr31 = {writeAddr[13:0]};
                readAddr30 = {writeAddr[13:0]};
                readAddr29 = {writeAddr[13:0]};
                readAddr28 = {writeAddr[13:0]};
                readAddr27 = {writeAddr[13:0]};
                readAddr26 = {writeAddr[13:0]};
                readAddr25 = {writeAddr[13:0]};
                readAddr24 = {writeAddr[13:0]};
                readAddr23 = {writeAddr[13:0]};
                readAddr22 = {writeAddr[13:0]};
                readAddr21 = {writeAddr[13:0]};
                readAddr20 = {writeAddr[13:0]};
                readAddr19 = {writeAddr[13:0]};
                readAddr18 = {writeAddr[13:0]};
                readAddr17 = {writeAddr[13:0]};
                readAddr16 = {writeAddr[13:0]};
                readAddr15 = {writeAddr[13:0]};
                readAddr14 = {writeAddr[13:0]};
                readAddr13 = {writeAddr[13:0]};
                readAddr12 = {writeAddr[13:0]};
                readAddr11 = {writeAddr[13:0]};
                readAddr10 = {writeAddr[13:0]};
                readAddr9 = {writeAddr[13:0]};
                readAddr8 = {writeAddr[13:0]};
                readAddr7 = {writeAddr[13:0]};
                readAddr6 = {writeAddr[13:0]};
                readAddr5 = {writeAddr[13:0]};
                readAddr4  = {readAddr[10:0],  3'b0};
                readAddr3  = {readAddr[10:0],  3'b0};
                readAddr2  = {readAddr[10:0],  3'b0};
                readAddr1  = {readAddr[10:0],  3'b0};
                readAddr0  = {readAddr[8:0],  5'b0};

                writeData36 = {17'b0, writeData[31]};
                writeData35 = {17'b0, writeData[30]};
                writeData34 = {17'b0, writeData[29]};
                writeData33 = {17'b0, writeData[28]};
                writeData32 = {17'b0, writeData[27]};
                writeData31 = {17'b0, writeData[26]};
                writeData30 = {17'b0, writeData[25]};
                writeData29 = {17'b0, writeData[24]};
                writeData28 = {17'b0, writeData[23]};
                writeData27 = {17'b0, writeData[22]};
                writeData26 = {17'b0, writeData[21]};
                writeData25 = {17'b0, writeData[20]};
                writeData24 = {17'b0, writeData[19]};
                writeData23 = {17'b0, writeData[18]};
                writeData22 = {17'b0, writeData[17]};
                writeData21 = {17'b0, writeData[16]};
                writeData20 = {17'b0, writeData[15]};
                writeData19 = {17'b0, writeData[14]};
                writeData18 = {17'b0, writeData[13]};
                writeData17 = {17'b0, writeData[12]};
                writeData16 = {17'b0, writeData[11]};
                writeData15 = {17'b0, writeData[10]};
                writeData14 = {17'b0, writeData[9]};
                writeData13 = {17'b0, writeData[8]};
                writeData12 = {17'b0, writeData[7]};
                writeData11 = {17'b0, writeData[6]};
                writeData10 = {17'b0, writeData[5]};
                writeData9 = {17'b0, writeData[4]};
                writeData8 = {17'b0, writeData[3]};
                writeData7 = {17'b0, writeData[2]};
                writeData6 = {17'b0, writeData[1]};
                writeData5 = {17'b0, writeData[0]};
                writeData4 = {10'b0, writeData[31:24]};
                writeData3 = {10'b0, writeData[23:16]};
                writeData2 = {10'b0, writeData[15:8]};
                writeData1 = {10'b0, writeData[7:0]};
                writeData0 = {1'b0, writeData[31:24], 1'b0, writeData[23:16], 1'b0, writeData[15:8], 1'b0, writeData[7:0]};

                case (writeAddr[14:9])
                    6'b000000, 6'b000001, 6'b000010, 6'b000011,
                    6'b000100, 6'b000101, 6'b000110, 6'b000111,
                    6'b001000, 6'b001001, 6'b001010, 6'b001011,
                    6'b001100, 6'b001101, 6'b001110, 6'b001111,
                    6'b010000, 6'b010001, 6'b010010, 6'b010011,
                    6'b010100, 6'b010101, 6'b010110, 6'b010111,
                    6'b011000, 6'b011001, 6'b011010, 6'b011011,
                    6'b011100, 6'b011101, 6'b011110, 6'b011111 : begin
                        wen_a36 = {1'b0, wen};
                        wen_a35 = {1'b0, wen};
                        wen_a34 = {1'b0, wen};
                        wen_a33 = {1'b0, wen};
                        wen_a32 = {1'b0, wen};
                        wen_a31 = {1'b0, wen};
                        wen_a30 = {1'b0, wen};
                        wen_a29 = {1'b0, wen};
                        wen_a28 = {1'b0, wen};
                        wen_a27 = {1'b0, wen};
                        wen_a26 = {1'b0, wen};
                        wen_a25 = {1'b0, wen};
                        wen_a24 = {1'b0, wen};
                        wen_a23 = {1'b0, wen};
                        wen_a22 = {1'b0, wen};
                        wen_a21 = {1'b0, wen};
                        wen_a20 = {1'b0, wen};
                        wen_a19 = {1'b0, wen};
                        wen_a18 = {1'b0, wen};
                        wen_a17 = {1'b0, wen};
                        wen_a16 = {1'b0, wen};
                        wen_a15 = {1'b0, wen};
                        wen_a14 = {1'b0, wen};
                        wen_a13 = {1'b0, wen};
                        wen_a12 = {1'b0, wen};
                        wen_a11 = {1'b0, wen};
                        wen_a10 = {1'b0, wen};
                        wen_a9 = {1'b0, wen};
                        wen_a8 = {1'b0, wen};
                        wen_a7 = {1'b0, wen};
                        wen_a6 = {1'b0, wen};
                        wen_a5 = {1'b0, wen};
                        wen_a4 = {1'b0, 1'b0};
                        wen_a3 = {1'b0, 1'b0};
                        wen_a2 = {1'b0, 1'b0};
                        wen_a1 = {1'b0, 1'b0};
                        wen_a0 = {1'b0, 1'b0};
                        wen_b0 = {1'b0, 1'b0};
                    end
                    6'b100000, 6'b100001, 6'b100010, 6'b100011 : begin
                        wen_a36 = {1'b0, 1'b0};
                        wen_a35 = {1'b0, 1'b0};
                        wen_a34 = {1'b0, 1'b0};
                        wen_a33 = {1'b0, 1'b0};
                        wen_a32 = {1'b0, 1'b0};
                        wen_a31 = {1'b0, 1'b0};
                        wen_a30 = {1'b0, 1'b0};
                        wen_a29 = {1'b0, 1'b0};
                        wen_a28 = {1'b0, 1'b0};
                        wen_a27 = {1'b0, 1'b0};
                        wen_a26 = {1'b0, 1'b0};
                        wen_a25 = {1'b0, 1'b0};
                        wen_a24 = {1'b0, 1'b0};
                        wen_a23 = {1'b0, 1'b0};
                        wen_a22 = {1'b0, 1'b0};
                        wen_a21 = {1'b0, 1'b0};
                        wen_a20 = {1'b0, 1'b0};
                        wen_a19 = {1'b0, 1'b0};
                        wen_a18 = {1'b0, 1'b0};
                        wen_a17 = {1'b0, 1'b0};
                        wen_a16 = {1'b0, 1'b0};
                        wen_a15 = {1'b0, 1'b0};
                        wen_a14 = {1'b0, 1'b0};
                        wen_a13 = {1'b0, 1'b0};
                        wen_a12 = {1'b0, 1'b0};
                        wen_a11 = {1'b0, 1'b0};
                        wen_a10 = {1'b0, 1'b0};
                        wen_a9 = {1'b0, 1'b0};
                        wen_a8 = {1'b0, 1'b0};
                        wen_a7 = {1'b0, 1'b0};
                        wen_a6 = {1'b0, 1'b0};
                        wen_a5 = {1'b0, 1'b0};
                        wen_a4 = {1'b0, wen};
                        wen_a3 = {1'b0, wen};
                        wen_a2 = {1'b0, wen};
                        wen_a1 = {1'b0, wen};
                        wen_a0 = {1'b0, 1'b0};
                        wen_b0 = {1'b0, 1'b0};
                    end
                    6'b100100 : begin
                        wen_a36 = {1'b0, 1'b0};
                        wen_a35 = {1'b0, 1'b0};
                        wen_a34 = {1'b0, 1'b0};
                        wen_a33 = {1'b0, 1'b0};
                        wen_a32 = {1'b0, 1'b0};
                        wen_a31 = {1'b0, 1'b0};
                        wen_a30 = {1'b0, 1'b0};
                        wen_a29 = {1'b0, 1'b0};
                        wen_a28 = {1'b0, 1'b0};
                        wen_a27 = {1'b0, 1'b0};
                        wen_a26 = {1'b0, 1'b0};
                        wen_a25 = {1'b0, 1'b0};
                        wen_a24 = {1'b0, 1'b0};
                        wen_a23 = {1'b0, 1'b0};
                        wen_a22 = {1'b0, 1'b0};
                        wen_a21 = {1'b0, 1'b0};
                        wen_a20 = {1'b0, 1'b0};
                        wen_a19 = {1'b0, 1'b0};
                        wen_a18 = {1'b0, 1'b0};
                        wen_a17 = {1'b0, 1'b0};
                        wen_a16 = {1'b0, 1'b0};
                        wen_a15 = {1'b0, 1'b0};
                        wen_a14 = {1'b0, 1'b0};
                        wen_a13 = {1'b0, 1'b0};
                        wen_a12 = {1'b0, 1'b0};
                        wen_a11 = {1'b0, 1'b0};
                        wen_a10 = {1'b0, 1'b0};
                        wen_a9 = {1'b0, 1'b0};
                        wen_a8 = {1'b0, 1'b0};
                        wen_a7 = {1'b0, 1'b0};
                        wen_a6 = {1'b0, 1'b0};
                        wen_a5 = {1'b0, 1'b0};
                        wen_a4 = {1'b0, 1'b0};
                        wen_a3 = {1'b0, 1'b0};
                        wen_a2 = {1'b0, 1'b0};
                        wen_a1 = {1'b0, 1'b0};
                        wen_a0 = {wen,  wen};
                        wen_b0 = {wen,  wen};
                    end
                    default : begin
                        wen_a36 = {1'b0, 1'b0};
                        wen_a35 = {1'b0, 1'b0};
                        wen_a34 = {1'b0, 1'b0};
                        wen_a33 = {1'b0, 1'b0};
                        wen_a32 = {1'b0, 1'b0};
                        wen_a31 = {1'b0, 1'b0};
                        wen_a30 = {1'b0, 1'b0};
                        wen_a29 = {1'b0, 1'b0};
                        wen_a28 = {1'b0, 1'b0};
                        wen_a27 = {1'b0, 1'b0};
                        wen_a26 = {1'b0, 1'b0};
                        wen_a25 = {1'b0, 1'b0};
                        wen_a24 = {1'b0, 1'b0};
                        wen_a23 = {1'b0, 1'b0};
                        wen_a22 = {1'b0, 1'b0};
                        wen_a21 = {1'b0, 1'b0};
                        wen_a20 = {1'b0, 1'b0};
                        wen_a19 = {1'b0, 1'b0};
                        wen_a18 = {1'b0, 1'b0};
                        wen_a17 = {1'b0, 1'b0};
                        wen_a16 = {1'b0, 1'b0};
                        wen_a15 = {1'b0, 1'b0};
                        wen_a14 = {1'b0, 1'b0};
                        wen_a13 = {1'b0, 1'b0};
                        wen_a12 = {1'b0, 1'b0};
                        wen_a11 = {1'b0, 1'b0};
                        wen_a10 = {1'b0, 1'b0};
                        wen_a9 = {1'b0, 1'b0};
                        wen_a8 = {1'b0, 1'b0};
                        wen_a7 = {1'b0, 1'b0};
                        wen_a6 = {1'b0, 1'b0};
                        wen_a5 = {1'b0, 1'b0};
                        wen_a4 = {1'b0, 1'b0};
                        wen_a3 = {1'b0, 1'b0};
                        wen_a2 = {1'b0, 1'b0};
                        wen_a1 = {1'b0, 1'b0};
                        wen_a0 = {1'b0, 1'b0};
                        wen_b0 = {1'b0, 1'b0};
                    end
                endcase

                case (ckRdAddr[14:9])
                    6'b000000, 6'b000001, 6'b000010, 6'b000011,
                    6'b000100, 6'b000101, 6'b000110, 6'b000111,
                    6'b001000, 6'b001001, 6'b001010, 6'b001011,
                    6'b001100, 6'b001101, 6'b001110, 6'b001111,
                    6'b010000, 6'b010001, 6'b010010, 6'b010011,
                    6'b010100, 6'b010101, 6'b010110, 6'b010111,
                    6'b011000, 6'b011001, 6'b011010, 6'b011011,
                    6'b011100, 6'b011101, 6'b011110, 6'b011111 : begin
                        readData = {
                                        readData36[0],
                                        readData35[0],
                                        readData34[0],
                                        readData33[0],
                                        readData32[0],
                                        readData31[0],
                                        readData30[0],
                                        readData29[0],
                                        readData28[0],
                                        readData27[0],
                                        readData26[0],
                                        readData25[0],
                                        readData24[0],
                                        readData23[0],
                                        readData22[0],
                                        readData21[0],
                                        readData20[0],
                                        readData19[0],
                                        readData18[0],
                                        readData17[0],
                                        readData16[0],
                                        readData15[0],
                                        readData14[0],
                                        readData13[0],
                                        readData12[0],
                                        readData11[0],
                                        readData10[0],
                                        readData9[0],
                                        readData8[0],
                                        readData7[0],
                                        readData6[0],
                                        readData5[0]
                        };
                    end
                    6'b100000, 6'b100001, 6'b100010, 6'b100011 : begin
                        readData = {readData4[7:0],readData3[7:0],readData2[7:0],readData1[7:0]};
                    end
                    6'b100100 : begin
                        readData = {readData0[34:27],readData0[25:18],readData0[16:9],readData0[7:0]};
                    end
                    default : begin
                        readData = 32'b0;
                    end
                endcase
            end
            19456: begin
                width38 = 3'b000;
                width37 = 3'b000;
                width36 = 3'b000;
                width35 = 3'b000;
                width34 = 3'b000;
                width33 = 3'b000;
                width32 = 3'b000;
                width31 = 3'b000;
                width30 = 3'b000;
                width29 = 3'b000;
                width28 = 3'b000;
                width27 = 3'b000;
                width26 = 3'b000;
                width25 = 3'b000;
                width24 = 3'b000;
                width23 = 3'b000;
                width22 = 3'b000;
                width21 = 3'b000;
                width20 = 3'b000;
                width19 = 3'b000;
                width18 = 3'b000;
                width17 = 3'b000;
                width16 = 3'b000;
                width15 = 3'b000;
                width14 = 3'b000;
                width13 = 3'b000;
                width12 = 3'b000;
                width11 = 3'b000;
                width10 = 3'b000;
                width9 = 3'b000;
                width8 = 3'b000;
                width7 = 3'b000;
                width6 = 3'b011;
                width5 = 3'b011;
                width4 = 3'b011;
                width3 = 3'b011;
                width2 = 3'b100;
                width1 = 3'b100;

                writeAddr38 = {writeAddr[13:0]};
                writeAddr37 = {writeAddr[13:0]};
                writeAddr36 = {writeAddr[13:0]};
                writeAddr35 = {writeAddr[13:0]};
                writeAddr34 = {writeAddr[13:0]};
                writeAddr33 = {writeAddr[13:0]};
                writeAddr32 = {writeAddr[13:0]};
                writeAddr31 = {writeAddr[13:0]};
                writeAddr30 = {writeAddr[13:0]};
                writeAddr29 = {writeAddr[13:0]};
                writeAddr28 = {writeAddr[13:0]};
                writeAddr27 = {writeAddr[13:0]};
                writeAddr26 = {writeAddr[13:0]};
                writeAddr25 = {writeAddr[13:0]};
                writeAddr24 = {writeAddr[13:0]};
                writeAddr23 = {writeAddr[13:0]};
                writeAddr22 = {writeAddr[13:0]};
                writeAddr21 = {writeAddr[13:0]};
                writeAddr20 = {writeAddr[13:0]};
                writeAddr19 = {writeAddr[13:0]};
                writeAddr18 = {writeAddr[13:0]};
                writeAddr17 = {writeAddr[13:0]};
                writeAddr16 = {writeAddr[13:0]};
                writeAddr15 = {writeAddr[13:0]};
                writeAddr14 = {writeAddr[13:0]};
                writeAddr13 = {writeAddr[13:0]};
                writeAddr12 = {writeAddr[13:0]};
                writeAddr11 = {writeAddr[13:0]};
                writeAddr10 = {writeAddr[13:0]};
                writeAddr9 = {writeAddr[13:0]};
                writeAddr8 = {writeAddr[13:0]};
                writeAddr7 = {writeAddr[13:0]};
                writeAddr6 = {writeAddr[10:0], 3'b0};
                writeAddr5 = {writeAddr[10:0], 3'b0};
                writeAddr4 = {writeAddr[10:0], 3'b0};
                writeAddr3 = {writeAddr[10:0], 3'b0};
                writeAddr2 = {writeAddr[9:0], 4'b0};
                writeAddr1 = {writeAddr[9:0], 4'b0};

                readAddr38 = {writeAddr[13:0]};
                readAddr37 = {writeAddr[13:0]};
                readAddr36 = {writeAddr[13:0]};
                readAddr35 = {writeAddr[13:0]};
                readAddr34 = {writeAddr[13:0]};
                readAddr33 = {writeAddr[13:0]};
                readAddr32 = {writeAddr[13:0]};
                readAddr31 = {writeAddr[13:0]};
                readAddr30 = {writeAddr[13:0]};
                readAddr29 = {writeAddr[13:0]};
                readAddr28 = {writeAddr[13:0]};
                readAddr27 = {writeAddr[13:0]};
                readAddr26 = {writeAddr[13:0]};
                readAddr25 = {writeAddr[13:0]};
                readAddr24 = {writeAddr[13:0]};
                readAddr23 = {writeAddr[13:0]};
                readAddr22 = {writeAddr[13:0]};
                readAddr21 = {writeAddr[13:0]};
                readAddr20 = {writeAddr[13:0]};
                readAddr19 = {writeAddr[13:0]};
                readAddr18 = {writeAddr[13:0]};
                readAddr17 = {writeAddr[13:0]};
                readAddr16 = {writeAddr[13:0]};
                readAddr15 = {writeAddr[13:0]};
                readAddr14 = {writeAddr[13:0]};
                readAddr13 = {writeAddr[13:0]};
                readAddr12 = {writeAddr[13:0]};
                readAddr11 = {writeAddr[13:0]};
                readAddr10 = {writeAddr[13:0]};
                readAddr9 = {writeAddr[13:0]};
                readAddr8 = {writeAddr[13:0]};
                readAddr7 = {writeAddr[13:0]};
                readAddr6  = {readAddr[10:0],  3'b0};
                readAddr5  = {readAddr[10:0],  3'b0};
                readAddr4  = {readAddr[10:0],  3'b0};
                readAddr3  = {readAddr[10:0],  3'b0};
                readAddr2  = {readAddr[9:0],  4'b0};
                readAddr1  = {readAddr[9:0],  4'b0};

                writeData38 = {17'b0, writeData[31]};
                writeData37 = {17'b0, writeData[30]};
                writeData36 = {17'b0, writeData[29]};
                writeData35 = {17'b0, writeData[28]};
                writeData34 = {17'b0, writeData[27]};
                writeData33 = {17'b0, writeData[26]};
                writeData32 = {17'b0, writeData[25]};
                writeData31 = {17'b0, writeData[24]};
                writeData30 = {17'b0, writeData[23]};
                writeData29 = {17'b0, writeData[22]};
                writeData28 = {17'b0, writeData[21]};
                writeData27 = {17'b0, writeData[20]};
                writeData26 = {17'b0, writeData[19]};
                writeData25 = {17'b0, writeData[18]};
                writeData24 = {17'b0, writeData[17]};
                writeData23 = {17'b0, writeData[16]};
                writeData22 = {17'b0, writeData[15]};
                writeData21 = {17'b0, writeData[14]};
                writeData20 = {17'b0, writeData[13]};
                writeData19 = {17'b0, writeData[12]};
                writeData18 = {17'b0, writeData[11]};
                writeData17 = {17'b0, writeData[10]};
                writeData16 = {17'b0, writeData[9]};
                writeData15 = {17'b0, writeData[8]};
                writeData14 = {17'b0, writeData[7]};
                writeData13 = {17'b0, writeData[6]};
                writeData12 = {17'b0, writeData[5]};
                writeData11 = {17'b0, writeData[4]};
                writeData10 = {17'b0, writeData[3]};
                writeData9 = {17'b0, writeData[2]};
                writeData8 = {17'b0, writeData[1]};
                writeData7 = {17'b0, writeData[0]};
                writeData6 = {10'b0, writeData[31:24]};
                writeData5 = {10'b0, writeData[23:16]};
                writeData4 = {10'b0, writeData[15:8]};
                writeData3 = {10'b0, writeData[7:0]};
                writeData2 = {1'b0, writeData[31:24], 1'b0, writeData[23:16]};
                writeData1 = {1'b0, writeData[15:8], 1'b0, writeData[7:0]};

                case (writeAddr[14:9])
                    6'b000000, 6'b000001, 6'b000010, 6'b000011,
                    6'b000100, 6'b000101, 6'b000110, 6'b000111,
                    6'b001000, 6'b001001, 6'b001010, 6'b001011,
                    6'b001100, 6'b001101, 6'b001110, 6'b001111,
                    6'b010000, 6'b010001, 6'b010010, 6'b010011,
                    6'b010100, 6'b010101, 6'b010110, 6'b010111,
                    6'b011000, 6'b011001, 6'b011010, 6'b011011,
                    6'b011100, 6'b011101, 6'b011110, 6'b011111 : begin
                        wen_a38 = {1'b0, wen};
                        wen_a37 = {1'b0, wen};
                        wen_a36 = {1'b0, wen};
                        wen_a35 = {1'b0, wen};
                        wen_a34 = {1'b0, wen};
                        wen_a33 = {1'b0, wen};
                        wen_a32 = {1'b0, wen};
                        wen_a31 = {1'b0, wen};
                        wen_a30 = {1'b0, wen};
                        wen_a29 = {1'b0, wen};
                        wen_a28 = {1'b0, wen};
                        wen_a27 = {1'b0, wen};
                        wen_a26 = {1'b0, wen};
                        wen_a25 = {1'b0, wen};
                        wen_a24 = {1'b0, wen};
                        wen_a23 = {1'b0, wen};
                        wen_a22 = {1'b0, wen};
                        wen_a21 = {1'b0, wen};
                        wen_a20 = {1'b0, wen};
                        wen_a19 = {1'b0, wen};
                        wen_a18 = {1'b0, wen};
                        wen_a17 = {1'b0, wen};
                        wen_a16 = {1'b0, wen};
                        wen_a15 = {1'b0, wen};
                        wen_a14 = {1'b0, wen};
                        wen_a13 = {1'b0, wen};
                        wen_a12 = {1'b0, wen};
                        wen_a11 = {1'b0, wen};
                        wen_a10 = {1'b0, wen};
                        wen_a9 = {1'b0, wen};
                        wen_a8 = {1'b0, wen};
                        wen_a7 = {1'b0, wen};
                        wen_a6 = {1'b0, 1'b0};
                        wen_a5 = {1'b0, 1'b0};
                        wen_a4 = {1'b0, 1'b0};
                        wen_a3 = {1'b0, 1'b0};
                        wen_a2 = {1'b0, 1'b0};
                        wen_a1 = {1'b0, 1'b0};
                    end
                    6'b100000, 6'b100001, 6'b100010, 6'b100011 : begin
                        wen_a38 = {1'b0, 1'b0};
                        wen_a37 = {1'b0, 1'b0};
                        wen_a36 = {1'b0, 1'b0};
                        wen_a35 = {1'b0, 1'b0};
                        wen_a34 = {1'b0, 1'b0};
                        wen_a33 = {1'b0, 1'b0};
                        wen_a32 = {1'b0, 1'b0};
                        wen_a31 = {1'b0, 1'b0};
                        wen_a30 = {1'b0, 1'b0};
                        wen_a29 = {1'b0, 1'b0};
                        wen_a28 = {1'b0, 1'b0};
                        wen_a27 = {1'b0, 1'b0};
                        wen_a26 = {1'b0, 1'b0};
                        wen_a25 = {1'b0, 1'b0};
                        wen_a24 = {1'b0, 1'b0};
                        wen_a23 = {1'b0, 1'b0};
                        wen_a22 = {1'b0, 1'b0};
                        wen_a21 = {1'b0, 1'b0};
                        wen_a20 = {1'b0, 1'b0};
                        wen_a19 = {1'b0, 1'b0};
                        wen_a18 = {1'b0, 1'b0};
                        wen_a17 = {1'b0, 1'b0};
                        wen_a16 = {1'b0, 1'b0};
                        wen_a15 = {1'b0, 1'b0};
                        wen_a14 = {1'b0, 1'b0};
                        wen_a13 = {1'b0, 1'b0};
                        wen_a12 = {1'b0, 1'b0};
                        wen_a11 = {1'b0, 1'b0};
                        wen_a10 = {1'b0, 1'b0};
                        wen_a9 = {1'b0, 1'b0};
                        wen_a8 = {1'b0, 1'b0};
                        wen_a7 = {1'b0, 1'b0};
                        wen_a6 = {1'b0, wen};
                        wen_a5 = {1'b0, wen};
                        wen_a4 = {1'b0, wen};
                        wen_a3 = {1'b0, wen};
                        wen_a2 = {1'b0, 1'b0};
                        wen_a1 = {1'b0, 1'b0};
                    end
                    6'b100100, 6'b100101 : begin
                        wen_a38 = {1'b0, 1'b0};
                        wen_a37 = {1'b0, 1'b0};
                        wen_a36 = {1'b0, 1'b0};
                        wen_a35 = {1'b0, 1'b0};
                        wen_a34 = {1'b0, 1'b0};
                        wen_a33 = {1'b0, 1'b0};
                        wen_a32 = {1'b0, 1'b0};
                        wen_a31 = {1'b0, 1'b0};
                        wen_a30 = {1'b0, 1'b0};
                        wen_a29 = {1'b0, 1'b0};
                        wen_a28 = {1'b0, 1'b0};
                        wen_a27 = {1'b0, 1'b0};
                        wen_a26 = {1'b0, 1'b0};
                        wen_a25 = {1'b0, 1'b0};
                        wen_a24 = {1'b0, 1'b0};
                        wen_a23 = {1'b0, 1'b0};
                        wen_a22 = {1'b0, 1'b0};
                        wen_a21 = {1'b0, 1'b0};
                        wen_a20 = {1'b0, 1'b0};
                        wen_a19 = {1'b0, 1'b0};
                        wen_a18 = {1'b0, 1'b0};
                        wen_a17 = {1'b0, 1'b0};
                        wen_a16 = {1'b0, 1'b0};
                        wen_a15 = {1'b0, 1'b0};
                        wen_a14 = {1'b0, 1'b0};
                        wen_a13 = {1'b0, 1'b0};
                        wen_a12 = {1'b0, 1'b0};
                        wen_a11 = {1'b0, 1'b0};
                        wen_a10 = {1'b0, 1'b0};
                        wen_a9 = {1'b0, 1'b0};
                        wen_a8 = {1'b0, 1'b0};
                        wen_a7 = {1'b0, 1'b0};
                        wen_a6 = {1'b0, 1'b0};
                        wen_a5 = {1'b0, 1'b0};
                        wen_a4 = {1'b0, 1'b0};
                        wen_a3 = {1'b0, 1'b0};
                        wen_a2 = {wen, wen};
                        wen_a1 = {wen, wen};
                    end
                    default : begin
                        wen_a38 = {1'b0, 1'b0};
                        wen_a37 = {1'b0, 1'b0};
                        wen_a36 = {1'b0, 1'b0};
                        wen_a35 = {1'b0, 1'b0};
                        wen_a34 = {1'b0, 1'b0};
                        wen_a33 = {1'b0, 1'b0};
                        wen_a32 = {1'b0, 1'b0};
                        wen_a31 = {1'b0, 1'b0};
                        wen_a30 = {1'b0, 1'b0};
                        wen_a29 = {1'b0, 1'b0};
                        wen_a28 = {1'b0, 1'b0};
                        wen_a27 = {1'b0, 1'b0};
                        wen_a26 = {1'b0, 1'b0};
                        wen_a25 = {1'b0, 1'b0};
                        wen_a24 = {1'b0, 1'b0};
                        wen_a23 = {1'b0, 1'b0};
                        wen_a22 = {1'b0, 1'b0};
                        wen_a21 = {1'b0, 1'b0};
                        wen_a20 = {1'b0, 1'b0};
                        wen_a19 = {1'b0, 1'b0};
                        wen_a18 = {1'b0, 1'b0};
                        wen_a17 = {1'b0, 1'b0};
                        wen_a16 = {1'b0, 1'b0};
                        wen_a15 = {1'b0, 1'b0};
                        wen_a14 = {1'b0, 1'b0};
                        wen_a13 = {1'b0, 1'b0};
                        wen_a12 = {1'b0, 1'b0};
                        wen_a11 = {1'b0, 1'b0};
                        wen_a10 = {1'b0, 1'b0};
                        wen_a9 = {1'b0, 1'b0};
                        wen_a8 = {1'b0, 1'b0};
                        wen_a7 = {1'b0, 1'b0};
                        wen_a6 = {1'b0, 1'b0};
                        wen_a5 = {1'b0, 1'b0};
                        wen_a4 = {1'b0, 1'b0};
                        wen_a3 = {1'b0, 1'b0};
                        wen_a2 = {1'b0, 1'b0};
                        wen_a1 = {1'b0, 1'b0};
                    end
                endcase

                case (ckRdAddr[14:9])
                    6'b000000, 6'b000001, 6'b000010, 6'b000011,
                    6'b000100, 6'b000101, 6'b000110, 6'b000111,
                    6'b001000, 6'b001001, 6'b001010, 6'b001011,
                    6'b001100, 6'b001101, 6'b001110, 6'b001111,
                    6'b010000, 6'b010001, 6'b010010, 6'b010011,
                    6'b010100, 6'b010101, 6'b010110, 6'b010111,
                    6'b011000, 6'b011001, 6'b011010, 6'b011011,
                    6'b011100, 6'b011101, 6'b011110, 6'b011111 : begin
                        readData = {
                                        readData38[0],
                                        readData37[0],
                                        readData36[0],
                                        readData35[0],
                                        readData34[0],
                                        readData33[0],
                                        readData32[0],
                                        readData31[0],
                                        readData30[0],
                                        readData29[0],
                                        readData28[0],
                                        readData27[0],
                                        readData26[0],
                                        readData25[0],
                                        readData24[0],
                                        readData23[0],
                                        readData22[0],
                                        readData21[0],
                                        readData20[0],
                                        readData19[0],
                                        readData18[0],
                                        readData17[0],
                                        readData16[0],
                                        readData15[0],
                                        readData14[0],
                                        readData13[0],
                                        readData12[0],
                                        readData11[0],
                                        readData10[0],
                                        readData9[0],
                                        readData8[0],
                                        readData7[0]
                        };
                    end
                    6'b100000, 6'b100001, 6'b100010, 6'b100011 : begin
                        readData = {readData6[7:0],readData5[7:0],readData4[7:0],readData3[7:0]};
                    end
                    6'b100100, 6'b100101 : begin
                        readData = {readData2[16:9],readData2[7:0],readData1[16:9],readData1[7:0]};
                    end
                    default : begin
                        readData = 32'b0;
                    end
                endcase
            end
            19968: begin
                width38 = 3'b000;
                width37 = 3'b000;
                width36 = 3'b000;
                width35 = 3'b000;
                width34 = 3'b000;
                width33 = 3'b000;
                width32 = 3'b000;
                width31 = 3'b000;
                width30 = 3'b000;
                width29 = 3'b000;
                width28 = 3'b000;
                width27 = 3'b000;
                width26 = 3'b000;
                width25 = 3'b000;
                width24 = 3'b000;
                width23 = 3'b000;
                width22 = 3'b000;
                width21 = 3'b000;
                width20 = 3'b000;
                width19 = 3'b000;
                width18 = 3'b000;
                width17 = 3'b000;
                width16 = 3'b000;
                width15 = 3'b000;
                width14 = 3'b000;
                width13 = 3'b000;
                width12 = 3'b000;
                width11 = 3'b000;
                width10 = 3'b000;
                width9 = 3'b000;
                width8 = 3'b000;
                width7 = 3'b000;
                width6 = 3'b011;
                width5 = 3'b011;
                width4 = 3'b011;
                width3 = 3'b011;
                width2 = 3'b100;
                width1 = 3'b100;
                width0 = 3'b101;

                writeAddr38 = {writeAddr[13:0]};
                writeAddr37 = {writeAddr[13:0]};
                writeAddr36 = {writeAddr[13:0]};
                writeAddr35 = {writeAddr[13:0]};
                writeAddr34 = {writeAddr[13:0]};
                writeAddr33 = {writeAddr[13:0]};
                writeAddr32 = {writeAddr[13:0]};
                writeAddr31 = {writeAddr[13:0]};
                writeAddr30 = {writeAddr[13:0]};
                writeAddr29 = {writeAddr[13:0]};
                writeAddr28 = {writeAddr[13:0]};
                writeAddr27 = {writeAddr[13:0]};
                writeAddr26 = {writeAddr[13:0]};
                writeAddr25 = {writeAddr[13:0]};
                writeAddr24 = {writeAddr[13:0]};
                writeAddr23 = {writeAddr[13:0]};
                writeAddr22 = {writeAddr[13:0]};
                writeAddr21 = {writeAddr[13:0]};
                writeAddr20 = {writeAddr[13:0]};
                writeAddr19 = {writeAddr[13:0]};
                writeAddr18 = {writeAddr[13:0]};
                writeAddr17 = {writeAddr[13:0]};
                writeAddr16 = {writeAddr[13:0]};
                writeAddr15 = {writeAddr[13:0]};
                writeAddr14 = {writeAddr[13:0]};
                writeAddr13 = {writeAddr[13:0]};
                writeAddr12 = {writeAddr[13:0]};
                writeAddr11 = {writeAddr[13:0]};
                writeAddr10 = {writeAddr[13:0]};
                writeAddr9 = {writeAddr[13:0]};
                writeAddr8 = {writeAddr[13:0]};
                writeAddr7 = {writeAddr[13:0]};
                writeAddr6 = {writeAddr[10:0], 3'b0};
                writeAddr5 = {writeAddr[10:0], 3'b0};
                writeAddr4 = {writeAddr[10:0], 3'b0};
                writeAddr3 = {writeAddr[10:0], 3'b0};
                writeAddr2 = {writeAddr[9:0], 4'b0};
                writeAddr1 = {writeAddr[9:0], 4'b0};
                writeAddr0 = {writeAddr[8:0], 5'b0};

                readAddr38 = {writeAddr[13:0]};
                readAddr37 = {writeAddr[13:0]};
                readAddr36 = {writeAddr[13:0]};
                readAddr35 = {writeAddr[13:0]};
                readAddr34 = {writeAddr[13:0]};
                readAddr33 = {writeAddr[13:0]};
                readAddr32 = {writeAddr[13:0]};
                readAddr31 = {writeAddr[13:0]};
                readAddr30 = {writeAddr[13:0]};
                readAddr29 = {writeAddr[13:0]};
                readAddr28 = {writeAddr[13:0]};
                readAddr27 = {writeAddr[13:0]};
                readAddr26 = {writeAddr[13:0]};
                readAddr25 = {writeAddr[13:0]};
                readAddr24 = {writeAddr[13:0]};
                readAddr23 = {writeAddr[13:0]};
                readAddr22 = {writeAddr[13:0]};
                readAddr21 = {writeAddr[13:0]};
                readAddr20 = {writeAddr[13:0]};
                readAddr19 = {writeAddr[13:0]};
                readAddr18 = {writeAddr[13:0]};
                readAddr17 = {writeAddr[13:0]};
                readAddr16 = {writeAddr[13:0]};
                readAddr15 = {writeAddr[13:0]};
                readAddr14 = {writeAddr[13:0]};
                readAddr13 = {writeAddr[13:0]};
                readAddr12 = {writeAddr[13:0]};
                readAddr11 = {writeAddr[13:0]};
                readAddr10 = {writeAddr[13:0]};
                readAddr9 = {writeAddr[13:0]};
                readAddr8 = {writeAddr[13:0]};
                readAddr7 = {writeAddr[13:0]};
                readAddr6  = {readAddr[10:0],  3'b0};
                readAddr5  = {readAddr[10:0],  3'b0};
                readAddr4  = {readAddr[10:0],  3'b0};
                readAddr3  = {readAddr[10:0],  3'b0};
                readAddr2  = {readAddr[9:0],  4'b0};
                readAddr1  = {readAddr[9:0],  4'b0};
                readAddr0  = {readAddr[8:0],  5'b0};

                writeData38 = {17'b0, writeData[31]};
                writeData37 = {17'b0, writeData[30]};
                writeData36 = {17'b0, writeData[29]};
                writeData35 = {17'b0, writeData[28]};
                writeData34 = {17'b0, writeData[27]};
                writeData33 = {17'b0, writeData[26]};
                writeData32 = {17'b0, writeData[25]};
                writeData31 = {17'b0, writeData[24]};
                writeData30 = {17'b0, writeData[23]};
                writeData29 = {17'b0, writeData[22]};
                writeData28 = {17'b0, writeData[21]};
                writeData27 = {17'b0, writeData[20]};
                writeData26 = {17'b0, writeData[19]};
                writeData25 = {17'b0, writeData[18]};
                writeData24 = {17'b0, writeData[17]};
                writeData23 = {17'b0, writeData[16]};
                writeData22 = {17'b0, writeData[15]};
                writeData21 = {17'b0, writeData[14]};
                writeData20 = {17'b0, writeData[13]};
                writeData19 = {17'b0, writeData[12]};
                writeData18 = {17'b0, writeData[11]};
                writeData17 = {17'b0, writeData[10]};
                writeData16 = {17'b0, writeData[9]};
                writeData15 = {17'b0, writeData[8]};
                writeData14 = {17'b0, writeData[7]};
                writeData13 = {17'b0, writeData[6]};
                writeData12 = {17'b0, writeData[5]};
                writeData11 = {17'b0, writeData[4]};
                writeData10 = {17'b0, writeData[3]};
                writeData9 = {17'b0, writeData[2]};
                writeData8 = {17'b0, writeData[1]};
                writeData7 = {17'b0, writeData[0]};
                writeData6 = {10'b0, writeData[31:24]};
                writeData5 = {10'b0, writeData[23:16]};
                writeData4 = {10'b0, writeData[15:8]};
                writeData3 = {10'b0, writeData[7:0]};
                writeData2 = {1'b0, writeData[31:24], 1'b0, writeData[23:16]};
                writeData1 = {1'b0, writeData[15:8], 1'b0, writeData[7:0]};
                writeData0 = {1'b0, writeData[31:24], 1'b0, writeData[23:16], 1'b0, writeData[15:8], 1'b0, writeData[7:0]};

                case (writeAddr[14:9])
                    6'b000000, 6'b000001, 6'b000010, 6'b000011,
                    6'b000100, 6'b000101, 6'b000110, 6'b000111,
                    6'b001000, 6'b001001, 6'b001010, 6'b001011,
                    6'b001100, 6'b001101, 6'b001110, 6'b001111,
                    6'b010000, 6'b010001, 6'b010010, 6'b010011,
                    6'b010100, 6'b010101, 6'b010110, 6'b010111,
                    6'b011000, 6'b011001, 6'b011010, 6'b011011,
                    6'b011100, 6'b011101, 6'b011110, 6'b011111 : begin
                        wen_a38 = {1'b0, wen};
                        wen_a37 = {1'b0, wen};
                        wen_a36 = {1'b0, wen};
                        wen_a35 = {1'b0, wen};
                        wen_a34 = {1'b0, wen};
                        wen_a33 = {1'b0, wen};
                        wen_a32 = {1'b0, wen};
                        wen_a31 = {1'b0, wen};
                        wen_a30 = {1'b0, wen};
                        wen_a29 = {1'b0, wen};
                        wen_a28 = {1'b0, wen};
                        wen_a27 = {1'b0, wen};
                        wen_a26 = {1'b0, wen};
                        wen_a25 = {1'b0, wen};
                        wen_a24 = {1'b0, wen};
                        wen_a23 = {1'b0, wen};
                        wen_a22 = {1'b0, wen};
                        wen_a21 = {1'b0, wen};
                        wen_a20 = {1'b0, wen};
                        wen_a19 = {1'b0, wen};
                        wen_a18 = {1'b0, wen};
                        wen_a17 = {1'b0, wen};
                        wen_a16 = {1'b0, wen};
                        wen_a15 = {1'b0, wen};
                        wen_a14 = {1'b0, wen};
                        wen_a13 = {1'b0, wen};
                        wen_a12 = {1'b0, wen};
                        wen_a11 = {1'b0, wen};
                        wen_a10 = {1'b0, wen};
                        wen_a9 = {1'b0, wen};
                        wen_a8 = {1'b0, wen};
                        wen_a7 = {1'b0, wen};
                        wen_a6 = {1'b0, 1'b0};
                        wen_a5 = {1'b0, 1'b0};
                        wen_a4 = {1'b0, 1'b0};
                        wen_a3 = {1'b0, 1'b0};
                        wen_a2 = {1'b0, 1'b0};
                        wen_a1 = {1'b0, 1'b0};
                        wen_a0 = {1'b0, 1'b0};
                        wen_b0 = {1'b0, 1'b0};
                    end
                    6'b100000, 6'b100001, 6'b100010, 6'b100011 : begin
                        wen_a38 = {1'b0, 1'b0};
                        wen_a37 = {1'b0, 1'b0};
                        wen_a36 = {1'b0, 1'b0};
                        wen_a35 = {1'b0, 1'b0};
                        wen_a34 = {1'b0, 1'b0};
                        wen_a33 = {1'b0, 1'b0};
                        wen_a32 = {1'b0, 1'b0};
                        wen_a31 = {1'b0, 1'b0};
                        wen_a30 = {1'b0, 1'b0};
                        wen_a29 = {1'b0, 1'b0};
                        wen_a28 = {1'b0, 1'b0};
                        wen_a27 = {1'b0, 1'b0};
                        wen_a26 = {1'b0, 1'b0};
                        wen_a25 = {1'b0, 1'b0};
                        wen_a24 = {1'b0, 1'b0};
                        wen_a23 = {1'b0, 1'b0};
                        wen_a22 = {1'b0, 1'b0};
                        wen_a21 = {1'b0, 1'b0};
                        wen_a20 = {1'b0, 1'b0};
                        wen_a19 = {1'b0, 1'b0};
                        wen_a18 = {1'b0, 1'b0};
                        wen_a17 = {1'b0, 1'b0};
                        wen_a16 = {1'b0, 1'b0};
                        wen_a15 = {1'b0, 1'b0};
                        wen_a14 = {1'b0, 1'b0};
                        wen_a13 = {1'b0, 1'b0};
                        wen_a12 = {1'b0, 1'b0};
                        wen_a11 = {1'b0, 1'b0};
                        wen_a10 = {1'b0, 1'b0};
                        wen_a9 = {1'b0, 1'b0};
                        wen_a8 = {1'b0, 1'b0};
                        wen_a7 = {1'b0, 1'b0};
                        wen_a6 = {1'b0, wen};
                        wen_a5 = {1'b0, wen};
                        wen_a4 = {1'b0, wen};
                        wen_a3 = {1'b0, wen};
                        wen_a2 = {1'b0, 1'b0};
                        wen_a1 = {1'b0, 1'b0};
                        wen_a0 = {1'b0, 1'b0};
                        wen_b0 = {1'b0, 1'b0};
                    end
                    6'b100100, 6'b100101 : begin
                        wen_a38 = {1'b0, 1'b0};
                        wen_a37 = {1'b0, 1'b0};
                        wen_a36 = {1'b0, 1'b0};
                        wen_a35 = {1'b0, 1'b0};
                        wen_a34 = {1'b0, 1'b0};
                        wen_a33 = {1'b0, 1'b0};
                        wen_a32 = {1'b0, 1'b0};
                        wen_a31 = {1'b0, 1'b0};
                        wen_a30 = {1'b0, 1'b0};
                        wen_a29 = {1'b0, 1'b0};
                        wen_a28 = {1'b0, 1'b0};
                        wen_a27 = {1'b0, 1'b0};
                        wen_a26 = {1'b0, 1'b0};
                        wen_a25 = {1'b0, 1'b0};
                        wen_a24 = {1'b0, 1'b0};
                        wen_a23 = {1'b0, 1'b0};
                        wen_a22 = {1'b0, 1'b0};
                        wen_a21 = {1'b0, 1'b0};
                        wen_a20 = {1'b0, 1'b0};
                        wen_a19 = {1'b0, 1'b0};
                        wen_a18 = {1'b0, 1'b0};
                        wen_a17 = {1'b0, 1'b0};
                        wen_a16 = {1'b0, 1'b0};
                        wen_a15 = {1'b0, 1'b0};
                        wen_a14 = {1'b0, 1'b0};
                        wen_a13 = {1'b0, 1'b0};
                        wen_a12 = {1'b0, 1'b0};
                        wen_a11 = {1'b0, 1'b0};
                        wen_a10 = {1'b0, 1'b0};
                        wen_a9 = {1'b0, 1'b0};
                        wen_a8 = {1'b0, 1'b0};
                        wen_a7 = {1'b0, 1'b0};
                        wen_a6 = {1'b0, 1'b0};
                        wen_a5 = {1'b0, 1'b0};
                        wen_a4 = {1'b0, 1'b0};
                        wen_a3 = {1'b0, 1'b0};
                        wen_a2 = {wen, wen};
                        wen_a1 = {wen, wen};
                        wen_a0 = {1'b0, 1'b0};
                        wen_b0 = {1'b0, 1'b0};
                    end
                    6'b100110: begin
                        wen_a38 = {1'b0, 1'b0};
                        wen_a37 = {1'b0, 1'b0};
                        wen_a36 = {1'b0, 1'b0};
                        wen_a35 = {1'b0, 1'b0};
                        wen_a34 = {1'b0, 1'b0};
                        wen_a33 = {1'b0, 1'b0};
                        wen_a32 = {1'b0, 1'b0};
                        wen_a31 = {1'b0, 1'b0};
                        wen_a30 = {1'b0, 1'b0};
                        wen_a29 = {1'b0, 1'b0};
                        wen_a28 = {1'b0, 1'b0};
                        wen_a27 = {1'b0, 1'b0};
                        wen_a26 = {1'b0, 1'b0};
                        wen_a25 = {1'b0, 1'b0};
                        wen_a24 = {1'b0, 1'b0};
                        wen_a23 = {1'b0, 1'b0};
                        wen_a22 = {1'b0, 1'b0};
                        wen_a21 = {1'b0, 1'b0};
                        wen_a20 = {1'b0, 1'b0};
                        wen_a19 = {1'b0, 1'b0};
                        wen_a18 = {1'b0, 1'b0};
                        wen_a17 = {1'b0, 1'b0};
                        wen_a16 = {1'b0, 1'b0};
                        wen_a15 = {1'b0, 1'b0};
                        wen_a14 = {1'b0, 1'b0};
                        wen_a13 = {1'b0, 1'b0};
                        wen_a12 = {1'b0, 1'b0};
                        wen_a11 = {1'b0, 1'b0};
                        wen_a10 = {1'b0, 1'b0};
                        wen_a9 = {1'b0, 1'b0};
                        wen_a8 = {1'b0, 1'b0};
                        wen_a7 = {1'b0, 1'b0};
                        wen_a6 = {1'b0, 1'b0};
                        wen_a5 = {1'b0, 1'b0};
                        wen_a4 = {1'b0, 1'b0};
                        wen_a3 = {1'b0, 1'b0};
                        wen_a2 = {1'b0, 1'b0};
                        wen_a1 = {1'b0, 1'b0};
                        wen_a0 = {wen, wen};
                        wen_b0 = {wen, wen};
                    end
                    default : begin
                        wen_a38 = {1'b0, 1'b0};
                        wen_a37 = {1'b0, 1'b0};
                        wen_a36 = {1'b0, 1'b0};
                        wen_a35 = {1'b0, 1'b0};
                        wen_a34 = {1'b0, 1'b0};
                        wen_a33 = {1'b0, 1'b0};
                        wen_a32 = {1'b0, 1'b0};
                        wen_a31 = {1'b0, 1'b0};
                        wen_a30 = {1'b0, 1'b0};
                        wen_a29 = {1'b0, 1'b0};
                        wen_a28 = {1'b0, 1'b0};
                        wen_a27 = {1'b0, 1'b0};
                        wen_a26 = {1'b0, 1'b0};
                        wen_a25 = {1'b0, 1'b0};
                        wen_a24 = {1'b0, 1'b0};
                        wen_a23 = {1'b0, 1'b0};
                        wen_a22 = {1'b0, 1'b0};
                        wen_a21 = {1'b0, 1'b0};
                        wen_a20 = {1'b0, 1'b0};
                        wen_a19 = {1'b0, 1'b0};
                        wen_a18 = {1'b0, 1'b0};
                        wen_a17 = {1'b0, 1'b0};
                        wen_a16 = {1'b0, 1'b0};
                        wen_a15 = {1'b0, 1'b0};
                        wen_a14 = {1'b0, 1'b0};
                        wen_a13 = {1'b0, 1'b0};
                        wen_a12 = {1'b0, 1'b0};
                        wen_a11 = {1'b0, 1'b0};
                        wen_a10 = {1'b0, 1'b0};
                        wen_a9 = {1'b0, 1'b0};
                        wen_a8 = {1'b0, 1'b0};
                        wen_a7 = {1'b0, 1'b0};
                        wen_a6 = {1'b0, 1'b0};
                        wen_a5 = {1'b0, 1'b0};
                        wen_a4 = {1'b0, 1'b0};
                        wen_a3 = {1'b0, 1'b0};
                        wen_a2 = {1'b0, 1'b0};
                        wen_a1 = {1'b0, 1'b0};
                        wen_a0 = {1'b0, 1'b0};
                        wen_b0 = {1'b0, 1'b0};
                    end
                endcase

                case (ckRdAddr[14:9])
                    6'b000000, 6'b000001, 6'b000010, 6'b000011,
                    6'b000100, 6'b000101, 6'b000110, 6'b000111,
                    6'b001000, 6'b001001, 6'b001010, 6'b001011,
                    6'b001100, 6'b001101, 6'b001110, 6'b001111,
                    6'b010000, 6'b010001, 6'b010010, 6'b010011,
                    6'b010100, 6'b010101, 6'b010110, 6'b010111,
                    6'b011000, 6'b011001, 6'b011010, 6'b011011,
                    6'b011100, 6'b011101, 6'b011110, 6'b011111 : begin
                        readData = {
                                        readData38[0],
                                        readData37[0],
                                        readData36[0],
                                        readData35[0],
                                        readData34[0],
                                        readData33[0],
                                        readData32[0],
                                        readData31[0],
                                        readData30[0],
                                        readData29[0],
                                        readData28[0],
                                        readData27[0],
                                        readData26[0],
                                        readData25[0],
                                        readData24[0],
                                        readData23[0],
                                        readData22[0],
                                        readData21[0],
                                        readData20[0],
                                        readData19[0],
                                        readData18[0],
                                        readData17[0],
                                        readData16[0],
                                        readData15[0],
                                        readData14[0],
                                        readData13[0],
                                        readData12[0],
                                        readData11[0],
                                        readData10[0],
                                        readData9[0],
                                        readData8[0],
                                        readData7[0]
                        };
                    end
                    6'b100000, 6'b100001, 6'b100010, 6'b100011 : begin
                        readData = {readData6[7:0],readData5[7:0],readData4[7:0],readData3[7:0]};
                    end
                    6'b100100, 6'b100101 : begin
                        readData = {readData2[16:9],readData2[7:0],readData1[16:9],readData1[7:0]};
                    end
                    6'b100110: begin
                        readData = {readData0[34:27],readData0[25:18],readData0[16:9],readData0[7:0]};
                    end
                    default : begin
                        readData = 32'b0;
                    end
                endcase
            end
            20480: begin
                width40 = 3'b000;
                width39 = 3'b000;
                width38 = 3'b000;
                width37 = 3'b000;
                width36 = 3'b000;
                width35 = 3'b000;
                width34 = 3'b000;
                width33 = 3'b000;
                width32 = 3'b000;
                width31 = 3'b000;
                width30 = 3'b000;
                width29 = 3'b000;
                width28 = 3'b000;
                width27 = 3'b000;
                width26 = 3'b000;
                width25 = 3'b000;
                width24 = 3'b000;
                width23 = 3'b000;
                width22 = 3'b000;
                width21 = 3'b000;
                width20 = 3'b000;
                width19 = 3'b000;
                width18 = 3'b000;
                width17 = 3'b000;
                width16 = 3'b000;
                width15 = 3'b000;
                width14 = 3'b000;
                width13 = 3'b000;
                width12 = 3'b000;
                width11 = 3'b000;
                width10 = 3'b000;
                width9 = 3'b000;
                width8 = 3'b010;
                width7 = 3'b010;
                width6 = 3'b010;
                width5 = 3'b010;
                width4 = 3'b010;
                width3 = 3'b010;
                width2 = 3'b010;
                width1 = 3'b010;

                writeAddr40 = {writeAddr[13:0]};
                writeAddr39 = {writeAddr[13:0]};
                writeAddr38 = {writeAddr[13:0]};
                writeAddr37 = {writeAddr[13:0]};
                writeAddr36 = {writeAddr[13:0]};
                writeAddr35 = {writeAddr[13:0]};
                writeAddr34 = {writeAddr[13:0]};
                writeAddr33 = {writeAddr[13:0]};
                writeAddr32 = {writeAddr[13:0]};
                writeAddr31 = {writeAddr[13:0]};
                writeAddr30 = {writeAddr[13:0]};
                writeAddr29 = {writeAddr[13:0]};
                writeAddr28 = {writeAddr[13:0]};
                writeAddr27 = {writeAddr[13:0]};
                writeAddr26 = {writeAddr[13:0]};
                writeAddr25 = {writeAddr[13:0]};
                writeAddr24 = {writeAddr[13:0]};
                writeAddr23 = {writeAddr[13:0]};
                writeAddr22 = {writeAddr[13:0]};
                writeAddr21 = {writeAddr[13:0]};
                writeAddr20 = {writeAddr[13:0]};
                writeAddr19 = {writeAddr[13:0]};
                writeAddr18 = {writeAddr[13:0]};
                writeAddr17 = {writeAddr[13:0]};
                writeAddr16 = {writeAddr[13:0]};
                writeAddr15 = {writeAddr[13:0]};
                writeAddr14 = {writeAddr[13:0]};
                writeAddr13 = {writeAddr[13:0]};
                writeAddr12 = {writeAddr[13:0]};
                writeAddr11 = {writeAddr[13:0]};
                writeAddr10 = {writeAddr[13:0]};
                writeAddr9 = {writeAddr[13:0]};
                writeAddr8 = {writeAddr[11:0], 2'b0};
                writeAddr7 = {writeAddr[11:0], 2'b0};
                writeAddr6 = {writeAddr[11:0], 2'b0};
                writeAddr5 = {writeAddr[11:0], 2'b0};
                writeAddr4 = {writeAddr[11:0], 2'b0};
                writeAddr3 = {writeAddr[11:0], 2'b0};
                writeAddr2 = {writeAddr[11:0], 2'b0};
                writeAddr1 = {writeAddr[11:0], 2'b0};

                readAddr40 = {writeAddr[13:0]};
                readAddr39 = {writeAddr[13:0]};
                readAddr38 = {writeAddr[13:0]};
                readAddr37 = {writeAddr[13:0]};
                readAddr36 = {writeAddr[13:0]};
                readAddr35 = {writeAddr[13:0]};
                readAddr34 = {writeAddr[13:0]};
                readAddr33 = {writeAddr[13:0]};
                readAddr32 = {writeAddr[13:0]};
                readAddr31 = {writeAddr[13:0]};
                readAddr30 = {writeAddr[13:0]};
                readAddr29 = {writeAddr[13:0]};
                readAddr28 = {writeAddr[13:0]};
                readAddr27 = {writeAddr[13:0]};
                readAddr26 = {writeAddr[13:0]};
                readAddr25 = {writeAddr[13:0]};
                readAddr24 = {writeAddr[13:0]};
                readAddr23 = {writeAddr[13:0]};
                readAddr22 = {writeAddr[13:0]};
                readAddr21 = {writeAddr[13:0]};
                readAddr20 = {writeAddr[13:0]};
                readAddr19 = {writeAddr[13:0]};
                readAddr18 = {writeAddr[13:0]};
                readAddr17 = {writeAddr[13:0]};
                readAddr16 = {writeAddr[13:0]};
                readAddr15 = {writeAddr[13:0]};
                readAddr14 = {writeAddr[13:0]};
                readAddr13 = {writeAddr[13:0]};
                readAddr12 = {writeAddr[13:0]};
                readAddr11 = {writeAddr[13:0]};
                readAddr10 = {writeAddr[13:0]};
                readAddr9 = {writeAddr[13:0]};
                readAddr8  = {readAddr[11:0],  2'b0};
                readAddr7  = {readAddr[11:0],  2'b0};
                readAddr6  = {readAddr[11:0],  2'b0};
                readAddr5  = {readAddr[11:0],  2'b0};
                readAddr4  = {readAddr[11:0],  2'b0};
                readAddr3  = {readAddr[11:0],  2'b0};
                readAddr2  = {readAddr[11:0],  2'b0};
                readAddr1  = {readAddr[11:0],  2'b0};

                writeData40 = {17'b0, writeData[31]};
                writeData39 = {17'b0, writeData[30]};
                writeData38 = {17'b0, writeData[29]};
                writeData37 = {17'b0, writeData[28]};
                writeData36 = {17'b0, writeData[27]};
                writeData35 = {17'b0, writeData[26]};
                writeData34 = {17'b0, writeData[25]};
                writeData33 = {17'b0, writeData[24]};
                writeData32 = {17'b0, writeData[23]};
                writeData31 = {17'b0, writeData[22]};
                writeData30 = {17'b0, writeData[21]};
                writeData29 = {17'b0, writeData[20]};
                writeData28 = {17'b0, writeData[19]};
                writeData27 = {17'b0, writeData[18]};
                writeData26 = {17'b0, writeData[17]};
                writeData25 = {17'b0, writeData[16]};
                writeData24 = {17'b0, writeData[15]};
                writeData23 = {17'b0, writeData[14]};
                writeData22 = {17'b0, writeData[13]};
                writeData21 = {17'b0, writeData[12]};
                writeData20 = {17'b0, writeData[11]};
                writeData19 = {17'b0, writeData[10]};
                writeData18 = {17'b0, writeData[9]};
                writeData17 = {17'b0, writeData[8]};
                writeData16 = {17'b0, writeData[7]};
                writeData15 = {17'b0, writeData[6]};
                writeData14 = {17'b0, writeData[5]};
                writeData13 = {17'b0, writeData[4]};
                writeData12 = {17'b0, writeData[3]};
                writeData11 = {17'b0, writeData[2]};
                writeData10 = {17'b0, writeData[1]};
                writeData9 = {17'b0, writeData[0]};
                writeData8 = {14'b0, writeData[31:28]};
                writeData7 = {14'b0, writeData[27:24]};
                writeData6 = {14'b0, writeData[23:20]};
                writeData5 = {14'b0, writeData[19:16]};
                writeData4 = {14'b0, writeData[15:12]};
                writeData3 = {14'b0, writeData[11:8]};
                writeData2 = {14'b0, writeData[7:4]};
                writeData1 = {14'b0, writeData[3:0]};

                case (writeAddr[14:9])
                    6'b000000, 6'b000001, 6'b000010, 6'b000011,
                    6'b000100, 6'b000101, 6'b000110, 6'b000111,
                    6'b001000, 6'b001001, 6'b001010, 6'b001011,
                    6'b001100, 6'b001101, 6'b001110, 6'b001111,
                    6'b010000, 6'b010001, 6'b010010, 6'b010011,
                    6'b010100, 6'b010101, 6'b010110, 6'b010111,
                    6'b011000, 6'b011001, 6'b011010, 6'b011011,
                    6'b011100, 6'b011101, 6'b011110, 6'b011111 : begin
                        wen_a40 = {1'b0, wen};
                        wen_a39 = {1'b0, wen};
                        wen_a38 = {1'b0, wen};
                        wen_a37 = {1'b0, wen};
                        wen_a36 = {1'b0, wen};
                        wen_a35 = {1'b0, wen};
                        wen_a34 = {1'b0, wen};
                        wen_a33 = {1'b0, wen};
                        wen_a32 = {1'b0, wen};
                        wen_a31 = {1'b0, wen};
                        wen_a30 = {1'b0, wen};
                        wen_a29 = {1'b0, wen};
                        wen_a28 = {1'b0, wen};
                        wen_a27 = {1'b0, wen};
                        wen_a26 = {1'b0, wen};
                        wen_a25 = {1'b0, wen};
                        wen_a24 = {1'b0, wen};
                        wen_a23 = {1'b0, wen};
                        wen_a22 = {1'b0, wen};
                        wen_a21 = {1'b0, wen};
                        wen_a20 = {1'b0, wen};
                        wen_a19 = {1'b0, wen};
                        wen_a18 = {1'b0, wen};
                        wen_a17 = {1'b0, wen};
                        wen_a16 = {1'b0, wen};
                        wen_a15 = {1'b0, wen};
                        wen_a14 = {1'b0, wen};
                        wen_a13 = {1'b0, wen};
                        wen_a12 = {1'b0, wen};
                        wen_a11 = {1'b0, wen};
                        wen_a10 = {1'b0, wen};
                        wen_a9 = {1'b0, wen};
                        wen_a8 = {1'b0, 1'b0};
                        wen_a7 = {1'b0, 1'b0};
                        wen_a6 = {1'b0, 1'b0};
                        wen_a5 = {1'b0, 1'b0};
                        wen_a4 = {1'b0, 1'b0};
                        wen_a3 = {1'b0, 1'b0};
                        wen_a2 = {1'b0, 1'b0};
                        wen_a1 = {1'b0, 1'b0};
                    end
                    6'b100000, 6'b100001, 6'b100010, 6'b100011,
                    6'b100100, 6'b100101, 6'b100110, 6'b100111: begin
                        wen_a40 = {1'b0, 1'b0};
                        wen_a39 = {1'b0, 1'b0};
                        wen_a38 = {1'b0, 1'b0};
                        wen_a37 = {1'b0, 1'b0};
                        wen_a36 = {1'b0, 1'b0};
                        wen_a35 = {1'b0, 1'b0};
                        wen_a34 = {1'b0, 1'b0};
                        wen_a33 = {1'b0, 1'b0};
                        wen_a32 = {1'b0, 1'b0};
                        wen_a31 = {1'b0, 1'b0};
                        wen_a30 = {1'b0, 1'b0};
                        wen_a29 = {1'b0, 1'b0};
                        wen_a28 = {1'b0, 1'b0};
                        wen_a27 = {1'b0, 1'b0};
                        wen_a26 = {1'b0, 1'b0};
                        wen_a25 = {1'b0, 1'b0};
                        wen_a24 = {1'b0, 1'b0};
                        wen_a23 = {1'b0, 1'b0};
                        wen_a22 = {1'b0, 1'b0};
                        wen_a21 = {1'b0, 1'b0};
                        wen_a20 = {1'b0, 1'b0};
                        wen_a19 = {1'b0, 1'b0};
                        wen_a18 = {1'b0, 1'b0};
                        wen_a17 = {1'b0, 1'b0};
                        wen_a16 = {1'b0, 1'b0};
                        wen_a15 = {1'b0, 1'b0};
                        wen_a14 = {1'b0, 1'b0};
                        wen_a13 = {1'b0, 1'b0};
                        wen_a12 = {1'b0, 1'b0};
                        wen_a11 = {1'b0, 1'b0};
                        wen_a10 = {1'b0, 1'b0};
                        wen_a9 = {1'b0, 1'b0};
                        wen_a8 = {1'b0, wen};
                        wen_a7 = {1'b0, wen};
                        wen_a6 = {1'b0, wen};
                        wen_a5 = {1'b0, wen};
                        wen_a4 = {1'b0, wen};
                        wen_a3 = {1'b0, wen};
                        wen_a2 = {1'b0, wen};
                        wen_a1 = {1'b0, wen};
                    end
                    default : begin
                        wen_a40 = {1'b0, 1'b0};
                        wen_a39 = {1'b0, 1'b0};
                        wen_a38 = {1'b0, 1'b0};
                        wen_a37 = {1'b0, 1'b0};
                        wen_a36 = {1'b0, 1'b0};
                        wen_a35 = {1'b0, 1'b0};
                        wen_a34 = {1'b0, 1'b0};
                        wen_a33 = {1'b0, 1'b0};
                        wen_a32 = {1'b0, 1'b0};
                        wen_a31 = {1'b0, 1'b0};
                        wen_a30 = {1'b0, 1'b0};
                        wen_a29 = {1'b0, 1'b0};
                        wen_a28 = {1'b0, 1'b0};
                        wen_a27 = {1'b0, 1'b0};
                        wen_a26 = {1'b0, 1'b0};
                        wen_a25 = {1'b0, 1'b0};
                        wen_a24 = {1'b0, 1'b0};
                        wen_a23 = {1'b0, 1'b0};
                        wen_a22 = {1'b0, 1'b0};
                        wen_a21 = {1'b0, 1'b0};
                        wen_a20 = {1'b0, 1'b0};
                        wen_a19 = {1'b0, 1'b0};
                        wen_a18 = {1'b0, 1'b0};
                        wen_a17 = {1'b0, 1'b0};
                        wen_a16 = {1'b0, 1'b0};
                        wen_a15 = {1'b0, 1'b0};
                        wen_a14 = {1'b0, 1'b0};
                        wen_a13 = {1'b0, 1'b0};
                        wen_a12 = {1'b0, 1'b0};
                        wen_a11 = {1'b0, 1'b0};
                        wen_a10 = {1'b0, 1'b0};
                        wen_a9 = {1'b0, 1'b0};
                        wen_a8 = {1'b0, 1'b0};
                        wen_a7 = {1'b0, 1'b0};
                        wen_a6 = {1'b0, 1'b0};
                        wen_a5 = {1'b0, 1'b0};
                        wen_a4 = {1'b0, 1'b0};
                        wen_a3 = {1'b0, 1'b0};
                        wen_a2 = {1'b0, 1'b0};
                        wen_a1 = {1'b0, 1'b0};
                    end
                endcase

                case (ckRdAddr[14:9])
                    6'b000000, 6'b000001, 6'b000010, 6'b000011,
                    6'b000100, 6'b000101, 6'b000110, 6'b000111,
                    6'b001000, 6'b001001, 6'b001010, 6'b001011,
                    6'b001100, 6'b001101, 6'b001110, 6'b001111,
                    6'b010000, 6'b010001, 6'b010010, 6'b010011,
                    6'b010100, 6'b010101, 6'b010110, 6'b010111,
                    6'b011000, 6'b011001, 6'b011010, 6'b011011,
                    6'b011100, 6'b011101, 6'b011110, 6'b011111 : begin
                        readData = {
                                        readData40[0],
                                        readData39[0],
                                        readData38[0],
                                        readData37[0],
                                        readData36[0],
                                        readData35[0],
                                        readData34[0],
                                        readData33[0],
                                        readData32[0],
                                        readData31[0],
                                        readData30[0],
                                        readData29[0],
                                        readData28[0],
                                        readData27[0],
                                        readData26[0],
                                        readData25[0],
                                        readData24[0],
                                        readData23[0],
                                        readData22[0],
                                        readData21[0],
                                        readData20[0],
                                        readData19[0],
                                        readData18[0],
                                        readData17[0],
                                        readData16[0],
                                        readData15[0],
                                        readData14[0],
                                        readData13[0],
                                        readData12[0],
                                        readData11[0],
                                        readData10[0],
                                        readData9[0]
                        };
                    end
                    6'b100000, 6'b100001, 6'b100010, 6'b100011,
                    6'b100100, 6'b100101, 6'b100110, 6'b100111: begin
                        readData = {
                                        readData8[3:0],
                                        readData7[3:0],
                                        readData6[3:0],
                                        readData5[3:0],
                                        readData4[3:0],
                                        readData3[3:0],
                                        readData2[3:0],
                                        readData1[3:0]
                        };
                    end
                    default : begin
                        readData = 32'b0;
                    end
                endcase
            end
            20992: begin
                width40 = 3'b000;
                width39 = 3'b000;
                width38 = 3'b000;
                width37 = 3'b000;
                width36 = 3'b000;
                width35 = 3'b000;
                width34 = 3'b000;
                width33 = 3'b000;
                width32 = 3'b000;
                width31 = 3'b000;
                width30 = 3'b000;
                width29 = 3'b000;
                width28 = 3'b000;
                width27 = 3'b000;
                width26 = 3'b000;
                width25 = 3'b000;
                width24 = 3'b000;
                width23 = 3'b000;
                width22 = 3'b000;
                width21 = 3'b000;
                width20 = 3'b000;
                width19 = 3'b000;
                width18 = 3'b000;
                width17 = 3'b000;
                width16 = 3'b000;
                width15 = 3'b000;
                width14 = 3'b000;
                width13 = 3'b000;
                width12 = 3'b000;
                width11 = 3'b000;
                width10 = 3'b000;
                width9 = 3'b000;
                width8 = 3'b010;
                width7 = 3'b010;
                width6 = 3'b010;
                width5 = 3'b010;
                width4 = 3'b010;
                width3 = 3'b010;
                width2 = 3'b010;
                width1 = 3'b010;
                width0 = 3'b101;

                writeAddr40 = {writeAddr[13:0]};
                writeAddr39 = {writeAddr[13:0]};
                writeAddr38 = {writeAddr[13:0]};
                writeAddr37 = {writeAddr[13:0]};
                writeAddr36 = {writeAddr[13:0]};
                writeAddr35 = {writeAddr[13:0]};
                writeAddr34 = {writeAddr[13:0]};
                writeAddr33 = {writeAddr[13:0]};
                writeAddr32 = {writeAddr[13:0]};
                writeAddr31 = {writeAddr[13:0]};
                writeAddr30 = {writeAddr[13:0]};
                writeAddr29 = {writeAddr[13:0]};
                writeAddr28 = {writeAddr[13:0]};
                writeAddr27 = {writeAddr[13:0]};
                writeAddr26 = {writeAddr[13:0]};
                writeAddr25 = {writeAddr[13:0]};
                writeAddr24 = {writeAddr[13:0]};
                writeAddr23 = {writeAddr[13:0]};
                writeAddr22 = {writeAddr[13:0]};
                writeAddr21 = {writeAddr[13:0]};
                writeAddr20 = {writeAddr[13:0]};
                writeAddr19 = {writeAddr[13:0]};
                writeAddr18 = {writeAddr[13:0]};
                writeAddr17 = {writeAddr[13:0]};
                writeAddr16 = {writeAddr[13:0]};
                writeAddr15 = {writeAddr[13:0]};
                writeAddr14 = {writeAddr[13:0]};
                writeAddr13 = {writeAddr[13:0]};
                writeAddr12 = {writeAddr[13:0]};
                writeAddr11 = {writeAddr[13:0]};
                writeAddr10 = {writeAddr[13:0]};
                writeAddr9 = {writeAddr[13:0]};
                writeAddr8 = {writeAddr[11:0], 2'b0};
                writeAddr7 = {writeAddr[11:0], 2'b0};
                writeAddr6 = {writeAddr[11:0], 2'b0};
                writeAddr5 = {writeAddr[11:0], 2'b0};
                writeAddr4 = {writeAddr[11:0], 2'b0};
                writeAddr3 = {writeAddr[11:0], 2'b0};
                writeAddr2 = {writeAddr[11:0], 2'b0};
                writeAddr1 = {writeAddr[11:0], 2'b0};
                writeAddr0 = {writeAddr[8:0], 5'b0};

                readAddr40 = {writeAddr[13:0]};
                readAddr39 = {writeAddr[13:0]};
                readAddr38 = {writeAddr[13:0]};
                readAddr37 = {writeAddr[13:0]};
                readAddr36 = {writeAddr[13:0]};
                readAddr35 = {writeAddr[13:0]};
                readAddr34 = {writeAddr[13:0]};
                readAddr33 = {writeAddr[13:0]};
                readAddr32 = {writeAddr[13:0]};
                readAddr31 = {writeAddr[13:0]};
                readAddr30 = {writeAddr[13:0]};
                readAddr29 = {writeAddr[13:0]};
                readAddr28 = {writeAddr[13:0]};
                readAddr27 = {writeAddr[13:0]};
                readAddr26 = {writeAddr[13:0]};
                readAddr25 = {writeAddr[13:0]};
                readAddr24 = {writeAddr[13:0]};
                readAddr23 = {writeAddr[13:0]};
                readAddr22 = {writeAddr[13:0]};
                readAddr21 = {writeAddr[13:0]};
                readAddr20 = {writeAddr[13:0]};
                readAddr19 = {writeAddr[13:0]};
                readAddr18 = {writeAddr[13:0]};
                readAddr17 = {writeAddr[13:0]};
                readAddr16 = {writeAddr[13:0]};
                readAddr15 = {writeAddr[13:0]};
                readAddr14 = {writeAddr[13:0]};
                readAddr13 = {writeAddr[13:0]};
                readAddr12 = {writeAddr[13:0]};
                readAddr11 = {writeAddr[13:0]};
                readAddr10 = {writeAddr[13:0]};
                readAddr9 = {writeAddr[13:0]};
                readAddr8  = {readAddr[11:0],  2'b0};
                readAddr7  = {readAddr[11:0],  2'b0};
                readAddr6  = {readAddr[11:0],  2'b0};
                readAddr5  = {readAddr[11:0],  2'b0};
                readAddr4  = {readAddr[11:0],  2'b0};
                readAddr3  = {readAddr[11:0],  2'b0};
                readAddr2  = {readAddr[11:0],  2'b0};
                readAddr1  = {readAddr[11:0],  2'b0};
                readAddr0  = {readAddr[8:0],  5'b0};

                writeData40 = {17'b0, writeData[31]};
                writeData39 = {17'b0, writeData[30]};
                writeData38 = {17'b0, writeData[29]};
                writeData37 = {17'b0, writeData[28]};
                writeData36 = {17'b0, writeData[27]};
                writeData35 = {17'b0, writeData[26]};
                writeData34 = {17'b0, writeData[25]};
                writeData33 = {17'b0, writeData[24]};
                writeData32 = {17'b0, writeData[23]};
                writeData31 = {17'b0, writeData[22]};
                writeData30 = {17'b0, writeData[21]};
                writeData29 = {17'b0, writeData[20]};
                writeData28 = {17'b0, writeData[19]};
                writeData27 = {17'b0, writeData[18]};
                writeData26 = {17'b0, writeData[17]};
                writeData25 = {17'b0, writeData[16]};
                writeData24 = {17'b0, writeData[15]};
                writeData23 = {17'b0, writeData[14]};
                writeData22 = {17'b0, writeData[13]};
                writeData21 = {17'b0, writeData[12]};
                writeData20 = {17'b0, writeData[11]};
                writeData19 = {17'b0, writeData[10]};
                writeData18 = {17'b0, writeData[9]};
                writeData17 = {17'b0, writeData[8]};
                writeData16 = {17'b0, writeData[7]};
                writeData15 = {17'b0, writeData[6]};
                writeData14 = {17'b0, writeData[5]};
                writeData13 = {17'b0, writeData[4]};
                writeData12 = {17'b0, writeData[3]};
                writeData11 = {17'b0, writeData[2]};
                writeData10 = {17'b0, writeData[1]};
                writeData9 = {17'b0, writeData[0]};
                writeData8 = {14'b0, writeData[31:28]};
                writeData7 = {14'b0, writeData[27:24]};
                writeData6 = {14'b0, writeData[23:20]};
                writeData5 = {14'b0, writeData[19:16]};
                writeData4 = {14'b0, writeData[15:12]};
                writeData3 = {14'b0, writeData[11:8]};
                writeData2 = {14'b0, writeData[7:4]};
                writeData1 = {14'b0, writeData[3:0]};
                writeData0 = {1'b0, writeData[31:24], 1'b0, writeData[23:16], 1'b0, writeData[15:8], 1'b0, writeData[7:0]};

                case (writeAddr[14:9])
                    6'b000000, 6'b000001, 6'b000010, 6'b000011,
                    6'b000100, 6'b000101, 6'b000110, 6'b000111,
                    6'b001000, 6'b001001, 6'b001010, 6'b001011,
                    6'b001100, 6'b001101, 6'b001110, 6'b001111,
                    6'b010000, 6'b010001, 6'b010010, 6'b010011,
                    6'b010100, 6'b010101, 6'b010110, 6'b010111,
                    6'b011000, 6'b011001, 6'b011010, 6'b011011,
                    6'b011100, 6'b011101, 6'b011110, 6'b011111 : begin
                        wen_a40 = {1'b0, wen};
                        wen_a39 = {1'b0, wen};
                        wen_a38 = {1'b0, wen};
                        wen_a37 = {1'b0, wen};
                        wen_a36 = {1'b0, wen};
                        wen_a35 = {1'b0, wen};
                        wen_a34 = {1'b0, wen};
                        wen_a33 = {1'b0, wen};
                        wen_a32 = {1'b0, wen};
                        wen_a31 = {1'b0, wen};
                        wen_a30 = {1'b0, wen};
                        wen_a29 = {1'b0, wen};
                        wen_a28 = {1'b0, wen};
                        wen_a27 = {1'b0, wen};
                        wen_a26 = {1'b0, wen};
                        wen_a25 = {1'b0, wen};
                        wen_a24 = {1'b0, wen};
                        wen_a23 = {1'b0, wen};
                        wen_a22 = {1'b0, wen};
                        wen_a21 = {1'b0, wen};
                        wen_a20 = {1'b0, wen};
                        wen_a19 = {1'b0, wen};
                        wen_a18 = {1'b0, wen};
                        wen_a17 = {1'b0, wen};
                        wen_a16 = {1'b0, wen};
                        wen_a15 = {1'b0, wen};
                        wen_a14 = {1'b0, wen};
                        wen_a13 = {1'b0, wen};
                        wen_a12 = {1'b0, wen};
                        wen_a11 = {1'b0, wen};
                        wen_a10 = {1'b0, wen};
                        wen_a9 = {1'b0, wen};
                        wen_a8 = {1'b0, 1'b0};
                        wen_a7 = {1'b0, 1'b0};
                        wen_a6 = {1'b0, 1'b0};
                        wen_a5 = {1'b0, 1'b0};
                        wen_a4 = {1'b0, 1'b0};
                        wen_a3 = {1'b0, 1'b0};
                        wen_a2 = {1'b0, 1'b0};
                        wen_a1 = {1'b0, 1'b0};
                        wen_a0 = {1'b0, 1'b0};
                        wen_b0 = {1'b0, 1'b0};
                    end
                    6'b100000, 6'b100001, 6'b100010, 6'b100011,
                    6'b100100, 6'b100101, 6'b100110, 6'b100111: begin
                        wen_a40 = {1'b0, 1'b0};
                        wen_a39 = {1'b0, 1'b0};
                        wen_a38 = {1'b0, 1'b0};
                        wen_a37 = {1'b0, 1'b0};
                        wen_a36 = {1'b0, 1'b0};
                        wen_a35 = {1'b0, 1'b0};
                        wen_a34 = {1'b0, 1'b0};
                        wen_a33 = {1'b0, 1'b0};
                        wen_a32 = {1'b0, 1'b0};
                        wen_a31 = {1'b0, 1'b0};
                        wen_a30 = {1'b0, 1'b0};
                        wen_a29 = {1'b0, 1'b0};
                        wen_a28 = {1'b0, 1'b0};
                        wen_a27 = {1'b0, 1'b0};
                        wen_a26 = {1'b0, 1'b0};
                        wen_a25 = {1'b0, 1'b0};
                        wen_a24 = {1'b0, 1'b0};
                        wen_a23 = {1'b0, 1'b0};
                        wen_a22 = {1'b0, 1'b0};
                        wen_a21 = {1'b0, 1'b0};
                        wen_a20 = {1'b0, 1'b0};
                        wen_a19 = {1'b0, 1'b0};
                        wen_a18 = {1'b0, 1'b0};
                        wen_a17 = {1'b0, 1'b0};
                        wen_a16 = {1'b0, 1'b0};
                        wen_a15 = {1'b0, 1'b0};
                        wen_a14 = {1'b0, 1'b0};
                        wen_a13 = {1'b0, 1'b0};
                        wen_a12 = {1'b0, 1'b0};
                        wen_a11 = {1'b0, 1'b0};
                        wen_a10 = {1'b0, 1'b0};
                        wen_a9 = {1'b0, 1'b0};
                        wen_a8 = {1'b0, wen};
                        wen_a7 = {1'b0, wen};
                        wen_a6 = {1'b0, wen};
                        wen_a5 = {1'b0, wen};
                        wen_a4 = {1'b0, wen};
                        wen_a3 = {1'b0, wen};
                        wen_a2 = {1'b0, wen};
                        wen_a1 = {1'b0, wen};
                        wen_a0 = {1'b0, 1'b0};
                        wen_b0 = {1'b0, 1'b0};
                    end
                    6'b101000: begin
                        wen_a40 = {1'b0, 1'b0};
                        wen_a39 = {1'b0, 1'b0};
                        wen_a38 = {1'b0, 1'b0};
                        wen_a37 = {1'b0, 1'b0};
                        wen_a36 = {1'b0, 1'b0};
                        wen_a35 = {1'b0, 1'b0};
                        wen_a34 = {1'b0, 1'b0};
                        wen_a33 = {1'b0, 1'b0};
                        wen_a32 = {1'b0, 1'b0};
                        wen_a31 = {1'b0, 1'b0};
                        wen_a30 = {1'b0, 1'b0};
                        wen_a29 = {1'b0, 1'b0};
                        wen_a28 = {1'b0, 1'b0};
                        wen_a27 = {1'b0, 1'b0};
                        wen_a26 = {1'b0, 1'b0};
                        wen_a25 = {1'b0, 1'b0};
                        wen_a24 = {1'b0, 1'b0};
                        wen_a23 = {1'b0, 1'b0};
                        wen_a22 = {1'b0, 1'b0};
                        wen_a21 = {1'b0, 1'b0};
                        wen_a20 = {1'b0, 1'b0};
                        wen_a19 = {1'b0, 1'b0};
                        wen_a18 = {1'b0, 1'b0};
                        wen_a17 = {1'b0, 1'b0};
                        wen_a16 = {1'b0, 1'b0};
                        wen_a15 = {1'b0, 1'b0};
                        wen_a14 = {1'b0, 1'b0};
                        wen_a13 = {1'b0, 1'b0};
                        wen_a12 = {1'b0, 1'b0};
                        wen_a11 = {1'b0, 1'b0};
                        wen_a10 = {1'b0, 1'b0};
                        wen_a9 = {1'b0, 1'b0};
                        wen_a8 = {1'b0, 1'b0};
                        wen_a7 = {1'b0, 1'b0};
                        wen_a6 = {1'b0, 1'b0};
                        wen_a5 = {1'b0, 1'b0};
                        wen_a4 = {1'b0, 1'b0};
                        wen_a3 = {1'b0, 1'b0};
                        wen_a2 = {1'b0, 1'b0};
                        wen_a1 = {1'b0, 1'b0};
                        wen_a0 = {wen, wen};
                        wen_b0 = {wen, wen};
                    end
                    default : begin
                        wen_a40 = {1'b0, 1'b0};
                        wen_a39 = {1'b0, 1'b0};
                        wen_a38 = {1'b0, 1'b0};
                        wen_a37 = {1'b0, 1'b0};
                        wen_a36 = {1'b0, 1'b0};
                        wen_a35 = {1'b0, 1'b0};
                        wen_a34 = {1'b0, 1'b0};
                        wen_a33 = {1'b0, 1'b0};
                        wen_a32 = {1'b0, 1'b0};
                        wen_a31 = {1'b0, 1'b0};
                        wen_a30 = {1'b0, 1'b0};
                        wen_a29 = {1'b0, 1'b0};
                        wen_a28 = {1'b0, 1'b0};
                        wen_a27 = {1'b0, 1'b0};
                        wen_a26 = {1'b0, 1'b0};
                        wen_a25 = {1'b0, 1'b0};
                        wen_a24 = {1'b0, 1'b0};
                        wen_a23 = {1'b0, 1'b0};
                        wen_a22 = {1'b0, 1'b0};
                        wen_a21 = {1'b0, 1'b0};
                        wen_a20 = {1'b0, 1'b0};
                        wen_a19 = {1'b0, 1'b0};
                        wen_a18 = {1'b0, 1'b0};
                        wen_a17 = {1'b0, 1'b0};
                        wen_a16 = {1'b0, 1'b0};
                        wen_a15 = {1'b0, 1'b0};
                        wen_a14 = {1'b0, 1'b0};
                        wen_a13 = {1'b0, 1'b0};
                        wen_a12 = {1'b0, 1'b0};
                        wen_a11 = {1'b0, 1'b0};
                        wen_a10 = {1'b0, 1'b0};
                        wen_a9 = {1'b0, 1'b0};
                        wen_a8 = {1'b0, 1'b0};
                        wen_a7 = {1'b0, 1'b0};
                        wen_a6 = {1'b0, 1'b0};
                        wen_a5 = {1'b0, 1'b0};
                        wen_a4 = {1'b0, 1'b0};
                        wen_a3 = {1'b0, 1'b0};
                        wen_a2 = {1'b0, 1'b0};
                        wen_a1 = {1'b0, 1'b0};
                        wen_a0 = {1'b0, 1'b0};
                        wen_b0 = {1'b0, 1'b0};
                    end
                endcase

                case (ckRdAddr[14:9])
                    6'b000000, 6'b000001, 6'b000010, 6'b000011,
                    6'b000100, 6'b000101, 6'b000110, 6'b000111,
                    6'b001000, 6'b001001, 6'b001010, 6'b001011,
                    6'b001100, 6'b001101, 6'b001110, 6'b001111,
                    6'b010000, 6'b010001, 6'b010010, 6'b010011,
                    6'b010100, 6'b010101, 6'b010110, 6'b010111,
                    6'b011000, 6'b011001, 6'b011010, 6'b011011,
                    6'b011100, 6'b011101, 6'b011110, 6'b011111 : begin
                        readData = {
                                        readData40[0],
                                        readData39[0],
                                        readData38[0],
                                        readData37[0],
                                        readData36[0],
                                        readData35[0],
                                        readData34[0],
                                        readData33[0],
                                        readData32[0],
                                        readData31[0],
                                        readData30[0],
                                        readData29[0],
                                        readData28[0],
                                        readData27[0],
                                        readData26[0],
                                        readData25[0],
                                        readData24[0],
                                        readData23[0],
                                        readData22[0],
                                        readData21[0],
                                        readData20[0],
                                        readData19[0],
                                        readData18[0],
                                        readData17[0],
                                        readData16[0],
                                        readData15[0],
                                        readData14[0],
                                        readData13[0],
                                        readData12[0],
                                        readData11[0],
                                        readData10[0],
                                        readData9[0]
                        };
                    end
                    6'b100000, 6'b100001, 6'b100010, 6'b100011,
                    6'b100100, 6'b100101, 6'b100110, 6'b100111: begin
                        readData = {
                                        readData8[3:0],
                                        readData7[3:0],
                                        readData6[3:0],
                                        readData5[3:0],
                                        readData4[3:0],
                                        readData3[3:0],
                                        readData2[3:0],
                                        readData1[3:0]
                        };
                    end
                    6'b101000: begin
                        readData = {readData0[34:27],readData0[25:18],readData0[16:9],readData0[7:0]};
                    end
                    default : begin
                        readData = 32'b0;
                    end
                endcase
            end
            21504: begin
                width42 = 3'b000;
                width41 = 3'b000;
                width40 = 3'b000;
                width39 = 3'b000;
                width38 = 3'b000;
                width37 = 3'b000;
                width36 = 3'b000;
                width35 = 3'b000;
                width34 = 3'b000;
                width33 = 3'b000;
                width32 = 3'b000;
                width31 = 3'b000;
                width30 = 3'b000;
                width29 = 3'b000;
                width28 = 3'b000;
                width27 = 3'b000;
                width26 = 3'b000;
                width25 = 3'b000;
                width24 = 3'b000;
                width23 = 3'b000;
                width22 = 3'b000;
                width21 = 3'b000;
                width20 = 3'b000;
                width19 = 3'b000;
                width18 = 3'b000;
                width17 = 3'b000;
                width16 = 3'b000;
                width15 = 3'b000;
                width14 = 3'b000;
                width13 = 3'b000;
                width12 = 3'b000;
                width11 = 3'b000;
                width10 = 3'b010;
                width9 = 3'b010;
                width8 = 3'b010;
                width7 = 3'b010;
                width6 = 3'b010;
                width5 = 3'b010;
                width4 = 3'b010;
                width3 = 3'b010;
                width2 = 3'b100;
                width1 = 3'b100;

                writeAddr42 = {writeAddr[13:0]};
                writeAddr41 = {writeAddr[13:0]};
                writeAddr40 = {writeAddr[13:0]};
                writeAddr39 = {writeAddr[13:0]};
                writeAddr38 = {writeAddr[13:0]};
                writeAddr37 = {writeAddr[13:0]};
                writeAddr36 = {writeAddr[13:0]};
                writeAddr35 = {writeAddr[13:0]};
                writeAddr34 = {writeAddr[13:0]};
                writeAddr33 = {writeAddr[13:0]};
                writeAddr32 = {writeAddr[13:0]};
                writeAddr31 = {writeAddr[13:0]};
                writeAddr30 = {writeAddr[13:0]};
                writeAddr29 = {writeAddr[13:0]};
                writeAddr28 = {writeAddr[13:0]};
                writeAddr27 = {writeAddr[13:0]};
                writeAddr26 = {writeAddr[13:0]};
                writeAddr25 = {writeAddr[13:0]};
                writeAddr24 = {writeAddr[13:0]};
                writeAddr23 = {writeAddr[13:0]};
                writeAddr22 = {writeAddr[13:0]};
                writeAddr21 = {writeAddr[13:0]};
                writeAddr20 = {writeAddr[13:0]};
                writeAddr19 = {writeAddr[13:0]};
                writeAddr18 = {writeAddr[13:0]};
                writeAddr17 = {writeAddr[13:0]};
                writeAddr16 = {writeAddr[13:0]};
                writeAddr15 = {writeAddr[13:0]};
                writeAddr14 = {writeAddr[13:0]};
                writeAddr13 = {writeAddr[13:0]};
                writeAddr12 = {writeAddr[13:0]};
                writeAddr11 = {writeAddr[13:0]};
                writeAddr10 = {writeAddr[11:0], 2'b0};
                writeAddr9 = {writeAddr[11:0], 2'b0};
                writeAddr8 = {writeAddr[11:0], 2'b0};
                writeAddr7 = {writeAddr[11:0], 2'b0};
                writeAddr6 = {writeAddr[11:0], 2'b0};
                writeAddr5 = {writeAddr[11:0], 2'b0};
                writeAddr4 = {writeAddr[11:0], 2'b0};
                writeAddr3 = {writeAddr[11:0], 2'b0};
                writeAddr2 = {writeAddr[9:0], 4'b0};
                writeAddr1 = {writeAddr[9:0], 4'b0};

                readAddr42 = {writeAddr[13:0]};
                readAddr41 = {writeAddr[13:0]};
                readAddr40 = {writeAddr[13:0]};
                readAddr39 = {writeAddr[13:0]};
                readAddr38 = {writeAddr[13:0]};
                readAddr37 = {writeAddr[13:0]};
                readAddr36 = {writeAddr[13:0]};
                readAddr35 = {writeAddr[13:0]};
                readAddr34 = {writeAddr[13:0]};
                readAddr33 = {writeAddr[13:0]};
                readAddr32 = {writeAddr[13:0]};
                readAddr31 = {writeAddr[13:0]};
                readAddr30 = {writeAddr[13:0]};
                readAddr29 = {writeAddr[13:0]};
                readAddr28 = {writeAddr[13:0]};
                readAddr27 = {writeAddr[13:0]};
                readAddr26 = {writeAddr[13:0]};
                readAddr25 = {writeAddr[13:0]};
                readAddr24 = {writeAddr[13:0]};
                readAddr23 = {writeAddr[13:0]};
                readAddr22 = {writeAddr[13:0]};
                readAddr21 = {writeAddr[13:0]};
                readAddr20 = {writeAddr[13:0]};
                readAddr19 = {writeAddr[13:0]};
                readAddr18 = {writeAddr[13:0]};
                readAddr17 = {writeAddr[13:0]};
                readAddr16 = {writeAddr[13:0]};
                readAddr15 = {writeAddr[13:0]};
                readAddr14 = {writeAddr[13:0]};
                readAddr13 = {writeAddr[13:0]};
                readAddr12 = {writeAddr[13:0]};
                readAddr11 = {writeAddr[13:0]};
                readAddr10  = {readAddr[11:0],  2'b0};
                readAddr9  = {readAddr[11:0],  2'b0};
                readAddr8  = {readAddr[11:0],  2'b0};
                readAddr7  = {readAddr[11:0],  2'b0};
                readAddr6  = {readAddr[11:0],  2'b0};
                readAddr5  = {readAddr[11:0],  2'b0};
                readAddr4  = {readAddr[11:0],  2'b0};
                readAddr3  = {readAddr[11:0],  2'b0};
                readAddr2  = {readAddr[9:0],  4'b0};
                readAddr1  = {readAddr[9:0],  4'b0};

                writeData42 = {17'b0, writeData[31]};
                writeData41 = {17'b0, writeData[30]};
                writeData40 = {17'b0, writeData[29]};
                writeData39 = {17'b0, writeData[28]};
                writeData38 = {17'b0, writeData[27]};
                writeData37 = {17'b0, writeData[26]};
                writeData36 = {17'b0, writeData[25]};
                writeData35 = {17'b0, writeData[24]};
                writeData34 = {17'b0, writeData[23]};
                writeData33 = {17'b0, writeData[22]};
                writeData32 = {17'b0, writeData[21]};
                writeData31 = {17'b0, writeData[20]};
                writeData30 = {17'b0, writeData[19]};
                writeData29 = {17'b0, writeData[18]};
                writeData28 = {17'b0, writeData[17]};
                writeData27 = {17'b0, writeData[16]};
                writeData26 = {17'b0, writeData[15]};
                writeData25 = {17'b0, writeData[14]};
                writeData24 = {17'b0, writeData[13]};
                writeData23 = {17'b0, writeData[12]};
                writeData22 = {17'b0, writeData[11]};
                writeData21 = {17'b0, writeData[10]};
                writeData20 = {17'b0, writeData[9]};
                writeData19 = {17'b0, writeData[8]};
                writeData18 = {17'b0, writeData[7]};
                writeData17 = {17'b0, writeData[6]};
                writeData16 = {17'b0, writeData[5]};
                writeData15 = {17'b0, writeData[4]};
                writeData14 = {17'b0, writeData[3]};
                writeData13 = {17'b0, writeData[2]};
                writeData12 = {17'b0, writeData[1]};
                writeData11 = {17'b0, writeData[0]};
                writeData10 = {14'b0, writeData[31:28]};
                writeData9 = {14'b0, writeData[27:24]};
                writeData8 = {14'b0, writeData[23:20]};
                writeData7 = {14'b0, writeData[19:16]};
                writeData6 = {14'b0, writeData[15:12]};
                writeData5 = {14'b0, writeData[11:8]};
                writeData4 = {14'b0, writeData[7:4]};
                writeData3 = {14'b0, writeData[3:0]};
                writeData2 = {1'b0, writeData[31:24], 1'b0, writeData[23:16]};
                writeData1 = {1'b0, writeData[15:8], 1'b0, writeData[7:0]};

                case (writeAddr[14:9])
                    6'b000000, 6'b000001, 6'b000010, 6'b000011,
                    6'b000100, 6'b000101, 6'b000110, 6'b000111,
                    6'b001000, 6'b001001, 6'b001010, 6'b001011,
                    6'b001100, 6'b001101, 6'b001110, 6'b001111,
                    6'b010000, 6'b010001, 6'b010010, 6'b010011,
                    6'b010100, 6'b010101, 6'b010110, 6'b010111,
                    6'b011000, 6'b011001, 6'b011010, 6'b011011,
                    6'b011100, 6'b011101, 6'b011110, 6'b011111 : begin
                        wen_a42 = {1'b0, wen};
                        wen_a41 = {1'b0, wen};
                        wen_a40 = {1'b0, wen};
                        wen_a39 = {1'b0, wen};
                        wen_a38 = {1'b0, wen};
                        wen_a37 = {1'b0, wen};
                        wen_a36 = {1'b0, wen};
                        wen_a35 = {1'b0, wen};
                        wen_a34 = {1'b0, wen};
                        wen_a33 = {1'b0, wen};
                        wen_a32 = {1'b0, wen};
                        wen_a31 = {1'b0, wen};
                        wen_a30 = {1'b0, wen};
                        wen_a29 = {1'b0, wen};
                        wen_a28 = {1'b0, wen};
                        wen_a27 = {1'b0, wen};
                        wen_a26 = {1'b0, wen};
                        wen_a25 = {1'b0, wen};
                        wen_a24 = {1'b0, wen};
                        wen_a23 = {1'b0, wen};
                        wen_a22 = {1'b0, wen};
                        wen_a21 = {1'b0, wen};
                        wen_a20 = {1'b0, wen};
                        wen_a19 = {1'b0, wen};
                        wen_a18 = {1'b0, wen};
                        wen_a17 = {1'b0, wen};
                        wen_a16 = {1'b0, wen};
                        wen_a15 = {1'b0, wen};
                        wen_a14 = {1'b0, wen};
                        wen_a13 = {1'b0, wen};
                        wen_a12 = {1'b0, wen};
                        wen_a11 = {1'b0, wen};
                        wen_a10 = {1'b0, 1'b0};
                        wen_a9 = {1'b0, 1'b0};
                        wen_a8 = {1'b0, 1'b0};
                        wen_a7 = {1'b0, 1'b0};
                        wen_a6 = {1'b0, 1'b0};
                        wen_a5 = {1'b0, 1'b0};
                        wen_a4 = {1'b0, 1'b0};
                        wen_a3 = {1'b0, 1'b0};
                        wen_a2 = {1'b0, 1'b0};
                        wen_a1 = {1'b0, 1'b0};
                    end
                    6'b100000, 6'b100001, 6'b100010, 6'b100011,
                    6'b100100, 6'b100101, 6'b100110, 6'b100111: begin
                        wen_a42 = {1'b0, 1'b0};
                        wen_a41 = {1'b0, 1'b0};
                        wen_a40 = {1'b0, 1'b0};
                        wen_a39 = {1'b0, 1'b0};
                        wen_a38 = {1'b0, 1'b0};
                        wen_a37 = {1'b0, 1'b0};
                        wen_a36 = {1'b0, 1'b0};
                        wen_a35 = {1'b0, 1'b0};
                        wen_a34 = {1'b0, 1'b0};
                        wen_a33 = {1'b0, 1'b0};
                        wen_a32 = {1'b0, 1'b0};
                        wen_a31 = {1'b0, 1'b0};
                        wen_a30 = {1'b0, 1'b0};
                        wen_a29 = {1'b0, 1'b0};
                        wen_a28 = {1'b0, 1'b0};
                        wen_a27 = {1'b0, 1'b0};
                        wen_a26 = {1'b0, 1'b0};
                        wen_a25 = {1'b0, 1'b0};
                        wen_a24 = {1'b0, 1'b0};
                        wen_a23 = {1'b0, 1'b0};
                        wen_a22 = {1'b0, 1'b0};
                        wen_a21 = {1'b0, 1'b0};
                        wen_a20 = {1'b0, 1'b0};
                        wen_a19 = {1'b0, 1'b0};
                        wen_a18 = {1'b0, 1'b0};
                        wen_a17 = {1'b0, 1'b0};
                        wen_a16 = {1'b0, 1'b0};
                        wen_a15 = {1'b0, 1'b0};
                        wen_a14 = {1'b0, 1'b0};
                        wen_a13 = {1'b0, 1'b0};
                        wen_a12 = {1'b0, 1'b0};
                        wen_a11 = {1'b0, 1'b0};
                        wen_a10 = {1'b0, wen};
                        wen_a9 = {1'b0, wen};
                        wen_a8 = {1'b0, wen};
                        wen_a7 = {1'b0, wen};
                        wen_a6 = {1'b0, wen};
                        wen_a5 = {1'b0, wen};
                        wen_a4 = {1'b0, wen};
                        wen_a3 = {1'b0, wen};
                        wen_a2 = {1'b0, 1'b0};
                        wen_a1 = {1'b0, 1'b0};
                    end
                    6'b101000, 6'b101001 : begin
                        wen_a42 = {1'b0, 1'b0};
                        wen_a41 = {1'b0, 1'b0};
                        wen_a40 = {1'b0, 1'b0};
                        wen_a39 = {1'b0, 1'b0};
                        wen_a38 = {1'b0, 1'b0};
                        wen_a37 = {1'b0, 1'b0};
                        wen_a36 = {1'b0, 1'b0};
                        wen_a35 = {1'b0, 1'b0};
                        wen_a34 = {1'b0, 1'b0};
                        wen_a33 = {1'b0, 1'b0};
                        wen_a32 = {1'b0, 1'b0};
                        wen_a31 = {1'b0, 1'b0};
                        wen_a30 = {1'b0, 1'b0};
                        wen_a29 = {1'b0, 1'b0};
                        wen_a28 = {1'b0, 1'b0};
                        wen_a27 = {1'b0, 1'b0};
                        wen_a26 = {1'b0, 1'b0};
                        wen_a25 = {1'b0, 1'b0};
                        wen_a24 = {1'b0, 1'b0};
                        wen_a23 = {1'b0, 1'b0};
                        wen_a22 = {1'b0, 1'b0};
                        wen_a21 = {1'b0, 1'b0};
                        wen_a20 = {1'b0, 1'b0};
                        wen_a19 = {1'b0, 1'b0};
                        wen_a18 = {1'b0, 1'b0};
                        wen_a17 = {1'b0, 1'b0};
                        wen_a16 = {1'b0, 1'b0};
                        wen_a15 = {1'b0, 1'b0};
                        wen_a14 = {1'b0, 1'b0};
                        wen_a13 = {1'b0, 1'b0};
                        wen_a12 = {1'b0, 1'b0};
                        wen_a11 = {1'b0, 1'b0};
                        wen_a10 = {1'b0, 1'b0};
                        wen_a9 = {1'b0, 1'b0};
                        wen_a8 = {1'b0, 1'b0};
                        wen_a7 = {1'b0, 1'b0};
                        wen_a6 = {1'b0, 1'b0};
                        wen_a5 = {1'b0, 1'b0};
                        wen_a4 = {1'b0, 1'b0};
                        wen_a3 = {1'b0, 1'b0};
                        wen_a2 = {wen, wen};
                        wen_a1 = {wen, wen};
                    end
                    default : begin
                        wen_a42 = {1'b0, 1'b0};
                        wen_a41 = {1'b0, 1'b0};
                        wen_a40 = {1'b0, 1'b0};
                        wen_a39 = {1'b0, 1'b0};
                        wen_a38 = {1'b0, 1'b0};
                        wen_a37 = {1'b0, 1'b0};
                        wen_a36 = {1'b0, 1'b0};
                        wen_a35 = {1'b0, 1'b0};
                        wen_a34 = {1'b0, 1'b0};
                        wen_a33 = {1'b0, 1'b0};
                        wen_a32 = {1'b0, 1'b0};
                        wen_a31 = {1'b0, 1'b0};
                        wen_a30 = {1'b0, 1'b0};
                        wen_a29 = {1'b0, 1'b0};
                        wen_a28 = {1'b0, 1'b0};
                        wen_a27 = {1'b0, 1'b0};
                        wen_a26 = {1'b0, 1'b0};
                        wen_a25 = {1'b0, 1'b0};
                        wen_a24 = {1'b0, 1'b0};
                        wen_a23 = {1'b0, 1'b0};
                        wen_a22 = {1'b0, 1'b0};
                        wen_a21 = {1'b0, 1'b0};
                        wen_a20 = {1'b0, 1'b0};
                        wen_a19 = {1'b0, 1'b0};
                        wen_a18 = {1'b0, 1'b0};
                        wen_a17 = {1'b0, 1'b0};
                        wen_a16 = {1'b0, 1'b0};
                        wen_a15 = {1'b0, 1'b0};
                        wen_a14 = {1'b0, 1'b0};
                        wen_a13 = {1'b0, 1'b0};
                        wen_a12 = {1'b0, 1'b0};
                        wen_a11 = {1'b0, 1'b0};
                        wen_a10 = {1'b0, 1'b0};
                        wen_a9 = {1'b0, 1'b0};
                        wen_a8 = {1'b0, 1'b0};
                        wen_a7 = {1'b0, 1'b0};
                        wen_a6 = {1'b0, 1'b0};
                        wen_a5 = {1'b0, 1'b0};
                        wen_a4 = {1'b0, 1'b0};
                        wen_a3 = {1'b0, 1'b0};
                        wen_a2 = {1'b0, 1'b0};
                        wen_a1 = {1'b0, 1'b0};
                    end
                endcase

                case (ckRdAddr[14:9])
                    6'b000000, 6'b000001, 6'b000010, 6'b000011,
                    6'b000100, 6'b000101, 6'b000110, 6'b000111,
                    6'b001000, 6'b001001, 6'b001010, 6'b001011,
                    6'b001100, 6'b001101, 6'b001110, 6'b001111,
                    6'b010000, 6'b010001, 6'b010010, 6'b010011,
                    6'b010100, 6'b010101, 6'b010110, 6'b010111,
                    6'b011000, 6'b011001, 6'b011010, 6'b011011,
                    6'b011100, 6'b011101, 6'b011110, 6'b011111 : begin
                        readData = {
                                        readData42[0],
                                        readData41[0],
                                        readData40[0],
                                        readData39[0],
                                        readData38[0],
                                        readData37[0],
                                        readData36[0],
                                        readData35[0],
                                        readData34[0],
                                        readData33[0],
                                        readData32[0],
                                        readData31[0],
                                        readData30[0],
                                        readData29[0],
                                        readData28[0],
                                        readData27[0],
                                        readData26[0],
                                        readData25[0],
                                        readData24[0],
                                        readData23[0],
                                        readData22[0],
                                        readData21[0],
                                        readData20[0],
                                        readData19[0],
                                        readData18[0],
                                        readData17[0],
                                        readData16[0],
                                        readData15[0],
                                        readData14[0],
                                        readData13[0],
                                        readData12[0],
                                        readData11[0]
                        };
                    end
                    6'b100000, 6'b100001, 6'b100010, 6'b100011,
                    6'b100100, 6'b100101, 6'b100110, 6'b100111: begin
                        readData = {
                                        readData10[3:0],
                                        readData9[3:0],
                                        readData8[3:0],
                                        readData7[3:0],
                                        readData6[3:0],
                                        readData5[3:0],
                                        readData4[3:0],
                                        readData3[3:0]
                        };
                    end
                    6'b101000, 6'b101001 : begin
                        readData = {readData2[16:9],readData2[7:0],readData1[16:9],readData1[7:0]};
                    end
                    default : begin
                        readData = 32'b0;
                    end
                endcase
            end
            22016: begin
                width42 = 3'b000;
                width41 = 3'b000;
                width40 = 3'b000;
                width39 = 3'b000;
                width38 = 3'b000;
                width37 = 3'b000;
                width36 = 3'b000;
                width35 = 3'b000;
                width34 = 3'b000;
                width33 = 3'b000;
                width32 = 3'b000;
                width31 = 3'b000;
                width30 = 3'b000;
                width29 = 3'b000;
                width28 = 3'b000;
                width27 = 3'b000;
                width26 = 3'b000;
                width25 = 3'b000;
                width24 = 3'b000;
                width23 = 3'b000;
                width22 = 3'b000;
                width21 = 3'b000;
                width20 = 3'b000;
                width19 = 3'b000;
                width18 = 3'b000;
                width17 = 3'b000;
                width16 = 3'b000;
                width15 = 3'b000;
                width14 = 3'b000;
                width13 = 3'b000;
                width12 = 3'b000;
                width11 = 3'b000;
                width10 = 3'b010;
                width9 = 3'b010;
                width8 = 3'b010;
                width7 = 3'b010;
                width6 = 3'b010;
                width5 = 3'b010;
                width4 = 3'b010;
                width3 = 3'b010;
                width2 = 3'b100;
                width1 = 3'b100;
                width0 = 3'b101;

                writeAddr42 = {writeAddr[13:0]};
                writeAddr41 = {writeAddr[13:0]};
                writeAddr40 = {writeAddr[13:0]};
                writeAddr39 = {writeAddr[13:0]};
                writeAddr38 = {writeAddr[13:0]};
                writeAddr37 = {writeAddr[13:0]};
                writeAddr36 = {writeAddr[13:0]};
                writeAddr35 = {writeAddr[13:0]};
                writeAddr34 = {writeAddr[13:0]};
                writeAddr33 = {writeAddr[13:0]};
                writeAddr32 = {writeAddr[13:0]};
                writeAddr31 = {writeAddr[13:0]};
                writeAddr30 = {writeAddr[13:0]};
                writeAddr29 = {writeAddr[13:0]};
                writeAddr28 = {writeAddr[13:0]};
                writeAddr27 = {writeAddr[13:0]};
                writeAddr26 = {writeAddr[13:0]};
                writeAddr25 = {writeAddr[13:0]};
                writeAddr24 = {writeAddr[13:0]};
                writeAddr23 = {writeAddr[13:0]};
                writeAddr22 = {writeAddr[13:0]};
                writeAddr21 = {writeAddr[13:0]};
                writeAddr20 = {writeAddr[13:0]};
                writeAddr19 = {writeAddr[13:0]};
                writeAddr18 = {writeAddr[13:0]};
                writeAddr17 = {writeAddr[13:0]};
                writeAddr16 = {writeAddr[13:0]};
                writeAddr15 = {writeAddr[13:0]};
                writeAddr14 = {writeAddr[13:0]};
                writeAddr13 = {writeAddr[13:0]};
                writeAddr12 = {writeAddr[13:0]};
                writeAddr11 = {writeAddr[13:0]};
                writeAddr10 = {writeAddr[11:0], 2'b0};
                writeAddr9 = {writeAddr[11:0], 2'b0};
                writeAddr8 = {writeAddr[11:0], 2'b0};
                writeAddr7 = {writeAddr[11:0], 2'b0};
                writeAddr6 = {writeAddr[11:0], 2'b0};
                writeAddr5 = {writeAddr[11:0], 2'b0};
                writeAddr4 = {writeAddr[11:0], 2'b0};
                writeAddr3 = {writeAddr[11:0], 2'b0};
                writeAddr2 = {writeAddr[9:0], 4'b0};
                writeAddr1 = {writeAddr[9:0], 4'b0};
                writeAddr0 = {writeAddr[8:0], 5'b0};

                readAddr42 = {writeAddr[13:0]};
                readAddr41 = {writeAddr[13:0]};
                readAddr40 = {writeAddr[13:0]};
                readAddr39 = {writeAddr[13:0]};
                readAddr38 = {writeAddr[13:0]};
                readAddr37 = {writeAddr[13:0]};
                readAddr36 = {writeAddr[13:0]};
                readAddr35 = {writeAddr[13:0]};
                readAddr34 = {writeAddr[13:0]};
                readAddr33 = {writeAddr[13:0]};
                readAddr32 = {writeAddr[13:0]};
                readAddr31 = {writeAddr[13:0]};
                readAddr30 = {writeAddr[13:0]};
                readAddr29 = {writeAddr[13:0]};
                readAddr28 = {writeAddr[13:0]};
                readAddr27 = {writeAddr[13:0]};
                readAddr26 = {writeAddr[13:0]};
                readAddr25 = {writeAddr[13:0]};
                readAddr24 = {writeAddr[13:0]};
                readAddr23 = {writeAddr[13:0]};
                readAddr22 = {writeAddr[13:0]};
                readAddr21 = {writeAddr[13:0]};
                readAddr20 = {writeAddr[13:0]};
                readAddr19 = {writeAddr[13:0]};
                readAddr18 = {writeAddr[13:0]};
                readAddr17 = {writeAddr[13:0]};
                readAddr16 = {writeAddr[13:0]};
                readAddr15 = {writeAddr[13:0]};
                readAddr14 = {writeAddr[13:0]};
                readAddr13 = {writeAddr[13:0]};
                readAddr12 = {writeAddr[13:0]};
                readAddr11 = {writeAddr[13:0]};
                readAddr10  = {readAddr[11:0],  2'b0};
                readAddr9  = {readAddr[11:0],  2'b0};
                readAddr8  = {readAddr[11:0],  2'b0};
                readAddr7  = {readAddr[11:0],  2'b0};
                readAddr6  = {readAddr[11:0],  2'b0};
                readAddr5  = {readAddr[11:0],  2'b0};
                readAddr4  = {readAddr[11:0],  2'b0};
                readAddr3  = {readAddr[11:0],  2'b0};
                readAddr2  = {readAddr[9:0],  4'b0};
                readAddr1  = {readAddr[9:0],  4'b0};
                readAddr0  = {readAddr[8:0],  5'b0};

                writeData42 = {17'b0, writeData[31]};
                writeData41 = {17'b0, writeData[30]};
                writeData40 = {17'b0, writeData[29]};
                writeData39 = {17'b0, writeData[28]};
                writeData38 = {17'b0, writeData[27]};
                writeData37 = {17'b0, writeData[26]};
                writeData36 = {17'b0, writeData[25]};
                writeData35 = {17'b0, writeData[24]};
                writeData34 = {17'b0, writeData[23]};
                writeData33 = {17'b0, writeData[22]};
                writeData32 = {17'b0, writeData[21]};
                writeData31 = {17'b0, writeData[20]};
                writeData30 = {17'b0, writeData[19]};
                writeData29 = {17'b0, writeData[18]};
                writeData28 = {17'b0, writeData[17]};
                writeData27 = {17'b0, writeData[16]};
                writeData26 = {17'b0, writeData[15]};
                writeData25 = {17'b0, writeData[14]};
                writeData24 = {17'b0, writeData[13]};
                writeData23 = {17'b0, writeData[12]};
                writeData22 = {17'b0, writeData[11]};
                writeData21 = {17'b0, writeData[10]};
                writeData20 = {17'b0, writeData[9]};
                writeData19 = {17'b0, writeData[8]};
                writeData18 = {17'b0, writeData[7]};
                writeData17 = {17'b0, writeData[6]};
                writeData16 = {17'b0, writeData[5]};
                writeData15 = {17'b0, writeData[4]};
                writeData14 = {17'b0, writeData[3]};
                writeData13 = {17'b0, writeData[2]};
                writeData12 = {17'b0, writeData[1]};
                writeData11 = {17'b0, writeData[0]};
                writeData10 = {14'b0, writeData[31:28]};
                writeData9 = {14'b0, writeData[27:24]};
                writeData8 = {14'b0, writeData[23:20]};
                writeData7 = {14'b0, writeData[19:16]};
                writeData6 = {14'b0, writeData[15:12]};
                writeData5 = {14'b0, writeData[11:8]};
                writeData4 = {14'b0, writeData[7:4]};
                writeData3 = {14'b0, writeData[3:0]};
                writeData2 = {1'b0, writeData[31:24], 1'b0, writeData[23:16]};
                writeData1 = {1'b0, writeData[15:8], 1'b0, writeData[7:0]};
                writeData0 = {1'b0, writeData[31:24], 1'b0, writeData[23:16], 1'b0, writeData[15:8], 1'b0, writeData[7:0]};

                case (writeAddr[14:9])
                    6'b000000, 6'b000001, 6'b000010, 6'b000011,
                    6'b000100, 6'b000101, 6'b000110, 6'b000111,
                    6'b001000, 6'b001001, 6'b001010, 6'b001011,
                    6'b001100, 6'b001101, 6'b001110, 6'b001111,
                    6'b010000, 6'b010001, 6'b010010, 6'b010011,
                    6'b010100, 6'b010101, 6'b010110, 6'b010111,
                    6'b011000, 6'b011001, 6'b011010, 6'b011011,
                    6'b011100, 6'b011101, 6'b011110, 6'b011111 : begin
                        wen_a42 = {1'b0, wen};
                        wen_a41 = {1'b0, wen};
                        wen_a40 = {1'b0, wen};
                        wen_a39 = {1'b0, wen};
                        wen_a38 = {1'b0, wen};
                        wen_a37 = {1'b0, wen};
                        wen_a36 = {1'b0, wen};
                        wen_a35 = {1'b0, wen};
                        wen_a34 = {1'b0, wen};
                        wen_a33 = {1'b0, wen};
                        wen_a32 = {1'b0, wen};
                        wen_a31 = {1'b0, wen};
                        wen_a30 = {1'b0, wen};
                        wen_a29 = {1'b0, wen};
                        wen_a28 = {1'b0, wen};
                        wen_a27 = {1'b0, wen};
                        wen_a26 = {1'b0, wen};
                        wen_a25 = {1'b0, wen};
                        wen_a24 = {1'b0, wen};
                        wen_a23 = {1'b0, wen};
                        wen_a22 = {1'b0, wen};
                        wen_a21 = {1'b0, wen};
                        wen_a20 = {1'b0, wen};
                        wen_a19 = {1'b0, wen};
                        wen_a18 = {1'b0, wen};
                        wen_a17 = {1'b0, wen};
                        wen_a16 = {1'b0, wen};
                        wen_a15 = {1'b0, wen};
                        wen_a14 = {1'b0, wen};
                        wen_a13 = {1'b0, wen};
                        wen_a12 = {1'b0, wen};
                        wen_a11 = {1'b0, wen};
                        wen_a10 = {1'b0, 1'b0};
                        wen_a9 = {1'b0, 1'b0};
                        wen_a8 = {1'b0, 1'b0};
                        wen_a7 = {1'b0, 1'b0};
                        wen_a6 = {1'b0, 1'b0};
                        wen_a5 = {1'b0, 1'b0};
                        wen_a4 = {1'b0, 1'b0};
                        wen_a3 = {1'b0, 1'b0};
                        wen_a2 = {1'b0, 1'b0};
                        wen_a1 = {1'b0, 1'b0};
                        wen_a0 = {1'b0, 1'b0};
                        wen_b0 = {1'b0, 1'b0};
                    end
                    6'b100000, 6'b100001, 6'b100010, 6'b100011,
                    6'b100100, 6'b100101, 6'b100110, 6'b100111: begin
                        wen_a42 = {1'b0, 1'b0};
                        wen_a41 = {1'b0, 1'b0};
                        wen_a40 = {1'b0, 1'b0};
                        wen_a39 = {1'b0, 1'b0};
                        wen_a38 = {1'b0, 1'b0};
                        wen_a37 = {1'b0, 1'b0};
                        wen_a36 = {1'b0, 1'b0};
                        wen_a35 = {1'b0, 1'b0};
                        wen_a34 = {1'b0, 1'b0};
                        wen_a33 = {1'b0, 1'b0};
                        wen_a32 = {1'b0, 1'b0};
                        wen_a31 = {1'b0, 1'b0};
                        wen_a30 = {1'b0, 1'b0};
                        wen_a29 = {1'b0, 1'b0};
                        wen_a28 = {1'b0, 1'b0};
                        wen_a27 = {1'b0, 1'b0};
                        wen_a26 = {1'b0, 1'b0};
                        wen_a25 = {1'b0, 1'b0};
                        wen_a24 = {1'b0, 1'b0};
                        wen_a23 = {1'b0, 1'b0};
                        wen_a22 = {1'b0, 1'b0};
                        wen_a21 = {1'b0, 1'b0};
                        wen_a20 = {1'b0, 1'b0};
                        wen_a19 = {1'b0, 1'b0};
                        wen_a18 = {1'b0, 1'b0};
                        wen_a17 = {1'b0, 1'b0};
                        wen_a16 = {1'b0, 1'b0};
                        wen_a15 = {1'b0, 1'b0};
                        wen_a14 = {1'b0, 1'b0};
                        wen_a13 = {1'b0, 1'b0};
                        wen_a12 = {1'b0, 1'b0};
                        wen_a11 = {1'b0, 1'b0};
                        wen_a10 = {1'b0, wen};
                        wen_a9 = {1'b0, wen};
                        wen_a8 = {1'b0, wen};
                        wen_a7 = {1'b0, wen};
                        wen_a6 = {1'b0, wen};
                        wen_a5 = {1'b0, wen};
                        wen_a4 = {1'b0, wen};
                        wen_a3 = {1'b0, wen};
                        wen_a2 = {1'b0, 1'b0};
                        wen_a1 = {1'b0, 1'b0};
                        wen_a0 = {1'b0, 1'b0};
                        wen_b0 = {1'b0, 1'b0};
                    end
                    6'b101000, 6'b101001 : begin
                        wen_a42 = {1'b0, 1'b0};
                        wen_a41 = {1'b0, 1'b0};
                        wen_a40 = {1'b0, 1'b0};
                        wen_a39 = {1'b0, 1'b0};
                        wen_a38 = {1'b0, 1'b0};
                        wen_a37 = {1'b0, 1'b0};
                        wen_a36 = {1'b0, 1'b0};
                        wen_a35 = {1'b0, 1'b0};
                        wen_a34 = {1'b0, 1'b0};
                        wen_a33 = {1'b0, 1'b0};
                        wen_a32 = {1'b0, 1'b0};
                        wen_a31 = {1'b0, 1'b0};
                        wen_a30 = {1'b0, 1'b0};
                        wen_a29 = {1'b0, 1'b0};
                        wen_a28 = {1'b0, 1'b0};
                        wen_a27 = {1'b0, 1'b0};
                        wen_a26 = {1'b0, 1'b0};
                        wen_a25 = {1'b0, 1'b0};
                        wen_a24 = {1'b0, 1'b0};
                        wen_a23 = {1'b0, 1'b0};
                        wen_a22 = {1'b0, 1'b0};
                        wen_a21 = {1'b0, 1'b0};
                        wen_a20 = {1'b0, 1'b0};
                        wen_a19 = {1'b0, 1'b0};
                        wen_a18 = {1'b0, 1'b0};
                        wen_a17 = {1'b0, 1'b0};
                        wen_a16 = {1'b0, 1'b0};
                        wen_a15 = {1'b0, 1'b0};
                        wen_a14 = {1'b0, 1'b0};
                        wen_a13 = {1'b0, 1'b0};
                        wen_a12 = {1'b0, 1'b0};
                        wen_a11 = {1'b0, 1'b0};
                        wen_a10 = {1'b0, 1'b0};
                        wen_a9 = {1'b0, 1'b0};
                        wen_a8 = {1'b0, 1'b0};
                        wen_a7 = {1'b0, 1'b0};
                        wen_a6 = {1'b0, 1'b0};
                        wen_a5 = {1'b0, 1'b0};
                        wen_a4 = {1'b0, 1'b0};
                        wen_a3 = {1'b0, 1'b0};
                        wen_a2 = {wen, wen};
                        wen_a1 = {wen, wen};
                        wen_a0 = {1'b0, 1'b0};
                        wen_b0 = {1'b0, 1'b0};
                    end
                    6'b101010 : begin
                        wen_a42 = {1'b0, 1'b0};
                        wen_a41 = {1'b0, 1'b0};
                        wen_a40 = {1'b0, 1'b0};
                        wen_a39 = {1'b0, 1'b0};
                        wen_a38 = {1'b0, 1'b0};
                        wen_a37 = {1'b0, 1'b0};
                        wen_a36 = {1'b0, 1'b0};
                        wen_a35 = {1'b0, 1'b0};
                        wen_a34 = {1'b0, 1'b0};
                        wen_a33 = {1'b0, 1'b0};
                        wen_a32 = {1'b0, 1'b0};
                        wen_a31 = {1'b0, 1'b0};
                        wen_a30 = {1'b0, 1'b0};
                        wen_a29 = {1'b0, 1'b0};
                        wen_a28 = {1'b0, 1'b0};
                        wen_a27 = {1'b0, 1'b0};
                        wen_a26 = {1'b0, 1'b0};
                        wen_a25 = {1'b0, 1'b0};
                        wen_a24 = {1'b0, 1'b0};
                        wen_a23 = {1'b0, 1'b0};
                        wen_a22 = {1'b0, 1'b0};
                        wen_a21 = {1'b0, 1'b0};
                        wen_a20 = {1'b0, 1'b0};
                        wen_a19 = {1'b0, 1'b0};
                        wen_a18 = {1'b0, 1'b0};
                        wen_a17 = {1'b0, 1'b0};
                        wen_a16 = {1'b0, 1'b0};
                        wen_a15 = {1'b0, 1'b0};
                        wen_a14 = {1'b0, 1'b0};
                        wen_a13 = {1'b0, 1'b0};
                        wen_a12 = {1'b0, 1'b0};
                        wen_a11 = {1'b0, 1'b0};
                        wen_a10 = {1'b0, 1'b0};
                        wen_a9 = {1'b0, 1'b0};
                        wen_a8 = {1'b0, 1'b0};
                        wen_a7 = {1'b0, 1'b0};
                        wen_a6 = {1'b0, 1'b0};
                        wen_a5 = {1'b0, 1'b0};
                        wen_a4 = {1'b0, 1'b0};
                        wen_a3 = {1'b0, 1'b0};
                        wen_a2 = {1'b0, 1'b0};
                        wen_a1 = {1'b0, 1'b0};
                        wen_a0 = {wen, wen};
                        wen_b0 = {wen, wen};
                    end
                    default : begin
                        wen_a42 = {1'b0, 1'b0};
                        wen_a41 = {1'b0, 1'b0};
                        wen_a40 = {1'b0, 1'b0};
                        wen_a39 = {1'b0, 1'b0};
                        wen_a38 = {1'b0, 1'b0};
                        wen_a37 = {1'b0, 1'b0};
                        wen_a36 = {1'b0, 1'b0};
                        wen_a35 = {1'b0, 1'b0};
                        wen_a34 = {1'b0, 1'b0};
                        wen_a33 = {1'b0, 1'b0};
                        wen_a32 = {1'b0, 1'b0};
                        wen_a31 = {1'b0, 1'b0};
                        wen_a30 = {1'b0, 1'b0};
                        wen_a29 = {1'b0, 1'b0};
                        wen_a28 = {1'b0, 1'b0};
                        wen_a27 = {1'b0, 1'b0};
                        wen_a26 = {1'b0, 1'b0};
                        wen_a25 = {1'b0, 1'b0};
                        wen_a24 = {1'b0, 1'b0};
                        wen_a23 = {1'b0, 1'b0};
                        wen_a22 = {1'b0, 1'b0};
                        wen_a21 = {1'b0, 1'b0};
                        wen_a20 = {1'b0, 1'b0};
                        wen_a19 = {1'b0, 1'b0};
                        wen_a18 = {1'b0, 1'b0};
                        wen_a17 = {1'b0, 1'b0};
                        wen_a16 = {1'b0, 1'b0};
                        wen_a15 = {1'b0, 1'b0};
                        wen_a14 = {1'b0, 1'b0};
                        wen_a13 = {1'b0, 1'b0};
                        wen_a12 = {1'b0, 1'b0};
                        wen_a11 = {1'b0, 1'b0};
                        wen_a10 = {1'b0, 1'b0};
                        wen_a9 = {1'b0, 1'b0};
                        wen_a8 = {1'b0, 1'b0};
                        wen_a7 = {1'b0, 1'b0};
                        wen_a6 = {1'b0, 1'b0};
                        wen_a5 = {1'b0, 1'b0};
                        wen_a4 = {1'b0, 1'b0};
                        wen_a3 = {1'b0, 1'b0};
                        wen_a2 = {1'b0, 1'b0};
                        wen_a1 = {1'b0, 1'b0};
                        wen_a0 = {1'b0, 1'b0};
                        wen_b0 = {1'b0, 1'b0};
                    end
                endcase

                case (ckRdAddr[14:9])
                    6'b000000, 6'b000001, 6'b000010, 6'b000011,
                    6'b000100, 6'b000101, 6'b000110, 6'b000111,
                    6'b001000, 6'b001001, 6'b001010, 6'b001011,
                    6'b001100, 6'b001101, 6'b001110, 6'b001111,
                    6'b010000, 6'b010001, 6'b010010, 6'b010011,
                    6'b010100, 6'b010101, 6'b010110, 6'b010111,
                    6'b011000, 6'b011001, 6'b011010, 6'b011011,
                    6'b011100, 6'b011101, 6'b011110, 6'b011111 : begin
                        readData = {
                                        readData42[0],
                                        readData41[0],
                                        readData40[0],
                                        readData39[0],
                                        readData38[0],
                                        readData37[0],
                                        readData36[0],
                                        readData35[0],
                                        readData34[0],
                                        readData33[0],
                                        readData32[0],
                                        readData31[0],
                                        readData30[0],
                                        readData29[0],
                                        readData28[0],
                                        readData27[0],
                                        readData26[0],
                                        readData25[0],
                                        readData24[0],
                                        readData23[0],
                                        readData22[0],
                                        readData21[0],
                                        readData20[0],
                                        readData19[0],
                                        readData18[0],
                                        readData17[0],
                                        readData16[0],
                                        readData15[0],
                                        readData14[0],
                                        readData13[0],
                                        readData12[0],
                                        readData11[0]
                        };
                    end
                    6'b100000, 6'b100001, 6'b100010, 6'b100011,
                    6'b100100, 6'b100101, 6'b100110, 6'b100111: begin
                        readData = {
                                        readData10[3:0],
                                        readData9[3:0],
                                        readData8[3:0],
                                        readData7[3:0],
                                        readData6[3:0],
                                        readData5[3:0],
                                        readData4[3:0],
                                        readData3[3:0]
                        };
                    end
                    6'b101000, 6'b101001 : begin
                        readData = {readData2[16:9],readData2[7:0],readData1[16:9],readData1[7:0]};
                    end
                    6'b101010 : begin
                        readData = {readData0[34:27],readData0[25:18],readData0[16:9],readData0[7:0]};
                    end
                    default : begin
                        readData = 32'b0;
                    end
                endcase
            end
            22528: begin
                width44 = 3'b000;
                width43 = 3'b000;
                width42 = 3'b000;
                width41 = 3'b000;
                width40 = 3'b000;
                width39 = 3'b000;
                width38 = 3'b000;
                width37 = 3'b000;
                width36 = 3'b000;
                width35 = 3'b000;
                width34 = 3'b000;
                width33 = 3'b000;
                width32 = 3'b000;
                width31 = 3'b000;
                width30 = 3'b000;
                width29 = 3'b000;
                width28 = 3'b000;
                width27 = 3'b000;
                width26 = 3'b000;
                width25 = 3'b000;
                width24 = 3'b000;
                width23 = 3'b000;
                width22 = 3'b000;
                width21 = 3'b000;
                width20 = 3'b000;
                width19 = 3'b000;
                width18 = 3'b000;
                width17 = 3'b000;
                width16 = 3'b000;
                width15 = 3'b000;
                width14 = 3'b000;
                width13 = 3'b000;
                width12 = 3'b010;
                width11 = 3'b010;
                width10 = 3'b010;
                width9 = 3'b010;
                width8 = 3'b010;
                width7 = 3'b010;
                width6 = 3'b010;
                width5 = 3'b010;
                width4 = 3'b011;
                width3 = 3'b011;
                width2 = 3'b011;
                width1 = 3'b011;

                writeAddr44 = {writeAddr[13:0]};
                writeAddr43 = {writeAddr[13:0]};
                writeAddr42 = {writeAddr[13:0]};
                writeAddr41 = {writeAddr[13:0]};
                writeAddr40 = {writeAddr[13:0]};
                writeAddr39 = {writeAddr[13:0]};
                writeAddr38 = {writeAddr[13:0]};
                writeAddr37 = {writeAddr[13:0]};
                writeAddr36 = {writeAddr[13:0]};
                writeAddr35 = {writeAddr[13:0]};
                writeAddr34 = {writeAddr[13:0]};
                writeAddr33 = {writeAddr[13:0]};
                writeAddr32 = {writeAddr[13:0]};
                writeAddr31 = {writeAddr[13:0]};
                writeAddr30 = {writeAddr[13:0]};
                writeAddr29 = {writeAddr[13:0]};
                writeAddr28 = {writeAddr[13:0]};
                writeAddr27 = {writeAddr[13:0]};
                writeAddr26 = {writeAddr[13:0]};
                writeAddr25 = {writeAddr[13:0]};
                writeAddr24 = {writeAddr[13:0]};
                writeAddr23 = {writeAddr[13:0]};
                writeAddr22 = {writeAddr[13:0]};
                writeAddr21 = {writeAddr[13:0]};
                writeAddr20 = {writeAddr[13:0]};
                writeAddr19 = {writeAddr[13:0]};
                writeAddr18 = {writeAddr[13:0]};
                writeAddr17 = {writeAddr[13:0]};
                writeAddr16 = {writeAddr[13:0]};
                writeAddr15 = {writeAddr[13:0]};
                writeAddr14 = {writeAddr[13:0]};
                writeAddr13 = {writeAddr[13:0]};
                writeAddr12 = {writeAddr[11:0], 2'b0};
                writeAddr11 = {writeAddr[11:0], 2'b0};
                writeAddr10 = {writeAddr[11:0], 2'b0};
                writeAddr9 = {writeAddr[11:0], 2'b0};
                writeAddr8 = {writeAddr[11:0], 2'b0};
                writeAddr7 = {writeAddr[11:0], 2'b0};
                writeAddr6 = {writeAddr[11:0], 2'b0};
                writeAddr5 = {writeAddr[11:0], 2'b0};
                writeAddr4 = {writeAddr[10:0], 3'b0};
                writeAddr3 = {writeAddr[10:0], 3'b0};
                writeAddr2 = {writeAddr[10:0], 3'b0};
                writeAddr1 = {writeAddr[10:0], 3'b0};

                readAddr44 = {writeAddr[13:0]};
                readAddr43 = {writeAddr[13:0]};
                readAddr42 = {writeAddr[13:0]};
                readAddr41 = {writeAddr[13:0]};
                readAddr40 = {writeAddr[13:0]};
                readAddr39 = {writeAddr[13:0]};
                readAddr38 = {writeAddr[13:0]};
                readAddr37 = {writeAddr[13:0]};
                readAddr36 = {writeAddr[13:0]};
                readAddr35 = {writeAddr[13:0]};
                readAddr34 = {writeAddr[13:0]};
                readAddr33 = {writeAddr[13:0]};
                readAddr32 = {writeAddr[13:0]};
                readAddr31 = {writeAddr[13:0]};
                readAddr30 = {writeAddr[13:0]};
                readAddr29 = {writeAddr[13:0]};
                readAddr28 = {writeAddr[13:0]};
                readAddr27 = {writeAddr[13:0]};
                readAddr26 = {writeAddr[13:0]};
                readAddr25 = {writeAddr[13:0]};
                readAddr24 = {writeAddr[13:0]};
                readAddr23 = {writeAddr[13:0]};
                readAddr22 = {writeAddr[13:0]};
                readAddr21 = {writeAddr[13:0]};
                readAddr20 = {writeAddr[13:0]};
                readAddr19 = {writeAddr[13:0]};
                readAddr18 = {writeAddr[13:0]};
                readAddr17 = {writeAddr[13:0]};
                readAddr16 = {writeAddr[13:0]};
                readAddr15 = {writeAddr[13:0]};
                readAddr14 = {writeAddr[13:0]};
                readAddr13 = {writeAddr[13:0]};
                readAddr12  = {readAddr[11:0],  2'b0};
                readAddr11  = {readAddr[11:0],  2'b0};
                readAddr10  = {readAddr[11:0],  2'b0};
                readAddr9  = {readAddr[11:0],  2'b0};
                readAddr8  = {readAddr[11:0],  2'b0};
                readAddr7  = {readAddr[11:0],  2'b0};
                readAddr6  = {readAddr[11:0],  2'b0};
                readAddr5  = {readAddr[11:0],  2'b0};
                readAddr4  = {readAddr[10:0],  3'b0};
                readAddr3  = {readAddr[10:0],  3'b0};
                readAddr2  = {readAddr[10:0],  3'b0};
                readAddr1  = {readAddr[10:0],  3'b0};

                writeData44 = {17'b0, writeData[31]};
                writeData43 = {17'b0, writeData[30]};
                writeData42 = {17'b0, writeData[29]};
                writeData41 = {17'b0, writeData[28]};
                writeData40 = {17'b0, writeData[27]};
                writeData39 = {17'b0, writeData[26]};
                writeData38 = {17'b0, writeData[25]};
                writeData37 = {17'b0, writeData[24]};
                writeData36 = {17'b0, writeData[23]};
                writeData35 = {17'b0, writeData[22]};
                writeData34 = {17'b0, writeData[21]};
                writeData33 = {17'b0, writeData[20]};
                writeData32 = {17'b0, writeData[19]};
                writeData31 = {17'b0, writeData[18]};
                writeData30 = {17'b0, writeData[17]};
                writeData29 = {17'b0, writeData[16]};
                writeData28 = {17'b0, writeData[15]};
                writeData27 = {17'b0, writeData[14]};
                writeData26 = {17'b0, writeData[13]};
                writeData25 = {17'b0, writeData[12]};
                writeData24 = {17'b0, writeData[11]};
                writeData23 = {17'b0, writeData[10]};
                writeData22 = {17'b0, writeData[9]};
                writeData21 = {17'b0, writeData[8]};
                writeData20 = {17'b0, writeData[7]};
                writeData19 = {17'b0, writeData[6]};
                writeData18 = {17'b0, writeData[5]};
                writeData17 = {17'b0, writeData[4]};
                writeData16 = {17'b0, writeData[3]};
                writeData15 = {17'b0, writeData[2]};
                writeData14 = {17'b0, writeData[1]};
                writeData13 = {17'b0, writeData[0]};
                writeData12 = {14'b0, writeData[31:28]};
                writeData11 = {14'b0, writeData[27:24]};
                writeData10 = {14'b0, writeData[23:20]};
                writeData9 = {14'b0, writeData[19:16]};
                writeData8 = {14'b0, writeData[15:12]};
                writeData7 = {14'b0, writeData[11:8]};
                writeData6 = {14'b0, writeData[7:4]};
                writeData5 = {14'b0, writeData[3:0]};
                writeData4 = {10'b0, writeData[31:24]};
                writeData3 = {10'b0, writeData[23:16]};
                writeData2 = {10'b0, writeData[15:8]};
                writeData1 = {10'b0, writeData[7:0]};

                case (writeAddr[14:9])
                    6'b000000, 6'b000001, 6'b000010, 6'b000011,
                    6'b000100, 6'b000101, 6'b000110, 6'b000111,
                    6'b001000, 6'b001001, 6'b001010, 6'b001011,
                    6'b001100, 6'b001101, 6'b001110, 6'b001111,
                    6'b010000, 6'b010001, 6'b010010, 6'b010011,
                    6'b010100, 6'b010101, 6'b010110, 6'b010111,
                    6'b011000, 6'b011001, 6'b011010, 6'b011011,
                    6'b011100, 6'b011101, 6'b011110, 6'b011111 : begin
                        wen_a44 = {1'b0, wen};
                        wen_a43 = {1'b0, wen};
                        wen_a42 = {1'b0, wen};
                        wen_a41 = {1'b0, wen};
                        wen_a40 = {1'b0, wen};
                        wen_a39 = {1'b0, wen};
                        wen_a38 = {1'b0, wen};
                        wen_a37 = {1'b0, wen};
                        wen_a36 = {1'b0, wen};
                        wen_a35 = {1'b0, wen};
                        wen_a34 = {1'b0, wen};
                        wen_a33 = {1'b0, wen};
                        wen_a32 = {1'b0, wen};
                        wen_a31 = {1'b0, wen};
                        wen_a30 = {1'b0, wen};
                        wen_a29 = {1'b0, wen};
                        wen_a28 = {1'b0, wen};
                        wen_a27 = {1'b0, wen};
                        wen_a26 = {1'b0, wen};
                        wen_a25 = {1'b0, wen};
                        wen_a24 = {1'b0, wen};
                        wen_a23 = {1'b0, wen};
                        wen_a22 = {1'b0, wen};
                        wen_a21 = {1'b0, wen};
                        wen_a20 = {1'b0, wen};
                        wen_a19 = {1'b0, wen};
                        wen_a18 = {1'b0, wen};
                        wen_a17 = {1'b0, wen};
                        wen_a16 = {1'b0, wen};
                        wen_a15 = {1'b0, wen};
                        wen_a14 = {1'b0, wen};
                        wen_a13 = {1'b0, wen};
                        wen_a12 = {1'b0, 1'b0};
                        wen_a11 = {1'b0, 1'b0};
                        wen_a10 = {1'b0, 1'b0};
                        wen_a9 = {1'b0, 1'b0};
                        wen_a8 = {1'b0, 1'b0};
                        wen_a7 = {1'b0, 1'b0};
                        wen_a6 = {1'b0, 1'b0};
                        wen_a5 = {1'b0, 1'b0};
                        wen_a4 = {1'b0, 1'b0};
                        wen_a3 = {1'b0, 1'b0};
                        wen_a2 = {1'b0, 1'b0};
                        wen_a1 = {1'b0, 1'b0};
                    end
                    6'b100000, 6'b100001, 6'b100010, 6'b100011,
                    6'b100100, 6'b100101, 6'b100110, 6'b100111: begin
                        wen_a44 = {1'b0, 1'b0};
                        wen_a43 = {1'b0, 1'b0};
                        wen_a42 = {1'b0, 1'b0};
                        wen_a41 = {1'b0, 1'b0};
                        wen_a40 = {1'b0, 1'b0};
                        wen_a39 = {1'b0, 1'b0};
                        wen_a38 = {1'b0, 1'b0};
                        wen_a37 = {1'b0, 1'b0};
                        wen_a36 = {1'b0, 1'b0};
                        wen_a35 = {1'b0, 1'b0};
                        wen_a34 = {1'b0, 1'b0};
                        wen_a33 = {1'b0, 1'b0};
                        wen_a32 = {1'b0, 1'b0};
                        wen_a31 = {1'b0, 1'b0};
                        wen_a30 = {1'b0, 1'b0};
                        wen_a29 = {1'b0, 1'b0};
                        wen_a28 = {1'b0, 1'b0};
                        wen_a27 = {1'b0, 1'b0};
                        wen_a26 = {1'b0, 1'b0};
                        wen_a25 = {1'b0, 1'b0};
                        wen_a24 = {1'b0, 1'b0};
                        wen_a23 = {1'b0, 1'b0};
                        wen_a22 = {1'b0, 1'b0};
                        wen_a21 = {1'b0, 1'b0};
                        wen_a20 = {1'b0, 1'b0};
                        wen_a19 = {1'b0, 1'b0};
                        wen_a18 = {1'b0, 1'b0};
                        wen_a17 = {1'b0, 1'b0};
                        wen_a16 = {1'b0, 1'b0};
                        wen_a15 = {1'b0, 1'b0};
                        wen_a14 = {1'b0, 1'b0};
                        wen_a13 = {1'b0, 1'b0};
                        wen_a12 = {1'b0, wen};
                        wen_a11 = {1'b0, wen};
                        wen_a10 = {1'b0, wen};
                        wen_a9 = {1'b0, wen};
                        wen_a8 = {1'b0, wen};
                        wen_a7 = {1'b0, wen};
                        wen_a6 = {1'b0, wen};
                        wen_a5 = {1'b0, wen};
                        wen_a4 = {1'b0, 1'b0};
                        wen_a3 = {1'b0, 1'b0};
                        wen_a2 = {1'b0, 1'b0};
                        wen_a1 = {1'b0, 1'b0};
                    end
                    6'b101000, 6'b101001, 6'b101010, 6'b101011 : begin
                        wen_a44 = {1'b0, 1'b0};
                        wen_a43 = {1'b0, 1'b0};
                        wen_a42 = {1'b0, 1'b0};
                        wen_a41 = {1'b0, 1'b0};
                        wen_a40 = {1'b0, 1'b0};
                        wen_a39 = {1'b0, 1'b0};
                        wen_a38 = {1'b0, 1'b0};
                        wen_a37 = {1'b0, 1'b0};
                        wen_a36 = {1'b0, 1'b0};
                        wen_a35 = {1'b0, 1'b0};
                        wen_a34 = {1'b0, 1'b0};
                        wen_a33 = {1'b0, 1'b0};
                        wen_a32 = {1'b0, 1'b0};
                        wen_a31 = {1'b0, 1'b0};
                        wen_a30 = {1'b0, 1'b0};
                        wen_a29 = {1'b0, 1'b0};
                        wen_a28 = {1'b0, 1'b0};
                        wen_a27 = {1'b0, 1'b0};
                        wen_a26 = {1'b0, 1'b0};
                        wen_a25 = {1'b0, 1'b0};
                        wen_a24 = {1'b0, 1'b0};
                        wen_a23 = {1'b0, 1'b0};
                        wen_a22 = {1'b0, 1'b0};
                        wen_a21 = {1'b0, 1'b0};
                        wen_a20 = {1'b0, 1'b0};
                        wen_a19 = {1'b0, 1'b0};
                        wen_a18 = {1'b0, 1'b0};
                        wen_a17 = {1'b0, 1'b0};
                        wen_a16 = {1'b0, 1'b0};
                        wen_a15 = {1'b0, 1'b0};
                        wen_a14 = {1'b0, 1'b0};
                        wen_a13 = {1'b0, 1'b0};
                        wen_a12 = {1'b0, 1'b0};
                        wen_a11 = {1'b0, 1'b0};
                        wen_a10 = {1'b0, 1'b0};
                        wen_a9 = {1'b0, 1'b0};
                        wen_a8 = {1'b0, 1'b0};
                        wen_a7 = {1'b0, 1'b0};
                        wen_a6 = {1'b0, 1'b0};
                        wen_a5 = {1'b0, 1'b0};
                        wen_a4 = {1'b0, wen};
                        wen_a3 = {1'b0, wen};
                        wen_a2 = {1'b0, wen};
                        wen_a1 = {1'b0, wen};
                    end
                    default : begin
                        wen_a44 = {1'b0, 1'b0};
                        wen_a43 = {1'b0, 1'b0};
                        wen_a42 = {1'b0, 1'b0};
                        wen_a41 = {1'b0, 1'b0};
                        wen_a40 = {1'b0, 1'b0};
                        wen_a39 = {1'b0, 1'b0};
                        wen_a38 = {1'b0, 1'b0};
                        wen_a37 = {1'b0, 1'b0};
                        wen_a36 = {1'b0, 1'b0};
                        wen_a35 = {1'b0, 1'b0};
                        wen_a34 = {1'b0, 1'b0};
                        wen_a33 = {1'b0, 1'b0};
                        wen_a32 = {1'b0, 1'b0};
                        wen_a31 = {1'b0, 1'b0};
                        wen_a30 = {1'b0, 1'b0};
                        wen_a29 = {1'b0, 1'b0};
                        wen_a28 = {1'b0, 1'b0};
                        wen_a27 = {1'b0, 1'b0};
                        wen_a26 = {1'b0, 1'b0};
                        wen_a25 = {1'b0, 1'b0};
                        wen_a24 = {1'b0, 1'b0};
                        wen_a23 = {1'b0, 1'b0};
                        wen_a22 = {1'b0, 1'b0};
                        wen_a21 = {1'b0, 1'b0};
                        wen_a20 = {1'b0, 1'b0};
                        wen_a19 = {1'b0, 1'b0};
                        wen_a18 = {1'b0, 1'b0};
                        wen_a17 = {1'b0, 1'b0};
                        wen_a16 = {1'b0, 1'b0};
                        wen_a15 = {1'b0, 1'b0};
                        wen_a14 = {1'b0, 1'b0};
                        wen_a13 = {1'b0, 1'b0};
                        wen_a12 = {1'b0, 1'b0};
                        wen_a11 = {1'b0, 1'b0};
                        wen_a10 = {1'b0, 1'b0};
                        wen_a9 = {1'b0, 1'b0};
                        wen_a8 = {1'b0, 1'b0};
                        wen_a7 = {1'b0, 1'b0};
                        wen_a6 = {1'b0, 1'b0};
                        wen_a5 = {1'b0, 1'b0};
                        wen_a4 = {1'b0, 1'b0};
                        wen_a3 = {1'b0, 1'b0};
                        wen_a2 = {1'b0, 1'b0};
                        wen_a1 = {1'b0, 1'b0};
                    end
                endcase

                case (ckRdAddr[14:9])
                    6'b000000, 6'b000001, 6'b000010, 6'b000011,
                    6'b000100, 6'b000101, 6'b000110, 6'b000111,
                    6'b001000, 6'b001001, 6'b001010, 6'b001011,
                    6'b001100, 6'b001101, 6'b001110, 6'b001111,
                    6'b010000, 6'b010001, 6'b010010, 6'b010011,
                    6'b010100, 6'b010101, 6'b010110, 6'b010111,
                    6'b011000, 6'b011001, 6'b011010, 6'b011011,
                    6'b011100, 6'b011101, 6'b011110, 6'b011111 : begin
                        readData = {
                                        readData44[0],
                                        readData43[0],
                                        readData42[0],
                                        readData41[0],
                                        readData40[0],
                                        readData39[0],
                                        readData38[0],
                                        readData37[0],
                                        readData36[0],
                                        readData35[0],
                                        readData34[0],
                                        readData33[0],
                                        readData32[0],
                                        readData31[0],
                                        readData30[0],
                                        readData29[0],
                                        readData28[0],
                                        readData27[0],
                                        readData26[0],
                                        readData25[0],
                                        readData24[0],
                                        readData23[0],
                                        readData22[0],
                                        readData21[0],
                                        readData20[0],
                                        readData19[0],
                                        readData18[0],
                                        readData17[0],
                                        readData16[0],
                                        readData15[0],
                                        readData14[0],
                                        readData13[0]
                        };
                    end
                    6'b100000, 6'b100001, 6'b100010, 6'b100011,
                    6'b100100, 6'b100101, 6'b100110, 6'b100111: begin
                        readData = {
                                        readData12[3:0],
                                        readData11[3:0],
                                        readData10[3:0],
                                        readData9[3:0],
                                        readData8[3:0],
                                        readData7[3:0],
                                        readData6[3:0],
                                        readData5[3:0]
                        };
                    end
                    6'b101000, 6'b101001, 6'b101010, 6'b101011: begin
                        readData = {readData4[7:0],readData3[7:0],readData2[7:0],readData1[7:0]};
                    end
                    default : begin
                        readData = 32'b0;
                    end
                endcase
            end
            23040: begin
                width44 = 3'b000;
                width43 = 3'b000;
                width42 = 3'b000;
                width41 = 3'b000;
                width40 = 3'b000;
                width39 = 3'b000;
                width38 = 3'b000;
                width37 = 3'b000;
                width36 = 3'b000;
                width35 = 3'b000;
                width34 = 3'b000;
                width33 = 3'b000;
                width32 = 3'b000;
                width31 = 3'b000;
                width30 = 3'b000;
                width29 = 3'b000;
                width28 = 3'b000;
                width27 = 3'b000;
                width26 = 3'b000;
                width25 = 3'b000;
                width24 = 3'b000;
                width23 = 3'b000;
                width22 = 3'b000;
                width21 = 3'b000;
                width20 = 3'b000;
                width19 = 3'b000;
                width18 = 3'b000;
                width17 = 3'b000;
                width16 = 3'b000;
                width15 = 3'b000;
                width14 = 3'b000;
                width13 = 3'b000;
                width12 = 3'b010;
                width11 = 3'b010;
                width10 = 3'b010;
                width9 = 3'b010;
                width8 = 3'b010;
                width7 = 3'b010;
                width6 = 3'b010;
                width5 = 3'b010;
                width4 = 3'b011;
                width3 = 3'b011;
                width2 = 3'b011;
                width1 = 3'b011;
                width0 = 3'b101;

                writeAddr44 = {writeAddr[13:0]};
                writeAddr43 = {writeAddr[13:0]};
                writeAddr42 = {writeAddr[13:0]};
                writeAddr41 = {writeAddr[13:0]};
                writeAddr40 = {writeAddr[13:0]};
                writeAddr39 = {writeAddr[13:0]};
                writeAddr38 = {writeAddr[13:0]};
                writeAddr37 = {writeAddr[13:0]};
                writeAddr36 = {writeAddr[13:0]};
                writeAddr35 = {writeAddr[13:0]};
                writeAddr34 = {writeAddr[13:0]};
                writeAddr33 = {writeAddr[13:0]};
                writeAddr32 = {writeAddr[13:0]};
                writeAddr31 = {writeAddr[13:0]};
                writeAddr30 = {writeAddr[13:0]};
                writeAddr29 = {writeAddr[13:0]};
                writeAddr28 = {writeAddr[13:0]};
                writeAddr27 = {writeAddr[13:0]};
                writeAddr26 = {writeAddr[13:0]};
                writeAddr25 = {writeAddr[13:0]};
                writeAddr24 = {writeAddr[13:0]};
                writeAddr23 = {writeAddr[13:0]};
                writeAddr22 = {writeAddr[13:0]};
                writeAddr21 = {writeAddr[13:0]};
                writeAddr20 = {writeAddr[13:0]};
                writeAddr19 = {writeAddr[13:0]};
                writeAddr18 = {writeAddr[13:0]};
                writeAddr17 = {writeAddr[13:0]};
                writeAddr16 = {writeAddr[13:0]};
                writeAddr15 = {writeAddr[13:0]};
                writeAddr14 = {writeAddr[13:0]};
                writeAddr13 = {writeAddr[13:0]};
                writeAddr12 = {writeAddr[11:0], 2'b0};
                writeAddr11 = {writeAddr[11:0], 2'b0};
                writeAddr10 = {writeAddr[11:0], 2'b0};
                writeAddr9 = {writeAddr[11:0], 2'b0};
                writeAddr8 = {writeAddr[11:0], 2'b0};
                writeAddr7 = {writeAddr[11:0], 2'b0};
                writeAddr6 = {writeAddr[11:0], 2'b0};
                writeAddr5 = {writeAddr[11:0], 2'b0};
                writeAddr4 = {writeAddr[10:0], 3'b0};
                writeAddr3 = {writeAddr[10:0], 3'b0};
                writeAddr2 = {writeAddr[10:0], 3'b0};
                writeAddr1 = {writeAddr[10:0], 3'b0};
                writeAddr0 = {writeAddr[8:0], 5'b0};

                readAddr44 = {writeAddr[13:0]};
                readAddr43 = {writeAddr[13:0]};
                readAddr42 = {writeAddr[13:0]};
                readAddr41 = {writeAddr[13:0]};
                readAddr40 = {writeAddr[13:0]};
                readAddr39 = {writeAddr[13:0]};
                readAddr38 = {writeAddr[13:0]};
                readAddr37 = {writeAddr[13:0]};
                readAddr36 = {writeAddr[13:0]};
                readAddr35 = {writeAddr[13:0]};
                readAddr34 = {writeAddr[13:0]};
                readAddr33 = {writeAddr[13:0]};
                readAddr32 = {writeAddr[13:0]};
                readAddr31 = {writeAddr[13:0]};
                readAddr30 = {writeAddr[13:0]};
                readAddr29 = {writeAddr[13:0]};
                readAddr28 = {writeAddr[13:0]};
                readAddr27 = {writeAddr[13:0]};
                readAddr26 = {writeAddr[13:0]};
                readAddr25 = {writeAddr[13:0]};
                readAddr24 = {writeAddr[13:0]};
                readAddr23 = {writeAddr[13:0]};
                readAddr22 = {writeAddr[13:0]};
                readAddr21 = {writeAddr[13:0]};
                readAddr20 = {writeAddr[13:0]};
                readAddr19 = {writeAddr[13:0]};
                readAddr18 = {writeAddr[13:0]};
                readAddr17 = {writeAddr[13:0]};
                readAddr16 = {writeAddr[13:0]};
                readAddr15 = {writeAddr[13:0]};
                readAddr14 = {writeAddr[13:0]};
                readAddr13 = {writeAddr[13:0]};
                readAddr12  = {readAddr[11:0],  2'b0};
                readAddr11  = {readAddr[11:0],  2'b0};
                readAddr10  = {readAddr[11:0],  2'b0};
                readAddr9  = {readAddr[11:0],  2'b0};
                readAddr8  = {readAddr[11:0],  2'b0};
                readAddr7  = {readAddr[11:0],  2'b0};
                readAddr6  = {readAddr[11:0],  2'b0};
                readAddr5  = {readAddr[11:0],  2'b0};
                readAddr4  = {readAddr[10:0],  3'b0};
                readAddr3  = {readAddr[10:0],  3'b0};
                readAddr2  = {readAddr[10:0],  3'b0};
                readAddr1  = {readAddr[10:0],  3'b0};
                readAddr0  = {readAddr[8:0],  5'b0};

                writeData44 = {17'b0, writeData[31]};
                writeData43 = {17'b0, writeData[30]};
                writeData42 = {17'b0, writeData[29]};
                writeData41 = {17'b0, writeData[28]};
                writeData40 = {17'b0, writeData[27]};
                writeData39 = {17'b0, writeData[26]};
                writeData38 = {17'b0, writeData[25]};
                writeData37 = {17'b0, writeData[24]};
                writeData36 = {17'b0, writeData[23]};
                writeData35 = {17'b0, writeData[22]};
                writeData34 = {17'b0, writeData[21]};
                writeData33 = {17'b0, writeData[20]};
                writeData32 = {17'b0, writeData[19]};
                writeData31 = {17'b0, writeData[18]};
                writeData30 = {17'b0, writeData[17]};
                writeData29 = {17'b0, writeData[16]};
                writeData28 = {17'b0, writeData[15]};
                writeData27 = {17'b0, writeData[14]};
                writeData26 = {17'b0, writeData[13]};
                writeData25 = {17'b0, writeData[12]};
                writeData24 = {17'b0, writeData[11]};
                writeData23 = {17'b0, writeData[10]};
                writeData22 = {17'b0, writeData[9]};
                writeData21 = {17'b0, writeData[8]};
                writeData20 = {17'b0, writeData[7]};
                writeData19 = {17'b0, writeData[6]};
                writeData18 = {17'b0, writeData[5]};
                writeData17 = {17'b0, writeData[4]};
                writeData16 = {17'b0, writeData[3]};
                writeData15 = {17'b0, writeData[2]};
                writeData14 = {17'b0, writeData[1]};
                writeData13 = {17'b0, writeData[0]};
                writeData12 = {14'b0, writeData[31:28]};
                writeData11 = {14'b0, writeData[27:24]};
                writeData10 = {14'b0, writeData[23:20]};
                writeData9 = {14'b0, writeData[19:16]};
                writeData8 = {14'b0, writeData[15:12]};
                writeData7 = {14'b0, writeData[11:8]};
                writeData6 = {14'b0, writeData[7:4]};
                writeData5 = {14'b0, writeData[3:0]};
                writeData4 = {10'b0, writeData[31:24]};
                writeData3 = {10'b0, writeData[23:16]};
                writeData2 = {10'b0, writeData[15:8]};
                writeData1 = {10'b0, writeData[7:0]};
                writeData0 = {1'b0, writeData[31:24], 1'b0, writeData[23:16], 1'b0, writeData[15:8], 1'b0, writeData[7:0]};

                case (writeAddr[14:9])
                    6'b000000, 6'b000001, 6'b000010, 6'b000011,
                    6'b000100, 6'b000101, 6'b000110, 6'b000111,
                    6'b001000, 6'b001001, 6'b001010, 6'b001011,
                    6'b001100, 6'b001101, 6'b001110, 6'b001111,
                    6'b010000, 6'b010001, 6'b010010, 6'b010011,
                    6'b010100, 6'b010101, 6'b010110, 6'b010111,
                    6'b011000, 6'b011001, 6'b011010, 6'b011011,
                    6'b011100, 6'b011101, 6'b011110, 6'b011111 : begin
                        wen_a44 = {1'b0, wen};
                        wen_a43 = {1'b0, wen};
                        wen_a42 = {1'b0, wen};
                        wen_a41 = {1'b0, wen};
                        wen_a40 = {1'b0, wen};
                        wen_a39 = {1'b0, wen};
                        wen_a38 = {1'b0, wen};
                        wen_a37 = {1'b0, wen};
                        wen_a36 = {1'b0, wen};
                        wen_a35 = {1'b0, wen};
                        wen_a34 = {1'b0, wen};
                        wen_a33 = {1'b0, wen};
                        wen_a32 = {1'b0, wen};
                        wen_a31 = {1'b0, wen};
                        wen_a30 = {1'b0, wen};
                        wen_a29 = {1'b0, wen};
                        wen_a28 = {1'b0, wen};
                        wen_a27 = {1'b0, wen};
                        wen_a26 = {1'b0, wen};
                        wen_a25 = {1'b0, wen};
                        wen_a24 = {1'b0, wen};
                        wen_a23 = {1'b0, wen};
                        wen_a22 = {1'b0, wen};
                        wen_a21 = {1'b0, wen};
                        wen_a20 = {1'b0, wen};
                        wen_a19 = {1'b0, wen};
                        wen_a18 = {1'b0, wen};
                        wen_a17 = {1'b0, wen};
                        wen_a16 = {1'b0, wen};
                        wen_a15 = {1'b0, wen};
                        wen_a14 = {1'b0, wen};
                        wen_a13 = {1'b0, wen};
                        wen_a12 = {1'b0, 1'b0};
                        wen_a11 = {1'b0, 1'b0};
                        wen_a10 = {1'b0, 1'b0};
                        wen_a9 = {1'b0, 1'b0};
                        wen_a8 = {1'b0, 1'b0};
                        wen_a7 = {1'b0, 1'b0};
                        wen_a6 = {1'b0, 1'b0};
                        wen_a5 = {1'b0, 1'b0};
                        wen_a4 = {1'b0, 1'b0};
                        wen_a3 = {1'b0, 1'b0};
                        wen_a2 = {1'b0, 1'b0};
                        wen_a1 = {1'b0, 1'b0};
                        wen_a0 = {1'b0, 1'b0};
                        wen_b0 = {1'b0, 1'b0};
                    end
                    6'b100000, 6'b100001, 6'b100010, 6'b100011,
                    6'b100100, 6'b100101, 6'b100110, 6'b100111: begin
                        wen_a44 = {1'b0, 1'b0};
                        wen_a43 = {1'b0, 1'b0};
                        wen_a42 = {1'b0, 1'b0};
                        wen_a41 = {1'b0, 1'b0};
                        wen_a40 = {1'b0, 1'b0};
                        wen_a39 = {1'b0, 1'b0};
                        wen_a38 = {1'b0, 1'b0};
                        wen_a37 = {1'b0, 1'b0};
                        wen_a36 = {1'b0, 1'b0};
                        wen_a35 = {1'b0, 1'b0};
                        wen_a34 = {1'b0, 1'b0};
                        wen_a33 = {1'b0, 1'b0};
                        wen_a32 = {1'b0, 1'b0};
                        wen_a31 = {1'b0, 1'b0};
                        wen_a30 = {1'b0, 1'b0};
                        wen_a29 = {1'b0, 1'b0};
                        wen_a28 = {1'b0, 1'b0};
                        wen_a27 = {1'b0, 1'b0};
                        wen_a26 = {1'b0, 1'b0};
                        wen_a25 = {1'b0, 1'b0};
                        wen_a24 = {1'b0, 1'b0};
                        wen_a23 = {1'b0, 1'b0};
                        wen_a22 = {1'b0, 1'b0};
                        wen_a21 = {1'b0, 1'b0};
                        wen_a20 = {1'b0, 1'b0};
                        wen_a19 = {1'b0, 1'b0};
                        wen_a18 = {1'b0, 1'b0};
                        wen_a17 = {1'b0, 1'b0};
                        wen_a16 = {1'b0, 1'b0};
                        wen_a15 = {1'b0, 1'b0};
                        wen_a14 = {1'b0, 1'b0};
                        wen_a13 = {1'b0, 1'b0};
                        wen_a12 = {1'b0, wen};
                        wen_a11 = {1'b0, wen};
                        wen_a10 = {1'b0, wen};
                        wen_a9 = {1'b0, wen};
                        wen_a8 = {1'b0, wen};
                        wen_a7 = {1'b0, wen};
                        wen_a6 = {1'b0, wen};
                        wen_a5 = {1'b0, wen};
                        wen_a4 = {1'b0, 1'b0};
                        wen_a3 = {1'b0, 1'b0};
                        wen_a2 = {1'b0, 1'b0};
                        wen_a1 = {1'b0, 1'b0};
                        wen_a0 = {1'b0, 1'b0};
                        wen_b0 = {1'b0, 1'b0};
                    end
                    6'b101000, 6'b101001, 6'b101010, 6'b101011 : begin
                        wen_a44 = {1'b0, 1'b0};
                        wen_a43 = {1'b0, 1'b0};
                        wen_a42 = {1'b0, 1'b0};
                        wen_a41 = {1'b0, 1'b0};
                        wen_a40 = {1'b0, 1'b0};
                        wen_a39 = {1'b0, 1'b0};
                        wen_a38 = {1'b0, 1'b0};
                        wen_a37 = {1'b0, 1'b0};
                        wen_a36 = {1'b0, 1'b0};
                        wen_a35 = {1'b0, 1'b0};
                        wen_a34 = {1'b0, 1'b0};
                        wen_a33 = {1'b0, 1'b0};
                        wen_a32 = {1'b0, 1'b0};
                        wen_a31 = {1'b0, 1'b0};
                        wen_a30 = {1'b0, 1'b0};
                        wen_a29 = {1'b0, 1'b0};
                        wen_a28 = {1'b0, 1'b0};
                        wen_a27 = {1'b0, 1'b0};
                        wen_a26 = {1'b0, 1'b0};
                        wen_a25 = {1'b0, 1'b0};
                        wen_a24 = {1'b0, 1'b0};
                        wen_a23 = {1'b0, 1'b0};
                        wen_a22 = {1'b0, 1'b0};
                        wen_a21 = {1'b0, 1'b0};
                        wen_a20 = {1'b0, 1'b0};
                        wen_a19 = {1'b0, 1'b0};
                        wen_a18 = {1'b0, 1'b0};
                        wen_a17 = {1'b0, 1'b0};
                        wen_a16 = {1'b0, 1'b0};
                        wen_a15 = {1'b0, 1'b0};
                        wen_a14 = {1'b0, 1'b0};
                        wen_a13 = {1'b0, 1'b0};
                        wen_a12 = {1'b0, 1'b0};
                        wen_a11 = {1'b0, 1'b0};
                        wen_a10 = {1'b0, 1'b0};
                        wen_a9 = {1'b0, 1'b0};
                        wen_a8 = {1'b0, 1'b0};
                        wen_a7 = {1'b0, 1'b0};
                        wen_a6 = {1'b0, 1'b0};
                        wen_a5 = {1'b0, 1'b0};
                        wen_a4 = {1'b0, wen};
                        wen_a3 = {1'b0, wen};
                        wen_a2 = {1'b0, wen};
                        wen_a1 = {1'b0, wen};
                        wen_a0 = {1'b0, 1'b0};
                        wen_b0 = {1'b0, 1'b0};
                    end
                    6'b101100 : begin
                        wen_a44 = {1'b0, 1'b0};
                        wen_a43 = {1'b0, 1'b0};
                        wen_a42 = {1'b0, 1'b0};
                        wen_a41 = {1'b0, 1'b0};
                        wen_a40 = {1'b0, 1'b0};
                        wen_a39 = {1'b0, 1'b0};
                        wen_a38 = {1'b0, 1'b0};
                        wen_a37 = {1'b0, 1'b0};
                        wen_a36 = {1'b0, 1'b0};
                        wen_a35 = {1'b0, 1'b0};
                        wen_a34 = {1'b0, 1'b0};
                        wen_a33 = {1'b0, 1'b0};
                        wen_a32 = {1'b0, 1'b0};
                        wen_a31 = {1'b0, 1'b0};
                        wen_a30 = {1'b0, 1'b0};
                        wen_a29 = {1'b0, 1'b0};
                        wen_a28 = {1'b0, 1'b0};
                        wen_a27 = {1'b0, 1'b0};
                        wen_a26 = {1'b0, 1'b0};
                        wen_a25 = {1'b0, 1'b0};
                        wen_a24 = {1'b0, 1'b0};
                        wen_a23 = {1'b0, 1'b0};
                        wen_a22 = {1'b0, 1'b0};
                        wen_a21 = {1'b0, 1'b0};
                        wen_a20 = {1'b0, 1'b0};
                        wen_a19 = {1'b0, 1'b0};
                        wen_a18 = {1'b0, 1'b0};
                        wen_a17 = {1'b0, 1'b0};
                        wen_a16 = {1'b0, 1'b0};
                        wen_a15 = {1'b0, 1'b0};
                        wen_a14 = {1'b0, 1'b0};
                        wen_a13 = {1'b0, 1'b0};
                        wen_a12 = {1'b0, 1'b0};
                        wen_a11 = {1'b0, 1'b0};
                        wen_a10 = {1'b0, 1'b0};
                        wen_a9 = {1'b0, 1'b0};
                        wen_a8 = {1'b0, 1'b0};
                        wen_a7 = {1'b0, 1'b0};
                        wen_a6 = {1'b0, 1'b0};
                        wen_a5 = {1'b0, 1'b0};
                        wen_a4 = {1'b0, 1'b0};
                        wen_a3 = {1'b0, 1'b0};
                        wen_a2 = {1'b0, 1'b0};
                        wen_a1 = {1'b0, 1'b0};
                        wen_a0 = {wen, wen};
                        wen_b0 = {wen, wen};
                    end
                    default : begin
                        wen_a44 = {1'b0, 1'b0};
                        wen_a43 = {1'b0, 1'b0};
                        wen_a42 = {1'b0, 1'b0};
                        wen_a41 = {1'b0, 1'b0};
                        wen_a40 = {1'b0, 1'b0};
                        wen_a39 = {1'b0, 1'b0};
                        wen_a38 = {1'b0, 1'b0};
                        wen_a37 = {1'b0, 1'b0};
                        wen_a36 = {1'b0, 1'b0};
                        wen_a35 = {1'b0, 1'b0};
                        wen_a34 = {1'b0, 1'b0};
                        wen_a33 = {1'b0, 1'b0};
                        wen_a32 = {1'b0, 1'b0};
                        wen_a31 = {1'b0, 1'b0};
                        wen_a30 = {1'b0, 1'b0};
                        wen_a29 = {1'b0, 1'b0};
                        wen_a28 = {1'b0, 1'b0};
                        wen_a27 = {1'b0, 1'b0};
                        wen_a26 = {1'b0, 1'b0};
                        wen_a25 = {1'b0, 1'b0};
                        wen_a24 = {1'b0, 1'b0};
                        wen_a23 = {1'b0, 1'b0};
                        wen_a22 = {1'b0, 1'b0};
                        wen_a21 = {1'b0, 1'b0};
                        wen_a20 = {1'b0, 1'b0};
                        wen_a19 = {1'b0, 1'b0};
                        wen_a18 = {1'b0, 1'b0};
                        wen_a17 = {1'b0, 1'b0};
                        wen_a16 = {1'b0, 1'b0};
                        wen_a15 = {1'b0, 1'b0};
                        wen_a14 = {1'b0, 1'b0};
                        wen_a13 = {1'b0, 1'b0};
                        wen_a12 = {1'b0, 1'b0};
                        wen_a11 = {1'b0, 1'b0};
                        wen_a10 = {1'b0, 1'b0};
                        wen_a9 = {1'b0, 1'b0};
                        wen_a8 = {1'b0, 1'b0};
                        wen_a7 = {1'b0, 1'b0};
                        wen_a6 = {1'b0, 1'b0};
                        wen_a5 = {1'b0, 1'b0};
                        wen_a4 = {1'b0, 1'b0};
                        wen_a3 = {1'b0, 1'b0};
                        wen_a2 = {1'b0, 1'b0};
                        wen_a1 = {1'b0, 1'b0};
                        wen_a0 = {1'b0, 1'b0};
                        wen_b0 = {1'b0, 1'b0};
                    end
                endcase

                case (ckRdAddr[14:9])
                    6'b000000, 6'b000001, 6'b000010, 6'b000011,
                    6'b000100, 6'b000101, 6'b000110, 6'b000111,
                    6'b001000, 6'b001001, 6'b001010, 6'b001011,
                    6'b001100, 6'b001101, 6'b001110, 6'b001111,
                    6'b010000, 6'b010001, 6'b010010, 6'b010011,
                    6'b010100, 6'b010101, 6'b010110, 6'b010111,
                    6'b011000, 6'b011001, 6'b011010, 6'b011011,
                    6'b011100, 6'b011101, 6'b011110, 6'b011111 : begin
                        readData = {
                                        readData44[0],
                                        readData43[0],
                                        readData42[0],
                                        readData41[0],
                                        readData40[0],
                                        readData39[0],
                                        readData38[0],
                                        readData37[0],
                                        readData36[0],
                                        readData35[0],
                                        readData34[0],
                                        readData33[0],
                                        readData32[0],
                                        readData31[0],
                                        readData30[0],
                                        readData29[0],
                                        readData28[0],
                                        readData27[0],
                                        readData26[0],
                                        readData25[0],
                                        readData24[0],
                                        readData23[0],
                                        readData22[0],
                                        readData21[0],
                                        readData20[0],
                                        readData19[0],
                                        readData18[0],
                                        readData17[0],
                                        readData16[0],
                                        readData15[0],
                                        readData14[0],
                                        readData13[0]
                        };
                    end
                    6'b100000, 6'b100001, 6'b100010, 6'b100011,
                    6'b100100, 6'b100101, 6'b100110, 6'b100111: begin
                        readData = {
                                        readData12[3:0],
                                        readData11[3:0],
                                        readData10[3:0],
                                        readData9[3:0],
                                        readData8[3:0],
                                        readData7[3:0],
                                        readData6[3:0],
                                        readData5[3:0]
                        };
                    end
                    6'b101000, 6'b101001, 6'b101010, 6'b101011 : begin
                        readData = {readData4[7:0],readData3[7:0],readData2[7:0],readData1[7:0]};
                    end
                    6'b101100 : begin
                        readData = {readData0[34:27],readData0[25:18],readData0[16:9],readData0[7:0]};
                    end
                    default : begin
                        readData = 32'b0;
                    end
                endcase
            end
            23552: begin
                width46 = 3'b000;
                width45 = 3'b000;
                width44 = 3'b000;
                width43 = 3'b000;
                width42 = 3'b000;
                width41 = 3'b000;
                width40 = 3'b000;
                width39 = 3'b000;
                width38 = 3'b000;
                width37 = 3'b000;
                width36 = 3'b000;
                width35 = 3'b000;
                width34 = 3'b000;
                width33 = 3'b000;
                width32 = 3'b000;
                width31 = 3'b000;
                width30 = 3'b000;
                width29 = 3'b000;
                width28 = 3'b000;
                width27 = 3'b000;
                width26 = 3'b000;
                width25 = 3'b000;
                width24 = 3'b000;
                width23 = 3'b000;
                width22 = 3'b000;
                width21 = 3'b000;
                width20 = 3'b000;
                width19 = 3'b000;
                width18 = 3'b000;
                width17 = 3'b000;
                width16 = 3'b000;
                width15 = 3'b000;
                width14 = 3'b010;
                width13 = 3'b010;
                width12 = 3'b010;
                width11 = 3'b010;
                width10 = 3'b010;
                width9 = 3'b010;
                width8 = 3'b010;
                width7 = 3'b010;
                width6 = 3'b011;
                width5 = 3'b011;
                width4 = 3'b011;
                width3 = 3'b011;
                width2 = 3'b100;
                width1 = 3'b100;

                writeAddr46 = {writeAddr[13:0]};
                writeAddr45 = {writeAddr[13:0]};
                writeAddr44 = {writeAddr[13:0]};
                writeAddr43 = {writeAddr[13:0]};
                writeAddr42 = {writeAddr[13:0]};
                writeAddr41 = {writeAddr[13:0]};
                writeAddr40 = {writeAddr[13:0]};
                writeAddr39 = {writeAddr[13:0]};
                writeAddr38 = {writeAddr[13:0]};
                writeAddr37 = {writeAddr[13:0]};
                writeAddr36 = {writeAddr[13:0]};
                writeAddr35 = {writeAddr[13:0]};
                writeAddr34 = {writeAddr[13:0]};
                writeAddr33 = {writeAddr[13:0]};
                writeAddr32 = {writeAddr[13:0]};
                writeAddr31 = {writeAddr[13:0]};
                writeAddr30 = {writeAddr[13:0]};
                writeAddr29 = {writeAddr[13:0]};
                writeAddr28 = {writeAddr[13:0]};
                writeAddr27 = {writeAddr[13:0]};
                writeAddr26 = {writeAddr[13:0]};
                writeAddr25 = {writeAddr[13:0]};
                writeAddr24 = {writeAddr[13:0]};
                writeAddr23 = {writeAddr[13:0]};
                writeAddr22 = {writeAddr[13:0]};
                writeAddr21 = {writeAddr[13:0]};
                writeAddr20 = {writeAddr[13:0]};
                writeAddr19 = {writeAddr[13:0]};
                writeAddr18 = {writeAddr[13:0]};
                writeAddr17 = {writeAddr[13:0]};
                writeAddr16 = {writeAddr[13:0]};
                writeAddr15 = {writeAddr[13:0]};
                writeAddr14 = {writeAddr[11:0], 2'b0};
                writeAddr13 = {writeAddr[11:0], 2'b0};
                writeAddr12 = {writeAddr[11:0], 2'b0};
                writeAddr11 = {writeAddr[11:0], 2'b0};
                writeAddr10 = {writeAddr[11:0], 2'b0};
                writeAddr9 = {writeAddr[11:0], 2'b0};
                writeAddr8 = {writeAddr[11:0], 2'b0};
                writeAddr7 = {writeAddr[11:0], 2'b0};
                writeAddr6 = {writeAddr[10:0], 3'b0};
                writeAddr5 = {writeAddr[10:0], 3'b0};
                writeAddr4 = {writeAddr[10:0], 3'b0};
                writeAddr3 = {writeAddr[10:0], 3'b0};
                writeAddr2 = {writeAddr[9:0], 4'b0};
                writeAddr1 = {writeAddr[9:0], 4'b0};

                readAddr46 = {writeAddr[13:0]};
                readAddr45 = {writeAddr[13:0]};
                readAddr44 = {writeAddr[13:0]};
                readAddr43 = {writeAddr[13:0]};
                readAddr42 = {writeAddr[13:0]};
                readAddr41 = {writeAddr[13:0]};
                readAddr40 = {writeAddr[13:0]};
                readAddr39 = {writeAddr[13:0]};
                readAddr38 = {writeAddr[13:0]};
                readAddr37 = {writeAddr[13:0]};
                readAddr36 = {writeAddr[13:0]};
                readAddr35 = {writeAddr[13:0]};
                readAddr34 = {writeAddr[13:0]};
                readAddr33 = {writeAddr[13:0]};
                readAddr32 = {writeAddr[13:0]};
                readAddr31 = {writeAddr[13:0]};
                readAddr30 = {writeAddr[13:0]};
                readAddr29 = {writeAddr[13:0]};
                readAddr28 = {writeAddr[13:0]};
                readAddr27 = {writeAddr[13:0]};
                readAddr26 = {writeAddr[13:0]};
                readAddr25 = {writeAddr[13:0]};
                readAddr24 = {writeAddr[13:0]};
                readAddr23 = {writeAddr[13:0]};
                readAddr22 = {writeAddr[13:0]};
                readAddr21 = {writeAddr[13:0]};
                readAddr20 = {writeAddr[13:0]};
                readAddr19 = {writeAddr[13:0]};
                readAddr18 = {writeAddr[13:0]};
                readAddr17 = {writeAddr[13:0]};
                readAddr16 = {writeAddr[13:0]};
                readAddr15 = {writeAddr[13:0]};
                readAddr14  = {readAddr[11:0],  2'b0};
                readAddr13  = {readAddr[11:0],  2'b0};
                readAddr12  = {readAddr[11:0],  2'b0};
                readAddr11  = {readAddr[11:0],  2'b0};
                readAddr10  = {readAddr[11:0],  2'b0};
                readAddr9  = {readAddr[11:0],  2'b0};
                readAddr8  = {readAddr[11:0],  2'b0};
                readAddr7  = {readAddr[11:0],  2'b0};
                readAddr6  = {readAddr[10:0],  3'b0};
                readAddr5  = {readAddr[10:0],  3'b0};
                readAddr4  = {readAddr[10:0],  3'b0};
                readAddr3  = {readAddr[10:0],  3'b0};
                readAddr2  = {readAddr[9:0],  4'b0};
                readAddr1  = {readAddr[9:0],  4'b0};

                writeData46 = {17'b0, writeData[31]};
                writeData45 = {17'b0, writeData[30]};
                writeData44 = {17'b0, writeData[29]};
                writeData43 = {17'b0, writeData[28]};
                writeData42 = {17'b0, writeData[27]};
                writeData41 = {17'b0, writeData[26]};
                writeData40 = {17'b0, writeData[25]};
                writeData39 = {17'b0, writeData[24]};
                writeData38 = {17'b0, writeData[23]};
                writeData37 = {17'b0, writeData[22]};
                writeData36 = {17'b0, writeData[21]};
                writeData35 = {17'b0, writeData[20]};
                writeData34 = {17'b0, writeData[19]};
                writeData33 = {17'b0, writeData[18]};
                writeData32 = {17'b0, writeData[17]};
                writeData31 = {17'b0, writeData[16]};
                writeData30 = {17'b0, writeData[15]};
                writeData29 = {17'b0, writeData[14]};
                writeData28 = {17'b0, writeData[13]};
                writeData27 = {17'b0, writeData[12]};
                writeData26 = {17'b0, writeData[11]};
                writeData25 = {17'b0, writeData[10]};
                writeData24 = {17'b0, writeData[9]};
                writeData23 = {17'b0, writeData[8]};
                writeData22 = {17'b0, writeData[7]};
                writeData21 = {17'b0, writeData[6]};
                writeData20 = {17'b0, writeData[5]};
                writeData19 = {17'b0, writeData[4]};
                writeData18 = {17'b0, writeData[3]};
                writeData17 = {17'b0, writeData[2]};
                writeData16 = {17'b0, writeData[1]};
                writeData15 = {17'b0, writeData[0]};
                writeData14 = {14'b0, writeData[31:28]};
                writeData13 = {14'b0, writeData[27:24]};
                writeData12 = {14'b0, writeData[23:20]};
                writeData11 = {14'b0, writeData[19:16]};
                writeData10 = {14'b0, writeData[15:12]};
                writeData9 = {14'b0, writeData[11:8]};
                writeData8 = {14'b0, writeData[7:4]};
                writeData7 = {14'b0, writeData[3:0]};
                writeData6 = {10'b0, writeData[31:24]};
                writeData5 = {10'b0, writeData[23:16]};
                writeData4 = {10'b0, writeData[15:8]};
                writeData3 = {10'b0, writeData[7:0]};
                writeData2 = {1'b0, writeData[31:24], 1'b0, writeData[23:16]};
                writeData1 = {1'b0, writeData[15:8], 1'b0, writeData[7:0]};

                case (writeAddr[14:9])
                    6'b000000, 6'b000001, 6'b000010, 6'b000011,
                    6'b000100, 6'b000101, 6'b000110, 6'b000111,
                    6'b001000, 6'b001001, 6'b001010, 6'b001011,
                    6'b001100, 6'b001101, 6'b001110, 6'b001111,
                    6'b010000, 6'b010001, 6'b010010, 6'b010011,
                    6'b010100, 6'b010101, 6'b010110, 6'b010111,
                    6'b011000, 6'b011001, 6'b011010, 6'b011011,
                    6'b011100, 6'b011101, 6'b011110, 6'b011111 : begin
                        wen_a46 = {1'b0, wen};
                        wen_a45 = {1'b0, wen};
                        wen_a44 = {1'b0, wen};
                        wen_a43 = {1'b0, wen};
                        wen_a42 = {1'b0, wen};
                        wen_a41 = {1'b0, wen};
                        wen_a40 = {1'b0, wen};
                        wen_a39 = {1'b0, wen};
                        wen_a38 = {1'b0, wen};
                        wen_a37 = {1'b0, wen};
                        wen_a36 = {1'b0, wen};
                        wen_a35 = {1'b0, wen};
                        wen_a34 = {1'b0, wen};
                        wen_a33 = {1'b0, wen};
                        wen_a32 = {1'b0, wen};
                        wen_a31 = {1'b0, wen};
                        wen_a30 = {1'b0, wen};
                        wen_a29 = {1'b0, wen};
                        wen_a28 = {1'b0, wen};
                        wen_a27 = {1'b0, wen};
                        wen_a26 = {1'b0, wen};
                        wen_a25 = {1'b0, wen};
                        wen_a24 = {1'b0, wen};
                        wen_a23 = {1'b0, wen};
                        wen_a22 = {1'b0, wen};
                        wen_a21 = {1'b0, wen};
                        wen_a20 = {1'b0, wen};
                        wen_a19 = {1'b0, wen};
                        wen_a18 = {1'b0, wen};
                        wen_a17 = {1'b0, wen};
                        wen_a16 = {1'b0, wen};
                        wen_a15 = {1'b0, wen};
                        wen_a14 = {1'b0, 1'b0};
                        wen_a13 = {1'b0, 1'b0};
                        wen_a12 = {1'b0, 1'b0};
                        wen_a11 = {1'b0, 1'b0};
                        wen_a10 = {1'b0, 1'b0};
                        wen_a9 = {1'b0, 1'b0};
                        wen_a8 = {1'b0, 1'b0};
                        wen_a7 = {1'b0, 1'b0};
                        wen_a6 = {1'b0, 1'b0};
                        wen_a5 = {1'b0, 1'b0};
                        wen_a4 = {1'b0, 1'b0};
                        wen_a3 = {1'b0, 1'b0};
                        wen_a2 = {1'b0, 1'b0};
                        wen_a1 = {1'b0, 1'b0};
                    end
                    6'b100000, 6'b100001, 6'b100010, 6'b100011,
                    6'b100100, 6'b100101, 6'b100110, 6'b100111: begin
                        wen_a46 = {1'b0, 1'b0};
                        wen_a45 = {1'b0, 1'b0};
                        wen_a44 = {1'b0, 1'b0};
                        wen_a43 = {1'b0, 1'b0};
                        wen_a42 = {1'b0, 1'b0};
                        wen_a41 = {1'b0, 1'b0};
                        wen_a40 = {1'b0, 1'b0};
                        wen_a39 = {1'b0, 1'b0};
                        wen_a38 = {1'b0, 1'b0};
                        wen_a37 = {1'b0, 1'b0};
                        wen_a36 = {1'b0, 1'b0};
                        wen_a35 = {1'b0, 1'b0};
                        wen_a34 = {1'b0, 1'b0};
                        wen_a33 = {1'b0, 1'b0};
                        wen_a32 = {1'b0, 1'b0};
                        wen_a31 = {1'b0, 1'b0};
                        wen_a30 = {1'b0, 1'b0};
                        wen_a29 = {1'b0, 1'b0};
                        wen_a28 = {1'b0, 1'b0};
                        wen_a27 = {1'b0, 1'b0};
                        wen_a26 = {1'b0, 1'b0};
                        wen_a25 = {1'b0, 1'b0};
                        wen_a24 = {1'b0, 1'b0};
                        wen_a23 = {1'b0, 1'b0};
                        wen_a22 = {1'b0, 1'b0};
                        wen_a21 = {1'b0, 1'b0};
                        wen_a20 = {1'b0, 1'b0};
                        wen_a19 = {1'b0, 1'b0};
                        wen_a18 = {1'b0, 1'b0};
                        wen_a17 = {1'b0, 1'b0};
                        wen_a16 = {1'b0, 1'b0};
                        wen_a15 = {1'b0, 1'b0};
                        wen_a14 = {1'b0, wen};
                        wen_a13 = {1'b0, wen};
                        wen_a12 = {1'b0, wen};
                        wen_a11 = {1'b0, wen};
                        wen_a10 = {1'b0, wen};
                        wen_a9 = {1'b0, wen};
                        wen_a8 = {1'b0, wen};
                        wen_a7 = {1'b0, wen};
                        wen_a6 = {1'b0, 1'b0};
                        wen_a5 = {1'b0, 1'b0};
                        wen_a4 = {1'b0, 1'b0};
                        wen_a3 = {1'b0, 1'b0};
                        wen_a2 = {1'b0, 1'b0};
                        wen_a1 = {1'b0, 1'b0};
                    end
                    6'b101000, 6'b101001, 6'b101010, 6'b101011 : begin
                        wen_a46 = {1'b0, 1'b0};
                        wen_a45 = {1'b0, 1'b0};
                        wen_a44 = {1'b0, 1'b0};
                        wen_a43 = {1'b0, 1'b0};
                        wen_a42 = {1'b0, 1'b0};
                        wen_a41 = {1'b0, 1'b0};
                        wen_a40 = {1'b0, 1'b0};
                        wen_a39 = {1'b0, 1'b0};
                        wen_a38 = {1'b0, 1'b0};
                        wen_a37 = {1'b0, 1'b0};
                        wen_a36 = {1'b0, 1'b0};
                        wen_a35 = {1'b0, 1'b0};
                        wen_a34 = {1'b0, 1'b0};
                        wen_a33 = {1'b0, 1'b0};
                        wen_a32 = {1'b0, 1'b0};
                        wen_a31 = {1'b0, 1'b0};
                        wen_a30 = {1'b0, 1'b0};
                        wen_a29 = {1'b0, 1'b0};
                        wen_a28 = {1'b0, 1'b0};
                        wen_a27 = {1'b0, 1'b0};
                        wen_a26 = {1'b0, 1'b0};
                        wen_a25 = {1'b0, 1'b0};
                        wen_a24 = {1'b0, 1'b0};
                        wen_a23 = {1'b0, 1'b0};
                        wen_a22 = {1'b0, 1'b0};
                        wen_a21 = {1'b0, 1'b0};
                        wen_a20 = {1'b0, 1'b0};
                        wen_a19 = {1'b0, 1'b0};
                        wen_a18 = {1'b0, 1'b0};
                        wen_a17 = {1'b0, 1'b0};
                        wen_a16 = {1'b0, 1'b0};
                        wen_a15 = {1'b0, 1'b0};
                        wen_a14 = {1'b0, 1'b0};
                        wen_a13 = {1'b0, 1'b0};
                        wen_a12 = {1'b0, 1'b0};
                        wen_a11 = {1'b0, 1'b0};
                        wen_a10 = {1'b0, 1'b0};
                        wen_a9 = {1'b0, 1'b0};
                        wen_a8 = {1'b0, 1'b0};
                        wen_a7 = {1'b0, 1'b0};
                        wen_a6 = {1'b0, wen};
                        wen_a5 = {1'b0, wen};
                        wen_a4 = {1'b0, wen};
                        wen_a3 = {1'b0, wen};
                        wen_a2 = {1'b0, 1'b0};
                        wen_a1 = {1'b0, 1'b0};
                    end
                    6'b101100, 6'b101101 : begin
                        wen_a46 = {1'b0, 1'b0};
                        wen_a45 = {1'b0, 1'b0};
                        wen_a44 = {1'b0, 1'b0};
                        wen_a43 = {1'b0, 1'b0};
                        wen_a42 = {1'b0, 1'b0};
                        wen_a41 = {1'b0, 1'b0};
                        wen_a40 = {1'b0, 1'b0};
                        wen_a39 = {1'b0, 1'b0};
                        wen_a38 = {1'b0, 1'b0};
                        wen_a37 = {1'b0, 1'b0};
                        wen_a36 = {1'b0, 1'b0};
                        wen_a35 = {1'b0, 1'b0};
                        wen_a34 = {1'b0, 1'b0};
                        wen_a33 = {1'b0, 1'b0};
                        wen_a32 = {1'b0, 1'b0};
                        wen_a31 = {1'b0, 1'b0};
                        wen_a30 = {1'b0, 1'b0};
                        wen_a29 = {1'b0, 1'b0};
                        wen_a28 = {1'b0, 1'b0};
                        wen_a27 = {1'b0, 1'b0};
                        wen_a26 = {1'b0, 1'b0};
                        wen_a25 = {1'b0, 1'b0};
                        wen_a24 = {1'b0, 1'b0};
                        wen_a23 = {1'b0, 1'b0};
                        wen_a22 = {1'b0, 1'b0};
                        wen_a21 = {1'b0, 1'b0};
                        wen_a20 = {1'b0, 1'b0};
                        wen_a19 = {1'b0, 1'b0};
                        wen_a18 = {1'b0, 1'b0};
                        wen_a17 = {1'b0, 1'b0};
                        wen_a16 = {1'b0, 1'b0};
                        wen_a15 = {1'b0, 1'b0};
                        wen_a14 = {1'b0, 1'b0};
                        wen_a13 = {1'b0, 1'b0};
                        wen_a12 = {1'b0, 1'b0};
                        wen_a11 = {1'b0, 1'b0};
                        wen_a10 = {1'b0, 1'b0};
                        wen_a9 = {1'b0, 1'b0};
                        wen_a8 = {1'b0, 1'b0};
                        wen_a7 = {1'b0, 1'b0};
                        wen_a6 = {1'b0, 1'b0};
                        wen_a5 = {1'b0, 1'b0};
                        wen_a4 = {1'b0, 1'b0};
                        wen_a3 = {1'b0, 1'b0};
                        wen_a2 = {wen, wen};
                        wen_a1 = {wen, wen};
                    end
                    default : begin
                        wen_a46 = {1'b0, 1'b0};
                        wen_a45 = {1'b0, 1'b0};
                        wen_a44 = {1'b0, 1'b0};
                        wen_a43 = {1'b0, 1'b0};
                        wen_a42 = {1'b0, 1'b0};
                        wen_a41 = {1'b0, 1'b0};
                        wen_a40 = {1'b0, 1'b0};
                        wen_a39 = {1'b0, 1'b0};
                        wen_a38 = {1'b0, 1'b0};
                        wen_a37 = {1'b0, 1'b0};
                        wen_a36 = {1'b0, 1'b0};
                        wen_a35 = {1'b0, 1'b0};
                        wen_a34 = {1'b0, 1'b0};
                        wen_a33 = {1'b0, 1'b0};
                        wen_a32 = {1'b0, 1'b0};
                        wen_a31 = {1'b0, 1'b0};
                        wen_a30 = {1'b0, 1'b0};
                        wen_a29 = {1'b0, 1'b0};
                        wen_a28 = {1'b0, 1'b0};
                        wen_a27 = {1'b0, 1'b0};
                        wen_a26 = {1'b0, 1'b0};
                        wen_a25 = {1'b0, 1'b0};
                        wen_a24 = {1'b0, 1'b0};
                        wen_a23 = {1'b0, 1'b0};
                        wen_a22 = {1'b0, 1'b0};
                        wen_a21 = {1'b0, 1'b0};
                        wen_a20 = {1'b0, 1'b0};
                        wen_a19 = {1'b0, 1'b0};
                        wen_a18 = {1'b0, 1'b0};
                        wen_a17 = {1'b0, 1'b0};
                        wen_a16 = {1'b0, 1'b0};
                        wen_a15 = {1'b0, 1'b0};
                        wen_a14 = {1'b0, 1'b0};
                        wen_a13 = {1'b0, 1'b0};
                        wen_a12 = {1'b0, 1'b0};
                        wen_a11 = {1'b0, 1'b0};
                        wen_a10 = {1'b0, 1'b0};
                        wen_a9 = {1'b0, 1'b0};
                        wen_a8 = {1'b0, 1'b0};
                        wen_a7 = {1'b0, 1'b0};
                        wen_a6 = {1'b0, 1'b0};
                        wen_a5 = {1'b0, 1'b0};
                        wen_a4 = {1'b0, 1'b0};
                        wen_a3 = {1'b0, 1'b0};
                        wen_a2 = {1'b0, 1'b0};
                        wen_a1 = {1'b0, 1'b0};
                    end
                endcase

                case (ckRdAddr[14:9])
                    6'b000000, 6'b000001, 6'b000010, 6'b000011,
                    6'b000100, 6'b000101, 6'b000110, 6'b000111,
                    6'b001000, 6'b001001, 6'b001010, 6'b001011,
                    6'b001100, 6'b001101, 6'b001110, 6'b001111,
                    6'b010000, 6'b010001, 6'b010010, 6'b010011,
                    6'b010100, 6'b010101, 6'b010110, 6'b010111,
                    6'b011000, 6'b011001, 6'b011010, 6'b011011,
                    6'b011100, 6'b011101, 6'b011110, 6'b011111 : begin
                        readData = {
                                        readData46[0],
                                        readData45[0],
                                        readData44[0],
                                        readData43[0],
                                        readData42[0],
                                        readData41[0],
                                        readData40[0],
                                        readData39[0],
                                        readData38[0],
                                        readData37[0],
                                        readData36[0],
                                        readData35[0],
                                        readData34[0],
                                        readData33[0],
                                        readData32[0],
                                        readData31[0],
                                        readData30[0],
                                        readData29[0],
                                        readData28[0],
                                        readData27[0],
                                        readData26[0],
                                        readData25[0],
                                        readData24[0],
                                        readData23[0],
                                        readData22[0],
                                        readData21[0],
                                        readData20[0],
                                        readData19[0],
                                        readData18[0],
                                        readData17[0],
                                        readData16[0],
                                        readData15[0]
                        };
                    end
                    6'b100000, 6'b100001, 6'b100010, 6'b100011,
                    6'b100100, 6'b100101, 6'b100110, 6'b100111: begin
                        readData = {
                                        readData14[3:0],
                                        readData13[3:0],
                                        readData12[3:0],
                                        readData11[3:0],
                                        readData10[3:0],
                                        readData9[3:0],
                                        readData8[3:0],
                                        readData7[3:0]
                        };
                    end
                    6'b101000, 6'b101001, 6'b101010, 6'b101011: begin
                        readData = {readData6[7:0],readData5[7:0],readData4[7:0],readData3[7:0]};
                    end
                    6'b101100, 6'b101101 : begin
                        readData = {readData2[16:9],readData2[7:0],readData1[16:9],readData1[7:0]};
                    end
                    default : begin
                        readData = 32'b0;
                    end
                endcase
            end        
            24064: begin
                width46 = 3'b000;
                width45 = 3'b000;
                width44 = 3'b000;
                width43 = 3'b000;
                width42 = 3'b000;
                width41 = 3'b000;
                width40 = 3'b000;
                width39 = 3'b000;
                width38 = 3'b000;
                width37 = 3'b000;
                width36 = 3'b000;
                width35 = 3'b000;
                width34 = 3'b000;
                width33 = 3'b000;
                width32 = 3'b000;
                width31 = 3'b000;
                width30 = 3'b000;
                width29 = 3'b000;
                width28 = 3'b000;
                width27 = 3'b000;
                width26 = 3'b000;
                width25 = 3'b000;
                width24 = 3'b000;
                width23 = 3'b000;
                width22 = 3'b000;
                width21 = 3'b000;
                width20 = 3'b000;
                width19 = 3'b000;
                width18 = 3'b000;
                width17 = 3'b000;
                width16 = 3'b000;
                width15 = 3'b000;
                width14 = 3'b010;
                width13 = 3'b010;
                width12 = 3'b010;
                width11 = 3'b010;
                width10 = 3'b010;
                width9 = 3'b010;
                width8 = 3'b010;
                width7 = 3'b010;
                width6 = 3'b011;
                width5 = 3'b011;
                width4 = 3'b011;
                width3 = 3'b011;
                width2 = 3'b100;
                width1 = 3'b100;
                width0 = 3'b101;

                writeAddr46 = {writeAddr[13:0]};
                writeAddr45 = {writeAddr[13:0]};
                writeAddr44 = {writeAddr[13:0]};
                writeAddr43 = {writeAddr[13:0]};
                writeAddr42 = {writeAddr[13:0]};
                writeAddr41 = {writeAddr[13:0]};
                writeAddr40 = {writeAddr[13:0]};
                writeAddr39 = {writeAddr[13:0]};
                writeAddr38 = {writeAddr[13:0]};
                writeAddr37 = {writeAddr[13:0]};
                writeAddr36 = {writeAddr[13:0]};
                writeAddr35 = {writeAddr[13:0]};
                writeAddr34 = {writeAddr[13:0]};
                writeAddr33 = {writeAddr[13:0]};
                writeAddr32 = {writeAddr[13:0]};
                writeAddr31 = {writeAddr[13:0]};
                writeAddr30 = {writeAddr[13:0]};
                writeAddr29 = {writeAddr[13:0]};
                writeAddr28 = {writeAddr[13:0]};
                writeAddr27 = {writeAddr[13:0]};
                writeAddr26 = {writeAddr[13:0]};
                writeAddr25 = {writeAddr[13:0]};
                writeAddr24 = {writeAddr[13:0]};
                writeAddr23 = {writeAddr[13:0]};
                writeAddr22 = {writeAddr[13:0]};
                writeAddr21 = {writeAddr[13:0]};
                writeAddr20 = {writeAddr[13:0]};
                writeAddr19 = {writeAddr[13:0]};
                writeAddr18 = {writeAddr[13:0]};
                writeAddr17 = {writeAddr[13:0]};
                writeAddr16 = {writeAddr[13:0]};
                writeAddr15 = {writeAddr[13:0]};
                writeAddr14 = {writeAddr[11:0], 2'b0};
                writeAddr13 = {writeAddr[11:0], 2'b0};
                writeAddr12 = {writeAddr[11:0], 2'b0};
                writeAddr11 = {writeAddr[11:0], 2'b0};
                writeAddr10 = {writeAddr[11:0], 2'b0};
                writeAddr9 = {writeAddr[11:0], 2'b0};
                writeAddr8 = {writeAddr[11:0], 2'b0};
                writeAddr7 = {writeAddr[11:0], 2'b0};
                writeAddr6 = {writeAddr[10:0], 3'b0};
                writeAddr5 = {writeAddr[10:0], 3'b0};
                writeAddr4 = {writeAddr[10:0], 3'b0};
                writeAddr3 = {writeAddr[10:0], 3'b0};
                writeAddr2 = {writeAddr[9:0], 4'b0};
                writeAddr1 = {writeAddr[9:0], 4'b0};
                writeAddr0 = {writeAddr[8:0], 5'b0};

                readAddr46 = {writeAddr[13:0]};
                readAddr45 = {writeAddr[13:0]};
                readAddr44 = {writeAddr[13:0]};
                readAddr43 = {writeAddr[13:0]};
                readAddr42 = {writeAddr[13:0]};
                readAddr41 = {writeAddr[13:0]};
                readAddr40 = {writeAddr[13:0]};
                readAddr39 = {writeAddr[13:0]};
                readAddr38 = {writeAddr[13:0]};
                readAddr37 = {writeAddr[13:0]};
                readAddr36 = {writeAddr[13:0]};
                readAddr35 = {writeAddr[13:0]};
                readAddr34 = {writeAddr[13:0]};
                readAddr33 = {writeAddr[13:0]};
                readAddr32 = {writeAddr[13:0]};
                readAddr31 = {writeAddr[13:0]};
                readAddr30 = {writeAddr[13:0]};
                readAddr29 = {writeAddr[13:0]};
                readAddr28 = {writeAddr[13:0]};
                readAddr27 = {writeAddr[13:0]};
                readAddr26 = {writeAddr[13:0]};
                readAddr25 = {writeAddr[13:0]};
                readAddr24 = {writeAddr[13:0]};
                readAddr23 = {writeAddr[13:0]};
                readAddr22 = {writeAddr[13:0]};
                readAddr21 = {writeAddr[13:0]};
                readAddr20 = {writeAddr[13:0]};
                readAddr19 = {writeAddr[13:0]};
                readAddr18 = {writeAddr[13:0]};
                readAddr17 = {writeAddr[13:0]};
                readAddr16 = {writeAddr[13:0]};
                readAddr15 = {writeAddr[13:0]};
                readAddr14  = {readAddr[11:0],  2'b0};
                readAddr13  = {readAddr[11:0],  2'b0};
                readAddr12  = {readAddr[11:0],  2'b0};
                readAddr11  = {readAddr[11:0],  2'b0};
                readAddr10  = {readAddr[11:0],  2'b0};
                readAddr9  = {readAddr[11:0],  2'b0};
                readAddr8  = {readAddr[11:0],  2'b0};
                readAddr7  = {readAddr[11:0],  2'b0};
                readAddr6  = {readAddr[10:0],  3'b0};
                readAddr5  = {readAddr[10:0],  3'b0};
                readAddr4  = {readAddr[10:0],  3'b0};
                readAddr3  = {readAddr[10:0],  3'b0};
                readAddr2  = {readAddr[9:0],  4'b0};
                readAddr1  = {readAddr[9:0],  4'b0};
                readAddr0  = {readAddr[8:0],  5'b0};

                writeData46 = {17'b0, writeData[31]};
                writeData45 = {17'b0, writeData[30]};
                writeData44 = {17'b0, writeData[29]};
                writeData43 = {17'b0, writeData[28]};
                writeData42 = {17'b0, writeData[27]};
                writeData41 = {17'b0, writeData[26]};
                writeData40 = {17'b0, writeData[25]};
                writeData39 = {17'b0, writeData[24]};
                writeData38 = {17'b0, writeData[23]};
                writeData37 = {17'b0, writeData[22]};
                writeData36 = {17'b0, writeData[21]};
                writeData35 = {17'b0, writeData[20]};
                writeData34 = {17'b0, writeData[19]};
                writeData33 = {17'b0, writeData[18]};
                writeData32 = {17'b0, writeData[17]};
                writeData31 = {17'b0, writeData[16]};
                writeData30 = {17'b0, writeData[15]};
                writeData29 = {17'b0, writeData[14]};
                writeData28 = {17'b0, writeData[13]};
                writeData27 = {17'b0, writeData[12]};
                writeData26 = {17'b0, writeData[11]};
                writeData25 = {17'b0, writeData[10]};
                writeData24 = {17'b0, writeData[9]};
                writeData23 = {17'b0, writeData[8]};
                writeData22 = {17'b0, writeData[7]};
                writeData21 = {17'b0, writeData[6]};
                writeData20 = {17'b0, writeData[5]};
                writeData19 = {17'b0, writeData[4]};
                writeData18 = {17'b0, writeData[3]};
                writeData17 = {17'b0, writeData[2]};
                writeData16 = {17'b0, writeData[1]};
                writeData15 = {17'b0, writeData[0]};
                writeData14 = {14'b0, writeData[31:28]};
                writeData13 = {14'b0, writeData[27:24]};
                writeData12 = {14'b0, writeData[23:20]};
                writeData11 = {14'b0, writeData[19:16]};
                writeData10 = {14'b0, writeData[15:12]};
                writeData9 = {14'b0, writeData[11:8]};
                writeData8 = {14'b0, writeData[7:4]};
                writeData7 = {14'b0, writeData[3:0]};
                writeData6 = {10'b0, writeData[31:24]};
                writeData5 = {10'b0, writeData[23:16]};
                writeData4 = {10'b0, writeData[15:8]};
                writeData3 = {10'b0, writeData[7:0]};
                writeData2 = {1'b0, writeData[31:24], 1'b0, writeData[23:16]};
                writeData1 = {1'b0, writeData[15:8], 1'b0, writeData[7:0]};
                writeData0 = {1'b0, writeData[31:24], 1'b0, writeData[23:16], 1'b0, writeData[15:8], 1'b0, writeData[7:0]};

                case (writeAddr[14:9])
                    6'b000000, 6'b000001, 6'b000010, 6'b000011,
                    6'b000100, 6'b000101, 6'b000110, 6'b000111,
                    6'b001000, 6'b001001, 6'b001010, 6'b001011,
                    6'b001100, 6'b001101, 6'b001110, 6'b001111,
                    6'b010000, 6'b010001, 6'b010010, 6'b010011,
                    6'b010100, 6'b010101, 6'b010110, 6'b010111,
                    6'b011000, 6'b011001, 6'b011010, 6'b011011,
                    6'b011100, 6'b011101, 6'b011110, 6'b011111 : begin
                        wen_a46 = {1'b0, wen};
                        wen_a45 = {1'b0, wen};
                        wen_a44 = {1'b0, wen};
                        wen_a43 = {1'b0, wen};
                        wen_a42 = {1'b0, wen};
                        wen_a41 = {1'b0, wen};
                        wen_a40 = {1'b0, wen};
                        wen_a39 = {1'b0, wen};
                        wen_a38 = {1'b0, wen};
                        wen_a37 = {1'b0, wen};
                        wen_a36 = {1'b0, wen};
                        wen_a35 = {1'b0, wen};
                        wen_a34 = {1'b0, wen};
                        wen_a33 = {1'b0, wen};
                        wen_a32 = {1'b0, wen};
                        wen_a31 = {1'b0, wen};
                        wen_a30 = {1'b0, wen};
                        wen_a29 = {1'b0, wen};
                        wen_a28 = {1'b0, wen};
                        wen_a27 = {1'b0, wen};
                        wen_a26 = {1'b0, wen};
                        wen_a25 = {1'b0, wen};
                        wen_a24 = {1'b0, wen};
                        wen_a23 = {1'b0, wen};
                        wen_a22 = {1'b0, wen};
                        wen_a21 = {1'b0, wen};
                        wen_a20 = {1'b0, wen};
                        wen_a19 = {1'b0, wen};
                        wen_a18 = {1'b0, wen};
                        wen_a17 = {1'b0, wen};
                        wen_a16 = {1'b0, wen};
                        wen_a15 = {1'b0, wen};
                        wen_a14 = {1'b0, 1'b0};
                        wen_a13 = {1'b0, 1'b0};
                        wen_a12 = {1'b0, 1'b0};
                        wen_a11 = {1'b0, 1'b0};
                        wen_a10 = {1'b0, 1'b0};
                        wen_a9 = {1'b0, 1'b0};
                        wen_a8 = {1'b0, 1'b0};
                        wen_a7 = {1'b0, 1'b0};
                        wen_a6 = {1'b0, 1'b0};
                        wen_a5 = {1'b0, 1'b0};
                        wen_a4 = {1'b0, 1'b0};
                        wen_a3 = {1'b0, 1'b0};
                        wen_a2 = {1'b0, 1'b0};
                        wen_a1 = {1'b0, 1'b0};
                        wen_a0 = {1'b0, 1'b0};
                        wen_b0 = {1'b0, 1'b0};
                    end
                    6'b100000, 6'b100001, 6'b100010, 6'b100011,
                    6'b100100, 6'b100101, 6'b100110, 6'b100111: begin
                        wen_a46 = {1'b0, 1'b0};
                        wen_a45 = {1'b0, 1'b0};
                        wen_a44 = {1'b0, 1'b0};
                        wen_a43 = {1'b0, 1'b0};
                        wen_a42 = {1'b0, 1'b0};
                        wen_a41 = {1'b0, 1'b0};
                        wen_a40 = {1'b0, 1'b0};
                        wen_a39 = {1'b0, 1'b0};
                        wen_a38 = {1'b0, 1'b0};
                        wen_a37 = {1'b0, 1'b0};
                        wen_a36 = {1'b0, 1'b0};
                        wen_a35 = {1'b0, 1'b0};
                        wen_a34 = {1'b0, 1'b0};
                        wen_a33 = {1'b0, 1'b0};
                        wen_a32 = {1'b0, 1'b0};
                        wen_a31 = {1'b0, 1'b0};
                        wen_a30 = {1'b0, 1'b0};
                        wen_a29 = {1'b0, 1'b0};
                        wen_a28 = {1'b0, 1'b0};
                        wen_a27 = {1'b0, 1'b0};
                        wen_a26 = {1'b0, 1'b0};
                        wen_a25 = {1'b0, 1'b0};
                        wen_a24 = {1'b0, 1'b0};
                        wen_a23 = {1'b0, 1'b0};
                        wen_a22 = {1'b0, 1'b0};
                        wen_a21 = {1'b0, 1'b0};
                        wen_a20 = {1'b0, 1'b0};
                        wen_a19 = {1'b0, 1'b0};
                        wen_a18 = {1'b0, 1'b0};
                        wen_a17 = {1'b0, 1'b0};
                        wen_a16 = {1'b0, 1'b0};
                        wen_a15 = {1'b0, 1'b0};
                        wen_a14 = {1'b0, wen};
                        wen_a13 = {1'b0, wen};
                        wen_a12 = {1'b0, wen};
                        wen_a11 = {1'b0, wen};
                        wen_a10 = {1'b0, wen};
                        wen_a9 = {1'b0, wen};
                        wen_a8 = {1'b0, wen};
                        wen_a7 = {1'b0, wen};
                        wen_a6 = {1'b0, 1'b0};
                        wen_a5 = {1'b0, 1'b0};
                        wen_a4 = {1'b0, 1'b0};
                        wen_a3 = {1'b0, 1'b0};
                        wen_a2 = {1'b0, 1'b0};
                        wen_a1 = {1'b0, 1'b0};
                        wen_a0 = {1'b0, 1'b0};
                        wen_b0 = {1'b0, 1'b0};
                    end
                    6'b101000, 6'b101001, 6'b101010, 6'b101011 : begin
                        wen_a46 = {1'b0, 1'b0};
                        wen_a45 = {1'b0, 1'b0};
                        wen_a44 = {1'b0, 1'b0};
                        wen_a43 = {1'b0, 1'b0};
                        wen_a42 = {1'b0, 1'b0};
                        wen_a41 = {1'b0, 1'b0};
                        wen_a40 = {1'b0, 1'b0};
                        wen_a39 = {1'b0, 1'b0};
                        wen_a38 = {1'b0, 1'b0};
                        wen_a37 = {1'b0, 1'b0};
                        wen_a36 = {1'b0, 1'b0};
                        wen_a35 = {1'b0, 1'b0};
                        wen_a34 = {1'b0, 1'b0};
                        wen_a33 = {1'b0, 1'b0};
                        wen_a32 = {1'b0, 1'b0};
                        wen_a31 = {1'b0, 1'b0};
                        wen_a30 = {1'b0, 1'b0};
                        wen_a29 = {1'b0, 1'b0};
                        wen_a28 = {1'b0, 1'b0};
                        wen_a27 = {1'b0, 1'b0};
                        wen_a26 = {1'b0, 1'b0};
                        wen_a25 = {1'b0, 1'b0};
                        wen_a24 = {1'b0, 1'b0};
                        wen_a23 = {1'b0, 1'b0};
                        wen_a22 = {1'b0, 1'b0};
                        wen_a21 = {1'b0, 1'b0};
                        wen_a20 = {1'b0, 1'b0};
                        wen_a19 = {1'b0, 1'b0};
                        wen_a18 = {1'b0, 1'b0};
                        wen_a17 = {1'b0, 1'b0};
                        wen_a16 = {1'b0, 1'b0};
                        wen_a15 = {1'b0, 1'b0};
                        wen_a14 = {1'b0, 1'b0};
                        wen_a13 = {1'b0, 1'b0};
                        wen_a12 = {1'b0, 1'b0};
                        wen_a11 = {1'b0, 1'b0};
                        wen_a10 = {1'b0, 1'b0};
                        wen_a9 = {1'b0, 1'b0};
                        wen_a8 = {1'b0, 1'b0};
                        wen_a7 = {1'b0, 1'b0};
                        wen_a6 = {1'b0, wen};
                        wen_a5 = {1'b0, wen};
                        wen_a4 = {1'b0, wen};
                        wen_a3 = {1'b0, wen};
                        wen_a2 = {1'b0, 1'b0};
                        wen_a1 = {1'b0, 1'b0};
                        wen_a0 = {1'b0, 1'b0};
                        wen_b0 = {1'b0, 1'b0};
                    end
                    6'b101100, 6'b101101 : begin
                        wen_a46 = {1'b0, 1'b0};
                        wen_a45 = {1'b0, 1'b0};
                        wen_a44 = {1'b0, 1'b0};
                        wen_a43 = {1'b0, 1'b0};
                        wen_a42 = {1'b0, 1'b0};
                        wen_a41 = {1'b0, 1'b0};
                        wen_a40 = {1'b0, 1'b0};
                        wen_a39 = {1'b0, 1'b0};
                        wen_a38 = {1'b0, 1'b0};
                        wen_a37 = {1'b0, 1'b0};
                        wen_a36 = {1'b0, 1'b0};
                        wen_a35 = {1'b0, 1'b0};
                        wen_a34 = {1'b0, 1'b0};
                        wen_a33 = {1'b0, 1'b0};
                        wen_a32 = {1'b0, 1'b0};
                        wen_a31 = {1'b0, 1'b0};
                        wen_a30 = {1'b0, 1'b0};
                        wen_a29 = {1'b0, 1'b0};
                        wen_a28 = {1'b0, 1'b0};
                        wen_a27 = {1'b0, 1'b0};
                        wen_a26 = {1'b0, 1'b0};
                        wen_a25 = {1'b0, 1'b0};
                        wen_a24 = {1'b0, 1'b0};
                        wen_a23 = {1'b0, 1'b0};
                        wen_a22 = {1'b0, 1'b0};
                        wen_a21 = {1'b0, 1'b0};
                        wen_a20 = {1'b0, 1'b0};
                        wen_a19 = {1'b0, 1'b0};
                        wen_a18 = {1'b0, 1'b0};
                        wen_a17 = {1'b0, 1'b0};
                        wen_a16 = {1'b0, 1'b0};
                        wen_a15 = {1'b0, 1'b0};
                        wen_a14 = {1'b0, 1'b0};
                        wen_a13 = {1'b0, 1'b0};
                        wen_a12 = {1'b0, 1'b0};
                        wen_a11 = {1'b0, 1'b0};
                        wen_a10 = {1'b0, 1'b0};
                        wen_a9 = {1'b0, 1'b0};
                        wen_a8 = {1'b0, 1'b0};
                        wen_a7 = {1'b0, 1'b0};
                        wen_a6 = {1'b0, 1'b0};
                        wen_a5 = {1'b0, 1'b0};
                        wen_a4 = {1'b0, 1'b0};
                        wen_a3 = {1'b0, 1'b0};
                        wen_a2 = {wen, wen};
                        wen_a1 = {wen, wen};
                        wen_a0 = {1'b0, 1'b0};
                        wen_b0 = {1'b0, 1'b0};
                    end
                    6'b101110 : begin
                        wen_a46 = {1'b0, 1'b0};
                        wen_a45 = {1'b0, 1'b0};
                        wen_a44 = {1'b0, 1'b0};
                        wen_a43 = {1'b0, 1'b0};
                        wen_a42 = {1'b0, 1'b0};
                        wen_a41 = {1'b0, 1'b0};
                        wen_a40 = {1'b0, 1'b0};
                        wen_a39 = {1'b0, 1'b0};
                        wen_a38 = {1'b0, 1'b0};
                        wen_a37 = {1'b0, 1'b0};
                        wen_a36 = {1'b0, 1'b0};
                        wen_a35 = {1'b0, 1'b0};
                        wen_a34 = {1'b0, 1'b0};
                        wen_a33 = {1'b0, 1'b0};
                        wen_a32 = {1'b0, 1'b0};
                        wen_a31 = {1'b0, 1'b0};
                        wen_a30 = {1'b0, 1'b0};
                        wen_a29 = {1'b0, 1'b0};
                        wen_a28 = {1'b0, 1'b0};
                        wen_a27 = {1'b0, 1'b0};
                        wen_a26 = {1'b0, 1'b0};
                        wen_a25 = {1'b0, 1'b0};
                        wen_a24 = {1'b0, 1'b0};
                        wen_a23 = {1'b0, 1'b0};
                        wen_a22 = {1'b0, 1'b0};
                        wen_a21 = {1'b0, 1'b0};
                        wen_a20 = {1'b0, 1'b0};
                        wen_a19 = {1'b0, 1'b0};
                        wen_a18 = {1'b0, 1'b0};
                        wen_a17 = {1'b0, 1'b0};
                        wen_a16 = {1'b0, 1'b0};
                        wen_a15 = {1'b0, 1'b0};
                        wen_a14 = {1'b0, 1'b0};
                        wen_a13 = {1'b0, 1'b0};
                        wen_a12 = {1'b0, 1'b0};
                        wen_a11 = {1'b0, 1'b0};
                        wen_a10 = {1'b0, 1'b0};
                        wen_a9 = {1'b0, 1'b0};
                        wen_a8 = {1'b0, 1'b0};
                        wen_a7 = {1'b0, 1'b0};
                        wen_a6 = {1'b0, 1'b0};
                        wen_a5 = {1'b0, 1'b0};
                        wen_a4 = {1'b0, 1'b0};
                        wen_a3 = {1'b0, 1'b0};
                        wen_a2 = {1'b0, 1'b0};
                        wen_a1 = {1'b0, 1'b0};
                        wen_a0 = {wen, wen};
                        wen_b0 = {wen, wen};
                    end
                    default : begin
                        wen_a46 = {1'b0, 1'b0};
                        wen_a45 = {1'b0, 1'b0};
                        wen_a44 = {1'b0, 1'b0};
                        wen_a43 = {1'b0, 1'b0};
                        wen_a42 = {1'b0, 1'b0};
                        wen_a41 = {1'b0, 1'b0};
                        wen_a40 = {1'b0, 1'b0};
                        wen_a39 = {1'b0, 1'b0};
                        wen_a38 = {1'b0, 1'b0};
                        wen_a37 = {1'b0, 1'b0};
                        wen_a36 = {1'b0, 1'b0};
                        wen_a35 = {1'b0, 1'b0};
                        wen_a34 = {1'b0, 1'b0};
                        wen_a33 = {1'b0, 1'b0};
                        wen_a32 = {1'b0, 1'b0};
                        wen_a31 = {1'b0, 1'b0};
                        wen_a30 = {1'b0, 1'b0};
                        wen_a29 = {1'b0, 1'b0};
                        wen_a28 = {1'b0, 1'b0};
                        wen_a27 = {1'b0, 1'b0};
                        wen_a26 = {1'b0, 1'b0};
                        wen_a25 = {1'b0, 1'b0};
                        wen_a24 = {1'b0, 1'b0};
                        wen_a23 = {1'b0, 1'b0};
                        wen_a22 = {1'b0, 1'b0};
                        wen_a21 = {1'b0, 1'b0};
                        wen_a20 = {1'b0, 1'b0};
                        wen_a19 = {1'b0, 1'b0};
                        wen_a18 = {1'b0, 1'b0};
                        wen_a17 = {1'b0, 1'b0};
                        wen_a16 = {1'b0, 1'b0};
                        wen_a15 = {1'b0, 1'b0};
                        wen_a14 = {1'b0, 1'b0};
                        wen_a13 = {1'b0, 1'b0};
                        wen_a12 = {1'b0, 1'b0};
                        wen_a11 = {1'b0, 1'b0};
                        wen_a10 = {1'b0, 1'b0};
                        wen_a9 = {1'b0, 1'b0};
                        wen_a8 = {1'b0, 1'b0};
                        wen_a7 = {1'b0, 1'b0};
                        wen_a6 = {1'b0, 1'b0};
                        wen_a5 = {1'b0, 1'b0};
                        wen_a4 = {1'b0, 1'b0};
                        wen_a3 = {1'b0, 1'b0};
                        wen_a2 = {1'b0, 1'b0};
                        wen_a1 = {1'b0, 1'b0};
                        wen_a0 = {1'b0, 1'b0};
                        wen_b0 = {1'b0, 1'b0};
                    end
                endcase

                case (ckRdAddr[14:9])
                    6'b000000, 6'b000001, 6'b000010, 6'b000011,
                    6'b000100, 6'b000101, 6'b000110, 6'b000111,
                    6'b001000, 6'b001001, 6'b001010, 6'b001011,
                    6'b001100, 6'b001101, 6'b001110, 6'b001111,
                    6'b010000, 6'b010001, 6'b010010, 6'b010011,
                    6'b010100, 6'b010101, 6'b010110, 6'b010111,
                    6'b011000, 6'b011001, 6'b011010, 6'b011011,
                    6'b011100, 6'b011101, 6'b011110, 6'b011111 : begin
                        readData = {
                                        readData46[0],
                                        readData45[0],
                                        readData44[0],
                                        readData43[0],
                                        readData42[0],
                                        readData41[0],
                                        readData40[0],
                                        readData39[0],
                                        readData38[0],
                                        readData37[0],
                                        readData36[0],
                                        readData35[0],
                                        readData34[0],
                                        readData33[0],
                                        readData32[0],
                                        readData31[0],
                                        readData30[0],
                                        readData29[0],
                                        readData28[0],
                                        readData27[0],
                                        readData26[0],
                                        readData25[0],
                                        readData24[0],
                                        readData23[0],
                                        readData22[0],
                                        readData21[0],
                                        readData20[0],
                                        readData19[0],
                                        readData18[0],
                                        readData17[0],
                                        readData16[0],
                                        readData15[0]
                        };
                    end
                    6'b100000, 6'b100001, 6'b100010, 6'b100011,
                    6'b100100, 6'b100101, 6'b100110, 6'b100111: begin
                        readData = {
                                        readData14[3:0],
                                        readData13[3:0],
                                        readData12[3:0],
                                        readData11[3:0],
                                        readData10[3:0],
                                        readData9[3:0],
                                        readData8[3:0],
                                        readData7[3:0]
                        };
                    end
                    6'b101000, 6'b101001, 6'b101010, 6'b101011: begin
                        readData = {readData6[7:0],readData5[7:0],readData4[7:0],readData3[7:0]};
                    end
                    6'b101100, 6'b101101 : begin
                        readData = {readData2[16:9],readData2[7:0],readData1[16:9],readData1[7:0]};
                    end
                    6'b101110 : begin
                        readData = {readData0[34:27],readData0[25:18],readData0[16:9],readData0[7:0]};
                    end
                    default : begin
                        readData = 32'b0;
                    end
                endcase
            end        
            24576: begin
                width48 = 3'b000;
                width47 = 3'b000;
                width46 = 3'b000;
                width45 = 3'b000;
                width44 = 3'b000;
                width43 = 3'b000;
                width42 = 3'b000;
                width41 = 3'b000;
                width40 = 3'b000;
                width39 = 3'b000;
                width38 = 3'b000;
                width37 = 3'b000;
                width36 = 3'b000;
                width35 = 3'b000;
                width34 = 3'b000;
                width33 = 3'b000;
                width32 = 3'b000;
                width31 = 3'b000;
                width30 = 3'b000;
                width29 = 3'b000;
                width28 = 3'b000;
                width27 = 3'b000;
                width26 = 3'b000;
                width25 = 3'b000;
                width24 = 3'b000;
                width23 = 3'b000;
                width22 = 3'b000;
                width21 = 3'b000;
                width20 = 3'b000;
                width19 = 3'b000;
                width18 = 3'b000;
                width17 = 3'b000;
                width16 = 3'b001;
                width15 = 3'b001;
                width14 = 3'b001;
                width13 = 3'b001;
                width12 = 3'b001;
                width11 = 3'b001;
                width10 = 3'b001;
                width9 = 3'b001;
                width8 = 3'b001;
                width7 = 3'b001;
                width6 = 3'b001;
                width5 = 3'b001;
                width4 = 3'b001;
                width3 = 3'b001;
                width2 = 3'b001;
                width1 = 3'b001;

                writeAddr48 = {writeAddr[13:0]};
                writeAddr47 = {writeAddr[13:0]};
                writeAddr46 = {writeAddr[13:0]};
                writeAddr45 = {writeAddr[13:0]};
                writeAddr44 = {writeAddr[13:0]};
                writeAddr43 = {writeAddr[13:0]};
                writeAddr42 = {writeAddr[13:0]};
                writeAddr41 = {writeAddr[13:0]};
                writeAddr40 = {writeAddr[13:0]};
                writeAddr39 = {writeAddr[13:0]};
                writeAddr38 = {writeAddr[13:0]};
                writeAddr37 = {writeAddr[13:0]};
                writeAddr36 = {writeAddr[13:0]};
                writeAddr35 = {writeAddr[13:0]};
                writeAddr34 = {writeAddr[13:0]};
                writeAddr33 = {writeAddr[13:0]};
                writeAddr32 = {writeAddr[13:0]};
                writeAddr31 = {writeAddr[13:0]};
                writeAddr30 = {writeAddr[13:0]};
                writeAddr29 = {writeAddr[13:0]};
                writeAddr28 = {writeAddr[13:0]};
                writeAddr27 = {writeAddr[13:0]};
                writeAddr26 = {writeAddr[13:0]};
                writeAddr25 = {writeAddr[13:0]};
                writeAddr24 = {writeAddr[13:0]};
                writeAddr23 = {writeAddr[13:0]};
                writeAddr22 = {writeAddr[13:0]};
                writeAddr21 = {writeAddr[13:0]};
                writeAddr20 = {writeAddr[13:0]};
                writeAddr19 = {writeAddr[13:0]};
                writeAddr18 = {writeAddr[13:0]};
                writeAddr17 = {writeAddr[13:0]};
                writeAddr16 = {writeAddr[12:0], 1'b0};
                writeAddr15 = {writeAddr[12:0], 1'b0};
                writeAddr14 = {writeAddr[12:0], 1'b0};
                writeAddr13 = {writeAddr[12:0], 1'b0};
                writeAddr12 = {writeAddr[12:0], 1'b0};
                writeAddr11 = {writeAddr[12:0], 1'b0};
                writeAddr10 = {writeAddr[12:0], 1'b0};
                writeAddr9 = {writeAddr[12:0], 1'b0};
                writeAddr8 = {writeAddr[12:0], 1'b0};
                writeAddr7 = {writeAddr[12:0], 1'b0};
                writeAddr6 = {writeAddr[12:0], 1'b0};
                writeAddr5 = {writeAddr[12:0], 1'b0};
                writeAddr4 = {writeAddr[12:0], 1'b0};
                writeAddr3 = {writeAddr[12:0], 1'b0};
                writeAddr2 = {writeAddr[12:0], 1'b0};
                writeAddr1 = {writeAddr[12:0], 1'b0};

                readAddr48 = {writeAddr[13:0]};
                readAddr47 = {writeAddr[13:0]};
                readAddr46 = {writeAddr[13:0]};
                readAddr45 = {writeAddr[13:0]};
                readAddr44 = {writeAddr[13:0]};
                readAddr43 = {writeAddr[13:0]};
                readAddr42 = {writeAddr[13:0]};
                readAddr41 = {writeAddr[13:0]};
                readAddr40 = {writeAddr[13:0]};
                readAddr39 = {writeAddr[13:0]};
                readAddr38 = {writeAddr[13:0]};
                readAddr37 = {writeAddr[13:0]};
                readAddr36 = {writeAddr[13:0]};
                readAddr35 = {writeAddr[13:0]};
                readAddr34 = {writeAddr[13:0]};
                readAddr33 = {writeAddr[13:0]};
                readAddr32 = {writeAddr[13:0]};
                readAddr31 = {writeAddr[13:0]};
                readAddr30 = {writeAddr[13:0]};
                readAddr29 = {writeAddr[13:0]};
                readAddr28 = {writeAddr[13:0]};
                readAddr27 = {writeAddr[13:0]};
                readAddr26 = {writeAddr[13:0]};
                readAddr25 = {writeAddr[13:0]};
                readAddr24 = {writeAddr[13:0]};
                readAddr23 = {writeAddr[13:0]};
                readAddr22 = {writeAddr[13:0]};
                readAddr21 = {writeAddr[13:0]};
                readAddr20 = {writeAddr[13:0]};
                readAddr19 = {writeAddr[13:0]};
                readAddr18 = {writeAddr[13:0]};
                readAddr17 = {writeAddr[13:0]};
                readAddr16  = {readAddr[12:0],  1'b0};
                readAddr15  = {readAddr[12:0],  1'b0};
                readAddr14  = {readAddr[12:0],  1'b0};
                readAddr13  = {readAddr[12:0],  1'b0};
                readAddr12  = {readAddr[12:0],  1'b0};
                readAddr11  = {readAddr[12:0],  1'b0};
                readAddr10  = {readAddr[12:0],  1'b0};
                readAddr9  = {readAddr[12:0],  1'b0};
                readAddr8  = {readAddr[12:0],  1'b0};
                readAddr7  = {readAddr[12:0],  1'b0};
                readAddr6  = {readAddr[12:0],  1'b0};
                readAddr5  = {readAddr[12:0],  1'b0};
                readAddr4  = {readAddr[12:0],  1'b0};
                readAddr3  = {readAddr[12:0],  1'b0};
                readAddr2  = {readAddr[12:0],  1'b0};
                readAddr1  = {readAddr[12:0],  1'b0};

                writeData48 = {17'b0, writeData[31]};
                writeData47 = {17'b0, writeData[30]};
                writeData46 = {17'b0, writeData[29]};
                writeData45 = {17'b0, writeData[28]};
                writeData44 = {17'b0, writeData[27]};
                writeData43 = {17'b0, writeData[26]};
                writeData42 = {17'b0, writeData[25]};
                writeData41 = {17'b0, writeData[24]};
                writeData40 = {17'b0, writeData[23]};
                writeData39 = {17'b0, writeData[22]};
                writeData38 = {17'b0, writeData[21]};
                writeData37 = {17'b0, writeData[20]};
                writeData36 = {17'b0, writeData[19]};
                writeData35 = {17'b0, writeData[18]};
                writeData34 = {17'b0, writeData[17]};
                writeData33 = {17'b0, writeData[16]};
                writeData32 = {17'b0, writeData[15]};
                writeData31 = {17'b0, writeData[14]};
                writeData30 = {17'b0, writeData[13]};
                writeData29 = {17'b0, writeData[12]};
                writeData28 = {17'b0, writeData[11]};
                writeData27 = {17'b0, writeData[10]};
                writeData26 = {17'b0, writeData[9]};
                writeData25 = {17'b0, writeData[8]};
                writeData24 = {17'b0, writeData[7]};
                writeData23 = {17'b0, writeData[6]};
                writeData22 = {17'b0, writeData[5]};
                writeData21 = {17'b0, writeData[4]};
                writeData20 = {17'b0, writeData[3]};
                writeData19 = {17'b0, writeData[2]};
                writeData18 = {17'b0, writeData[1]};
                writeData17 = {17'b0, writeData[0]};
                writeData16 = {16'b0, writeData[31:30]};
                writeData15 = {16'b0, writeData[29:28]};
                writeData14 = {16'b0, writeData[27:26]};
                writeData13 = {16'b0, writeData[25:24]};
                writeData12 = {16'b0, writeData[23:22]};
                writeData11 = {16'b0, writeData[21:20]};
                writeData10 = {16'b0, writeData[19:18]};
                writeData9 = {16'b0, writeData[17:16]};
                writeData8 = {16'b0, writeData[15:14]};
                writeData7 = {16'b0, writeData[13:12]};
                writeData6 = {16'b0, writeData[11:10]};
                writeData5 = {16'b0, writeData[9:8]};
                writeData4 = {16'b0, writeData[7:6]};
                writeData3 = {16'b0, writeData[5:4]};
                writeData2 = {16'b0, writeData[3:2]};
                writeData1 = {16'b0, writeData[1:0]};

                case (writeAddr[14:9])
                    6'b000000, 6'b000001, 6'b000010, 6'b000011,
                    6'b000100, 6'b000101, 6'b000110, 6'b000111,
                    6'b001000, 6'b001001, 6'b001010, 6'b001011,
                    6'b001100, 6'b001101, 6'b001110, 6'b001111,
                    6'b010000, 6'b010001, 6'b010010, 6'b010011,
                    6'b010100, 6'b010101, 6'b010110, 6'b010111,
                    6'b011000, 6'b011001, 6'b011010, 6'b011011,
                    6'b011100, 6'b011101, 6'b011110, 6'b011111 : begin
                        wen_a48 = {1'b0, wen};
                        wen_a47 = {1'b0, wen};
                        wen_a46 = {1'b0, wen};
                        wen_a45 = {1'b0, wen};
                        wen_a44 = {1'b0, wen};
                        wen_a43 = {1'b0, wen};
                        wen_a42 = {1'b0, wen};
                        wen_a41 = {1'b0, wen};
                        wen_a40 = {1'b0, wen};
                        wen_a39 = {1'b0, wen};
                        wen_a38 = {1'b0, wen};
                        wen_a37 = {1'b0, wen};
                        wen_a36 = {1'b0, wen};
                        wen_a35 = {1'b0, wen};
                        wen_a34 = {1'b0, wen};
                        wen_a33 = {1'b0, wen};
                        wen_a32 = {1'b0, wen};
                        wen_a31 = {1'b0, wen};
                        wen_a30 = {1'b0, wen};
                        wen_a29 = {1'b0, wen};
                        wen_a28 = {1'b0, wen};
                        wen_a27 = {1'b0, wen};
                        wen_a26 = {1'b0, wen};
                        wen_a25 = {1'b0, wen};
                        wen_a24 = {1'b0, wen};
                        wen_a23 = {1'b0, wen};
                        wen_a22 = {1'b0, wen};
                        wen_a21 = {1'b0, wen};
                        wen_a20 = {1'b0, wen};
                        wen_a19 = {1'b0, wen};
                        wen_a18 = {1'b0, wen};
                        wen_a17 = {1'b0, wen};
                        wen_a16 = {1'b0, 1'b0};
                        wen_a15 = {1'b0, 1'b0};
                        wen_a14 = {1'b0, 1'b0};
                        wen_a13 = {1'b0, 1'b0};
                        wen_a12 = {1'b0, 1'b0};
                        wen_a11 = {1'b0, 1'b0};
                        wen_a10 = {1'b0, 1'b0};
                        wen_a9 = {1'b0, 1'b0};
                        wen_a8 = {1'b0, 1'b0};
                        wen_a7 = {1'b0, 1'b0};
                        wen_a6 = {1'b0, 1'b0};
                        wen_a5 = {1'b0, 1'b0};
                        wen_a4 = {1'b0, 1'b0};
                        wen_a3 = {1'b0, 1'b0};
                        wen_a2 = {1'b0, 1'b0};
                        wen_a1 = {1'b0, 1'b0};
                    end
                    6'b100000, 6'b100001, 6'b100010, 6'b100011,
                    6'b100100, 6'b100101, 6'b100110, 6'b100111,
                    6'b101000, 6'b101001, 6'b101010, 6'b101011,
                    6'b101100, 6'b101101, 6'b101110, 6'b101111 : begin
                        wen_a48 = {1'b0, 1'b0};
                        wen_a47 = {1'b0, 1'b0};
                        wen_a46 = {1'b0, 1'b0};
                        wen_a45 = {1'b0, 1'b0};
                        wen_a44 = {1'b0, 1'b0};
                        wen_a43 = {1'b0, 1'b0};
                        wen_a42 = {1'b0, 1'b0};
                        wen_a41 = {1'b0, 1'b0};
                        wen_a40 = {1'b0, 1'b0};
                        wen_a39 = {1'b0, 1'b0};
                        wen_a38 = {1'b0, 1'b0};
                        wen_a37 = {1'b0, 1'b0};
                        wen_a36 = {1'b0, 1'b0};
                        wen_a35 = {1'b0, 1'b0};
                        wen_a34 = {1'b0, 1'b0};
                        wen_a33 = {1'b0, 1'b0};
                        wen_a32 = {1'b0, 1'b0};
                        wen_a31 = {1'b0, 1'b0};
                        wen_a30 = {1'b0, 1'b0};
                        wen_a29 = {1'b0, 1'b0};
                        wen_a28 = {1'b0, 1'b0};
                        wen_a27 = {1'b0, 1'b0};
                        wen_a26 = {1'b0, 1'b0};
                        wen_a25 = {1'b0, 1'b0};
                        wen_a24 = {1'b0, 1'b0};
                        wen_a23 = {1'b0, 1'b0};
                        wen_a22 = {1'b0, 1'b0};
                        wen_a21 = {1'b0, 1'b0};
                        wen_a20 = {1'b0, 1'b0};
                        wen_a19 = {1'b0, 1'b0};
                        wen_a18 = {1'b0, 1'b0};
                        wen_a17 = {1'b0, 1'b0};
                        wen_a16 = {1'b0, wen};
                        wen_a15 = {1'b0, wen};
                        wen_a14 = {1'b0, wen};
                        wen_a13 = {1'b0, wen};
                        wen_a12 = {1'b0, wen};
                        wen_a11 = {1'b0, wen};
                        wen_a10 = {1'b0, wen};
                        wen_a9 = {1'b0, wen};
                        wen_a8 = {1'b0, wen};
                        wen_a7 = {1'b0, wen};
                        wen_a6 = {1'b0, wen};
                        wen_a5 = {1'b0, wen};
                        wen_a4 = {1'b0, wen};
                        wen_a3 = {1'b0, wen};
                        wen_a2 = {1'b0, wen};
                        wen_a1 = {1'b0, wen};
                    end
                    default : begin
                        wen_a48 = {1'b0, 1'b0};
                        wen_a47 = {1'b0, 1'b0};
                        wen_a46 = {1'b0, 1'b0};
                        wen_a45 = {1'b0, 1'b0};
                        wen_a44 = {1'b0, 1'b0};
                        wen_a43 = {1'b0, 1'b0};
                        wen_a42 = {1'b0, 1'b0};
                        wen_a41 = {1'b0, 1'b0};
                        wen_a40 = {1'b0, 1'b0};
                        wen_a39 = {1'b0, 1'b0};
                        wen_a38 = {1'b0, 1'b0};
                        wen_a37 = {1'b0, 1'b0};
                        wen_a36 = {1'b0, 1'b0};
                        wen_a35 = {1'b0, 1'b0};
                        wen_a34 = {1'b0, 1'b0};
                        wen_a33 = {1'b0, 1'b0};
                        wen_a32 = {1'b0, 1'b0};
                        wen_a31 = {1'b0, 1'b0};
                        wen_a30 = {1'b0, 1'b0};
                        wen_a29 = {1'b0, 1'b0};
                        wen_a28 = {1'b0, 1'b0};
                        wen_a27 = {1'b0, 1'b0};
                        wen_a26 = {1'b0, 1'b0};
                        wen_a25 = {1'b0, 1'b0};
                        wen_a24 = {1'b0, 1'b0};
                        wen_a23 = {1'b0, 1'b0};
                        wen_a22 = {1'b0, 1'b0};
                        wen_a21 = {1'b0, 1'b0};
                        wen_a20 = {1'b0, 1'b0};
                        wen_a19 = {1'b0, 1'b0};
                        wen_a18 = {1'b0, 1'b0};
                        wen_a17 = {1'b0, 1'b0};
                        wen_a16 = {1'b0, 1'b0};
                        wen_a15 = {1'b0, 1'b0};
                        wen_a14 = {1'b0, 1'b0};
                        wen_a13 = {1'b0, 1'b0};
                        wen_a12 = {1'b0, 1'b0};
                        wen_a11 = {1'b0, 1'b0};
                        wen_a10 = {1'b0, 1'b0};
                        wen_a9 = {1'b0, 1'b0};
                        wen_a8 = {1'b0, 1'b0};
                        wen_a7 = {1'b0, 1'b0};
                        wen_a6 = {1'b0, 1'b0};
                        wen_a5 = {1'b0, 1'b0};
                        wen_a4 = {1'b0, 1'b0};
                        wen_a3 = {1'b0, 1'b0};
                        wen_a2 = {1'b0, 1'b0};
                        wen_a1 = {1'b0, 1'b0};
                    end
                endcase

                case (ckRdAddr[14:9])
                    6'b000000, 6'b000001, 6'b000010, 6'b000011,
                    6'b000100, 6'b000101, 6'b000110, 6'b000111,
                    6'b001000, 6'b001001, 6'b001010, 6'b001011,
                    6'b001100, 6'b001101, 6'b001110, 6'b001111,
                    6'b010000, 6'b010001, 6'b010010, 6'b010011,
                    6'b010100, 6'b010101, 6'b010110, 6'b010111,
                    6'b011000, 6'b011001, 6'b011010, 6'b011011,
                    6'b011100, 6'b011101, 6'b011110, 6'b011111 : begin
                        readData = {
                                        readData48[0],
                                        readData47[0],
                                        readData46[0],
                                        readData45[0],
                                        readData44[0],
                                        readData43[0],
                                        readData42[0],
                                        readData41[0],
                                        readData40[0],
                                        readData39[0],
                                        readData38[0],
                                        readData37[0],
                                        readData36[0],
                                        readData35[0],
                                        readData34[0],
                                        readData33[0],
                                        readData32[0],
                                        readData31[0],
                                        readData30[0],
                                        readData29[0],
                                        readData28[0],
                                        readData27[0],
                                        readData26[0],
                                        readData25[0],
                                        readData24[0],
                                        readData23[0],
                                        readData22[0],
                                        readData21[0],
                                        readData20[0],
                                        readData19[0],
                                        readData18[0],
                                        readData17[0]
                        };
                    end
                    6'b100000, 6'b100001, 6'b100010, 6'b100011,
                    6'b100100, 6'b100101, 6'b100110, 6'b100111,
                    6'b101000, 6'b101001, 6'b101010, 6'b101011,
                    6'b101100, 6'b101101, 6'b101110, 6'b101111 : begin
                        readData = {
                                        readData16[1:0],
                                        readData15[1:0],
                                        readData14[1:0],
                                        readData13[1:0],
                                        readData12[1:0],
                                        readData11[1:0],
                                        readData10[1:0],
                                        readData9[1:0],
                                        readData8[1:0],
                                        readData7[1:0],
                                        readData6[1:0],
                                        readData5[1:0],
                                        readData4[1:0],
                                        readData3[1:0],
                                        readData2[1:0],
                                        readData1[1:0]
                        };
                    end
                    default : begin
                        readData = 32'b0;
                    end
                endcase
            end        
            25088: begin
                width48 = 3'b000;
                width47 = 3'b000;
                width46 = 3'b000;
                width45 = 3'b000;
                width44 = 3'b000;
                width43 = 3'b000;
                width42 = 3'b000;
                width41 = 3'b000;
                width40 = 3'b000;
                width39 = 3'b000;
                width38 = 3'b000;
                width37 = 3'b000;
                width36 = 3'b000;
                width35 = 3'b000;
                width34 = 3'b000;
                width33 = 3'b000;
                width32 = 3'b000;
                width31 = 3'b000;
                width30 = 3'b000;
                width29 = 3'b000;
                width28 = 3'b000;
                width27 = 3'b000;
                width26 = 3'b000;
                width25 = 3'b000;
                width24 = 3'b000;
                width23 = 3'b000;
                width22 = 3'b000;
                width21 = 3'b000;
                width20 = 3'b000;
                width19 = 3'b000;
                width18 = 3'b000;
                width17 = 3'b000;
                width16 = 3'b001;
                width15 = 3'b001;
                width14 = 3'b001;
                width13 = 3'b001;
                width12 = 3'b001;
                width11 = 3'b001;
                width10 = 3'b001;
                width9 = 3'b001;
                width8 = 3'b001;
                width7 = 3'b001;
                width6 = 3'b001;
                width5 = 3'b001;
                width4 = 3'b001;
                width3 = 3'b001;
                width2 = 3'b001;
                width1 = 3'b001;
                width0 = 3'b101;

                writeAddr48 = {writeAddr[13:0]};
                writeAddr47 = {writeAddr[13:0]};
                writeAddr46 = {writeAddr[13:0]};
                writeAddr45 = {writeAddr[13:0]};
                writeAddr44 = {writeAddr[13:0]};
                writeAddr43 = {writeAddr[13:0]};
                writeAddr42 = {writeAddr[13:0]};
                writeAddr41 = {writeAddr[13:0]};
                writeAddr40 = {writeAddr[13:0]};
                writeAddr39 = {writeAddr[13:0]};
                writeAddr38 = {writeAddr[13:0]};
                writeAddr37 = {writeAddr[13:0]};
                writeAddr36 = {writeAddr[13:0]};
                writeAddr35 = {writeAddr[13:0]};
                writeAddr34 = {writeAddr[13:0]};
                writeAddr33 = {writeAddr[13:0]};
                writeAddr32 = {writeAddr[13:0]};
                writeAddr31 = {writeAddr[13:0]};
                writeAddr30 = {writeAddr[13:0]};
                writeAddr29 = {writeAddr[13:0]};
                writeAddr28 = {writeAddr[13:0]};
                writeAddr27 = {writeAddr[13:0]};
                writeAddr26 = {writeAddr[13:0]};
                writeAddr25 = {writeAddr[13:0]};
                writeAddr24 = {writeAddr[13:0]};
                writeAddr23 = {writeAddr[13:0]};
                writeAddr22 = {writeAddr[13:0]};
                writeAddr21 = {writeAddr[13:0]};
                writeAddr20 = {writeAddr[13:0]};
                writeAddr19 = {writeAddr[13:0]};
                writeAddr18 = {writeAddr[13:0]};
                writeAddr17 = {writeAddr[13:0]};
                writeAddr16 = {writeAddr[12:0], 1'b0};
                writeAddr15 = {writeAddr[12:0], 1'b0};
                writeAddr14 = {writeAddr[12:0], 1'b0};
                writeAddr13 = {writeAddr[12:0], 1'b0};
                writeAddr12 = {writeAddr[12:0], 1'b0};
                writeAddr11 = {writeAddr[12:0], 1'b0};
                writeAddr10 = {writeAddr[12:0], 1'b0};
                writeAddr9 = {writeAddr[12:0], 1'b0};
                writeAddr8 = {writeAddr[12:0], 1'b0};
                writeAddr7 = {writeAddr[12:0], 1'b0};
                writeAddr6 = {writeAddr[12:0], 1'b0};
                writeAddr5 = {writeAddr[12:0], 1'b0};
                writeAddr4 = {writeAddr[12:0], 1'b0};
                writeAddr3 = {writeAddr[12:0], 1'b0};
                writeAddr2 = {writeAddr[12:0], 1'b0};
                writeAddr1 = {writeAddr[12:0], 1'b0};
                writeAddr0 = {writeAddr[8:0], 5'b0};

                readAddr48 = {writeAddr[13:0]};
                readAddr47 = {writeAddr[13:0]};
                readAddr46 = {writeAddr[13:0]};
                readAddr45 = {writeAddr[13:0]};
                readAddr44 = {writeAddr[13:0]};
                readAddr43 = {writeAddr[13:0]};
                readAddr42 = {writeAddr[13:0]};
                readAddr41 = {writeAddr[13:0]};
                readAddr40 = {writeAddr[13:0]};
                readAddr39 = {writeAddr[13:0]};
                readAddr38 = {writeAddr[13:0]};
                readAddr37 = {writeAddr[13:0]};
                readAddr36 = {writeAddr[13:0]};
                readAddr35 = {writeAddr[13:0]};
                readAddr34 = {writeAddr[13:0]};
                readAddr33 = {writeAddr[13:0]};
                readAddr32 = {writeAddr[13:0]};
                readAddr31 = {writeAddr[13:0]};
                readAddr30 = {writeAddr[13:0]};
                readAddr29 = {writeAddr[13:0]};
                readAddr28 = {writeAddr[13:0]};
                readAddr27 = {writeAddr[13:0]};
                readAddr26 = {writeAddr[13:0]};
                readAddr25 = {writeAddr[13:0]};
                readAddr24 = {writeAddr[13:0]};
                readAddr23 = {writeAddr[13:0]};
                readAddr22 = {writeAddr[13:0]};
                readAddr21 = {writeAddr[13:0]};
                readAddr20 = {writeAddr[13:0]};
                readAddr19 = {writeAddr[13:0]};
                readAddr18 = {writeAddr[13:0]};
                readAddr17 = {writeAddr[13:0]};
                readAddr16  = {readAddr[12:0],  1'b0};
                readAddr15  = {readAddr[12:0],  1'b0};
                readAddr14  = {readAddr[12:0],  1'b0};
                readAddr13  = {readAddr[12:0],  1'b0};
                readAddr12  = {readAddr[12:0],  1'b0};
                readAddr11  = {readAddr[12:0],  1'b0};
                readAddr10  = {readAddr[12:0],  1'b0};
                readAddr9  = {readAddr[12:0],  1'b0};
                readAddr8  = {readAddr[12:0],  1'b0};
                readAddr7  = {readAddr[12:0],  1'b0};
                readAddr6  = {readAddr[12:0],  1'b0};
                readAddr5  = {readAddr[12:0],  1'b0};
                readAddr4  = {readAddr[12:0],  1'b0};
                readAddr3  = {readAddr[12:0],  1'b0};
                readAddr2  = {readAddr[12:0],  1'b0};
                readAddr1  = {readAddr[12:0],  1'b0};
                readAddr0  = {readAddr[8:0],  5'b0};

                writeData48 = {17'b0, writeData[31]};
                writeData47 = {17'b0, writeData[30]};
                writeData46 = {17'b0, writeData[29]};
                writeData45 = {17'b0, writeData[28]};
                writeData44 = {17'b0, writeData[27]};
                writeData43 = {17'b0, writeData[26]};
                writeData42 = {17'b0, writeData[25]};
                writeData41 = {17'b0, writeData[24]};
                writeData40 = {17'b0, writeData[23]};
                writeData39 = {17'b0, writeData[22]};
                writeData38 = {17'b0, writeData[21]};
                writeData37 = {17'b0, writeData[20]};
                writeData36 = {17'b0, writeData[19]};
                writeData35 = {17'b0, writeData[18]};
                writeData34 = {17'b0, writeData[17]};
                writeData33 = {17'b0, writeData[16]};
                writeData32 = {17'b0, writeData[15]};
                writeData31 = {17'b0, writeData[14]};
                writeData30 = {17'b0, writeData[13]};
                writeData29 = {17'b0, writeData[12]};
                writeData28 = {17'b0, writeData[11]};
                writeData27 = {17'b0, writeData[10]};
                writeData26 = {17'b0, writeData[9]};
                writeData25 = {17'b0, writeData[8]};
                writeData24 = {17'b0, writeData[7]};
                writeData23 = {17'b0, writeData[6]};
                writeData22 = {17'b0, writeData[5]};
                writeData21 = {17'b0, writeData[4]};
                writeData20 = {17'b0, writeData[3]};
                writeData19 = {17'b0, writeData[2]};
                writeData18 = {17'b0, writeData[1]};
                writeData17 = {17'b0, writeData[0]};
                writeData16 = {16'b0, writeData[31:30]};
                writeData15 = {16'b0, writeData[29:28]};
                writeData14 = {16'b0, writeData[27:26]};
                writeData13 = {16'b0, writeData[25:24]};
                writeData12 = {16'b0, writeData[23:22]};
                writeData11 = {16'b0, writeData[21:20]};
                writeData10 = {16'b0, writeData[19:18]};
                writeData9 = {16'b0, writeData[17:16]};
                writeData8 = {16'b0, writeData[15:14]};
                writeData7 = {16'b0, writeData[13:12]};
                writeData6 = {16'b0, writeData[11:10]};
                writeData5 = {16'b0, writeData[9:8]};
                writeData4 = {16'b0, writeData[7:6]};
                writeData3 = {16'b0, writeData[5:4]};
                writeData2 = {16'b0, writeData[3:2]};
                writeData1 = {16'b0, writeData[1:0]};
                writeData0 = {1'b0, writeData[31:24], 1'b0, writeData[23:16], 1'b0, writeData[15:8], 1'b0, writeData[7:0]};

                case (writeAddr[14:9])
                    6'b000000, 6'b000001, 6'b000010, 6'b000011,
                    6'b000100, 6'b000101, 6'b000110, 6'b000111,
                    6'b001000, 6'b001001, 6'b001010, 6'b001011,
                    6'b001100, 6'b001101, 6'b001110, 6'b001111,
                    6'b010000, 6'b010001, 6'b010010, 6'b010011,
                    6'b010100, 6'b010101, 6'b010110, 6'b010111,
                    6'b011000, 6'b011001, 6'b011010, 6'b011011,
                    6'b011100, 6'b011101, 6'b011110, 6'b011111 : begin
                        wen_a48 = {1'b0, wen};
                        wen_a47 = {1'b0, wen};
                        wen_a46 = {1'b0, wen};
                        wen_a45 = {1'b0, wen};
                        wen_a44 = {1'b0, wen};
                        wen_a43 = {1'b0, wen};
                        wen_a42 = {1'b0, wen};
                        wen_a41 = {1'b0, wen};
                        wen_a40 = {1'b0, wen};
                        wen_a39 = {1'b0, wen};
                        wen_a38 = {1'b0, wen};
                        wen_a37 = {1'b0, wen};
                        wen_a36 = {1'b0, wen};
                        wen_a35 = {1'b0, wen};
                        wen_a34 = {1'b0, wen};
                        wen_a33 = {1'b0, wen};
                        wen_a32 = {1'b0, wen};
                        wen_a31 = {1'b0, wen};
                        wen_a30 = {1'b0, wen};
                        wen_a29 = {1'b0, wen};
                        wen_a28 = {1'b0, wen};
                        wen_a27 = {1'b0, wen};
                        wen_a26 = {1'b0, wen};
                        wen_a25 = {1'b0, wen};
                        wen_a24 = {1'b0, wen};
                        wen_a23 = {1'b0, wen};
                        wen_a22 = {1'b0, wen};
                        wen_a21 = {1'b0, wen};
                        wen_a20 = {1'b0, wen};
                        wen_a19 = {1'b0, wen};
                        wen_a18 = {1'b0, wen};
                        wen_a17 = {1'b0, wen};
                        wen_a16 = {1'b0, 1'b0};
                        wen_a15 = {1'b0, 1'b0};
                        wen_a14 = {1'b0, 1'b0};
                        wen_a13 = {1'b0, 1'b0};
                        wen_a12 = {1'b0, 1'b0};
                        wen_a11 = {1'b0, 1'b0};
                        wen_a10 = {1'b0, 1'b0};
                        wen_a9 = {1'b0, 1'b0};
                        wen_a8 = {1'b0, 1'b0};
                        wen_a7 = {1'b0, 1'b0};
                        wen_a6 = {1'b0, 1'b0};
                        wen_a5 = {1'b0, 1'b0};
                        wen_a4 = {1'b0, 1'b0};
                        wen_a3 = {1'b0, 1'b0};
                        wen_a2 = {1'b0, 1'b0};
                        wen_a1 = {1'b0, 1'b0};
                        wen_a0 = {1'b0, 1'b0};
                        wen_b0 = {1'b0, 1'b0};
                    end
                    6'b100000, 6'b100001, 6'b100010, 6'b100011,
                    6'b100100, 6'b100101, 6'b100110, 6'b100111,
                    6'b101000, 6'b101001, 6'b101010, 6'b101011,
                    6'b101100, 6'b101101, 6'b101110, 6'b101111 : begin
                        wen_a48 = {1'b0, 1'b0};
                        wen_a47 = {1'b0, 1'b0};
                        wen_a46 = {1'b0, 1'b0};
                        wen_a45 = {1'b0, 1'b0};
                        wen_a44 = {1'b0, 1'b0};
                        wen_a43 = {1'b0, 1'b0};
                        wen_a42 = {1'b0, 1'b0};
                        wen_a41 = {1'b0, 1'b0};
                        wen_a40 = {1'b0, 1'b0};
                        wen_a39 = {1'b0, 1'b0};
                        wen_a38 = {1'b0, 1'b0};
                        wen_a37 = {1'b0, 1'b0};
                        wen_a36 = {1'b0, 1'b0};
                        wen_a35 = {1'b0, 1'b0};
                        wen_a34 = {1'b0, 1'b0};
                        wen_a33 = {1'b0, 1'b0};
                        wen_a32 = {1'b0, 1'b0};
                        wen_a31 = {1'b0, 1'b0};
                        wen_a30 = {1'b0, 1'b0};
                        wen_a29 = {1'b0, 1'b0};
                        wen_a28 = {1'b0, 1'b0};
                        wen_a27 = {1'b0, 1'b0};
                        wen_a26 = {1'b0, 1'b0};
                        wen_a25 = {1'b0, 1'b0};
                        wen_a24 = {1'b0, 1'b0};
                        wen_a23 = {1'b0, 1'b0};
                        wen_a22 = {1'b0, 1'b0};
                        wen_a21 = {1'b0, 1'b0};
                        wen_a20 = {1'b0, 1'b0};
                        wen_a19 = {1'b0, 1'b0};
                        wen_a18 = {1'b0, 1'b0};
                        wen_a17 = {1'b0, 1'b0};
                        wen_a16 = {1'b0, wen};
                        wen_a15 = {1'b0, wen};
                        wen_a14 = {1'b0, wen};
                        wen_a13 = {1'b0, wen};
                        wen_a12 = {1'b0, wen};
                        wen_a11 = {1'b0, wen};
                        wen_a10 = {1'b0, wen};
                        wen_a9 = {1'b0, wen};
                        wen_a8 = {1'b0, wen};
                        wen_a7 = {1'b0, wen};
                        wen_a6 = {1'b0, wen};
                        wen_a5 = {1'b0, wen};
                        wen_a4 = {1'b0, wen};
                        wen_a3 = {1'b0, wen};
                        wen_a2 = {1'b0, wen};
                        wen_a1 = {1'b0, wen};
                        wen_a0 = {1'b0, 1'b0};
                        wen_b0 = {1'b0, 1'b0};
                    end
                    6'b110000 : begin
                        wen_a48 = {1'b0, 1'b0};
                        wen_a47 = {1'b0, 1'b0};
                        wen_a46 = {1'b0, 1'b0};
                        wen_a45 = {1'b0, 1'b0};
                        wen_a44 = {1'b0, 1'b0};
                        wen_a43 = {1'b0, 1'b0};
                        wen_a42 = {1'b0, 1'b0};
                        wen_a41 = {1'b0, 1'b0};
                        wen_a40 = {1'b0, 1'b0};
                        wen_a39 = {1'b0, 1'b0};
                        wen_a38 = {1'b0, 1'b0};
                        wen_a37 = {1'b0, 1'b0};
                        wen_a36 = {1'b0, 1'b0};
                        wen_a35 = {1'b0, 1'b0};
                        wen_a34 = {1'b0, 1'b0};
                        wen_a33 = {1'b0, 1'b0};
                        wen_a32 = {1'b0, 1'b0};
                        wen_a31 = {1'b0, 1'b0};
                        wen_a30 = {1'b0, 1'b0};
                        wen_a29 = {1'b0, 1'b0};
                        wen_a28 = {1'b0, 1'b0};
                        wen_a27 = {1'b0, 1'b0};
                        wen_a26 = {1'b0, 1'b0};
                        wen_a25 = {1'b0, 1'b0};
                        wen_a24 = {1'b0, 1'b0};
                        wen_a23 = {1'b0, 1'b0};
                        wen_a22 = {1'b0, 1'b0};
                        wen_a21 = {1'b0, 1'b0};
                        wen_a20 = {1'b0, 1'b0};
                        wen_a19 = {1'b0, 1'b0};
                        wen_a18 = {1'b0, 1'b0};
                        wen_a17 = {1'b0, 1'b0};
                        wen_a16 = {1'b0, 1'b0};
                        wen_a15 = {1'b0, 1'b0};
                        wen_a14 = {1'b0, 1'b0};
                        wen_a13 = {1'b0, 1'b0};
                        wen_a12 = {1'b0, 1'b0};
                        wen_a11 = {1'b0, 1'b0};
                        wen_a10 = {1'b0, 1'b0};
                        wen_a9 = {1'b0, 1'b0};
                        wen_a8 = {1'b0, 1'b0};
                        wen_a7 = {1'b0, 1'b0};
                        wen_a6 = {1'b0, 1'b0};
                        wen_a5 = {1'b0, 1'b0};
                        wen_a4 = {1'b0, 1'b0};
                        wen_a3 = {1'b0, 1'b0};
                        wen_a2 = {1'b0, 1'b0};
                        wen_a1 = {1'b0, 1'b0};
                        wen_a0 = {wen, wen};
                        wen_b0 = {wen, wen};
                    end
                    default : begin
                        wen_a48 = {1'b0, 1'b0};
                        wen_a47 = {1'b0, 1'b0};
                        wen_a46 = {1'b0, 1'b0};
                        wen_a45 = {1'b0, 1'b0};
                        wen_a44 = {1'b0, 1'b0};
                        wen_a43 = {1'b0, 1'b0};
                        wen_a42 = {1'b0, 1'b0};
                        wen_a41 = {1'b0, 1'b0};
                        wen_a40 = {1'b0, 1'b0};
                        wen_a39 = {1'b0, 1'b0};
                        wen_a38 = {1'b0, 1'b0};
                        wen_a37 = {1'b0, 1'b0};
                        wen_a36 = {1'b0, 1'b0};
                        wen_a35 = {1'b0, 1'b0};
                        wen_a34 = {1'b0, 1'b0};
                        wen_a33 = {1'b0, 1'b0};
                        wen_a32 = {1'b0, 1'b0};
                        wen_a31 = {1'b0, 1'b0};
                        wen_a30 = {1'b0, 1'b0};
                        wen_a29 = {1'b0, 1'b0};
                        wen_a28 = {1'b0, 1'b0};
                        wen_a27 = {1'b0, 1'b0};
                        wen_a26 = {1'b0, 1'b0};
                        wen_a25 = {1'b0, 1'b0};
                        wen_a24 = {1'b0, 1'b0};
                        wen_a23 = {1'b0, 1'b0};
                        wen_a22 = {1'b0, 1'b0};
                        wen_a21 = {1'b0, 1'b0};
                        wen_a20 = {1'b0, 1'b0};
                        wen_a19 = {1'b0, 1'b0};
                        wen_a18 = {1'b0, 1'b0};
                        wen_a17 = {1'b0, 1'b0};
                        wen_a16 = {1'b0, 1'b0};
                        wen_a15 = {1'b0, 1'b0};
                        wen_a14 = {1'b0, 1'b0};
                        wen_a13 = {1'b0, 1'b0};
                        wen_a12 = {1'b0, 1'b0};
                        wen_a11 = {1'b0, 1'b0};
                        wen_a10 = {1'b0, 1'b0};
                        wen_a9 = {1'b0, 1'b0};
                        wen_a8 = {1'b0, 1'b0};
                        wen_a7 = {1'b0, 1'b0};
                        wen_a6 = {1'b0, 1'b0};
                        wen_a5 = {1'b0, 1'b0};
                        wen_a4 = {1'b0, 1'b0};
                        wen_a3 = {1'b0, 1'b0};
                        wen_a2 = {1'b0, 1'b0};
                        wen_a1 = {1'b0, 1'b0};
                        wen_a0 = {1'b0, 1'b0};
                        wen_b0 = {1'b0, 1'b0};
                    end
                endcase

                case (ckRdAddr[14:9])
                    6'b000000, 6'b000001, 6'b000010, 6'b000011,
                    6'b000100, 6'b000101, 6'b000110, 6'b000111,
                    6'b001000, 6'b001001, 6'b001010, 6'b001011,
                    6'b001100, 6'b001101, 6'b001110, 6'b001111,
                    6'b010000, 6'b010001, 6'b010010, 6'b010011,
                    6'b010100, 6'b010101, 6'b010110, 6'b010111,
                    6'b011000, 6'b011001, 6'b011010, 6'b011011,
                    6'b011100, 6'b011101, 6'b011110, 6'b011111 : begin
                        readData = {
                                        readData48[0],
                                        readData47[0],
                                        readData46[0],
                                        readData45[0],
                                        readData44[0],
                                        readData43[0],
                                        readData42[0],
                                        readData41[0],
                                        readData40[0],
                                        readData39[0],
                                        readData38[0],
                                        readData37[0],
                                        readData36[0],
                                        readData35[0],
                                        readData34[0],
                                        readData33[0],
                                        readData32[0],
                                        readData31[0],
                                        readData30[0],
                                        readData29[0],
                                        readData28[0],
                                        readData27[0],
                                        readData26[0],
                                        readData25[0],
                                        readData24[0],
                                        readData23[0],
                                        readData22[0],
                                        readData21[0],
                                        readData20[0],
                                        readData19[0],
                                        readData18[0],
                                        readData17[0]
                        };
                    end
                    6'b100000, 6'b100001, 6'b100010, 6'b100011,
                    6'b100100, 6'b100101, 6'b100110, 6'b100111,
                    6'b101000, 6'b101001, 6'b101010, 6'b101011,
                    6'b101100, 6'b101101, 6'b101110, 6'b101111 : begin
                        readData = {
                                        readData16[1:0],
                                        readData15[1:0],
                                        readData14[1:0],
                                        readData13[1:0],
                                        readData12[1:0],
                                        readData11[1:0],
                                        readData10[1:0],
                                        readData9[1:0],
                                        readData8[1:0],
                                        readData7[1:0],
                                        readData6[1:0],
                                        readData5[1:0],
                                        readData4[1:0],
                                        readData3[1:0],
                                        readData2[1:0],
                                        readData1[1:0]
                        };
                    end
                    6'b110000 : begin
                        readData = {readData0[34:27],readData0[25:18],readData0[16:9],readData0[7:0]};
                    end
                    default : begin
                        readData = 32'b0;
                    end
                endcase
            end        
            25600: begin
                width50 = 3'b000;
                width49 = 3'b000;
                width48 = 3'b000;
                width47 = 3'b000;
                width46 = 3'b000;
                width45 = 3'b000;
                width44 = 3'b000;
                width43 = 3'b000;
                width42 = 3'b000;
                width41 = 3'b000;
                width40 = 3'b000;
                width39 = 3'b000;
                width38 = 3'b000;
                width37 = 3'b000;
                width36 = 3'b000;
                width35 = 3'b000;
                width34 = 3'b000;
                width33 = 3'b000;
                width32 = 3'b000;
                width31 = 3'b000;
                width30 = 3'b000;
                width29 = 3'b000;
                width28 = 3'b000;
                width27 = 3'b000;
                width26 = 3'b000;
                width25 = 3'b000;
                width24 = 3'b000;
                width23 = 3'b000;
                width22 = 3'b000;
                width21 = 3'b000;
                width20 = 3'b000;
                width19 = 3'b000;
                width18 = 3'b001;
                width17 = 3'b001;
                width16 = 3'b001;
                width15 = 3'b001;
                width14 = 3'b001;
                width13 = 3'b001;
                width12 = 3'b001;
                width11 = 3'b001;
                width10 = 3'b001;
                width9 = 3'b001;
                width8 = 3'b001;
                width7 = 3'b001;
                width6 = 3'b001;
                width5 = 3'b001;
                width4 = 3'b001;
                width3 = 3'b001;
                width2 = 3'b100;
                width1 = 3'b100;

                writeAddr50 = {writeAddr[13:0]};
                writeAddr49 = {writeAddr[13:0]};
                writeAddr48 = {writeAddr[13:0]};
                writeAddr47 = {writeAddr[13:0]};
                writeAddr46 = {writeAddr[13:0]};
                writeAddr45 = {writeAddr[13:0]};
                writeAddr44 = {writeAddr[13:0]};
                writeAddr43 = {writeAddr[13:0]};
                writeAddr42 = {writeAddr[13:0]};
                writeAddr41 = {writeAddr[13:0]};
                writeAddr40 = {writeAddr[13:0]};
                writeAddr39 = {writeAddr[13:0]};
                writeAddr38 = {writeAddr[13:0]};
                writeAddr37 = {writeAddr[13:0]};
                writeAddr36 = {writeAddr[13:0]};
                writeAddr35 = {writeAddr[13:0]};
                writeAddr34 = {writeAddr[13:0]};
                writeAddr33 = {writeAddr[13:0]};
                writeAddr32 = {writeAddr[13:0]};
                writeAddr31 = {writeAddr[13:0]};
                writeAddr30 = {writeAddr[13:0]};
                writeAddr29 = {writeAddr[13:0]};
                writeAddr28 = {writeAddr[13:0]};
                writeAddr27 = {writeAddr[13:0]};
                writeAddr26 = {writeAddr[13:0]};
                writeAddr25 = {writeAddr[13:0]};
                writeAddr24 = {writeAddr[13:0]};
                writeAddr23 = {writeAddr[13:0]};
                writeAddr22 = {writeAddr[13:0]};
                writeAddr21 = {writeAddr[13:0]};
                writeAddr20 = {writeAddr[13:0]};
                writeAddr19 = {writeAddr[13:0]};
                writeAddr18 = {writeAddr[12:0], 1'b0};
                writeAddr17 = {writeAddr[12:0], 1'b0};
                writeAddr16 = {writeAddr[12:0], 1'b0};
                writeAddr15 = {writeAddr[12:0], 1'b0};
                writeAddr14 = {writeAddr[12:0], 1'b0};
                writeAddr13 = {writeAddr[12:0], 1'b0};
                writeAddr12 = {writeAddr[12:0], 1'b0};
                writeAddr11 = {writeAddr[12:0], 1'b0};
                writeAddr10 = {writeAddr[12:0], 1'b0};
                writeAddr9 = {writeAddr[12:0], 1'b0};
                writeAddr8 = {writeAddr[12:0], 1'b0};
                writeAddr7 = {writeAddr[12:0], 1'b0};
                writeAddr6 = {writeAddr[12:0], 1'b0};
                writeAddr5 = {writeAddr[12:0], 1'b0};
                writeAddr4 = {writeAddr[12:0], 1'b0};
                writeAddr3 = {writeAddr[12:0], 1'b0};
                writeAddr2 = {writeAddr[9:0], 4'b0};
                writeAddr1 = {writeAddr[9:0], 4'b0};

                readAddr50 = {writeAddr[13:0]};
                readAddr49 = {writeAddr[13:0]};
                readAddr48 = {writeAddr[13:0]};
                readAddr47 = {writeAddr[13:0]};
                readAddr46 = {writeAddr[13:0]};
                readAddr45 = {writeAddr[13:0]};
                readAddr44 = {writeAddr[13:0]};
                readAddr43 = {writeAddr[13:0]};
                readAddr42 = {writeAddr[13:0]};
                readAddr41 = {writeAddr[13:0]};
                readAddr40 = {writeAddr[13:0]};
                readAddr39 = {writeAddr[13:0]};
                readAddr38 = {writeAddr[13:0]};
                readAddr37 = {writeAddr[13:0]};
                readAddr36 = {writeAddr[13:0]};
                readAddr35 = {writeAddr[13:0]};
                readAddr34 = {writeAddr[13:0]};
                readAddr33 = {writeAddr[13:0]};
                readAddr32 = {writeAddr[13:0]};
                readAddr31 = {writeAddr[13:0]};
                readAddr30 = {writeAddr[13:0]};
                readAddr29 = {writeAddr[13:0]};
                readAddr28 = {writeAddr[13:0]};
                readAddr27 = {writeAddr[13:0]};
                readAddr26 = {writeAddr[13:0]};
                readAddr25 = {writeAddr[13:0]};
                readAddr24 = {writeAddr[13:0]};
                readAddr23 = {writeAddr[13:0]};
                readAddr22 = {writeAddr[13:0]};
                readAddr21 = {writeAddr[13:0]};
                readAddr20 = {writeAddr[13:0]};
                readAddr19 = {writeAddr[13:0]};
                readAddr18  = {readAddr[12:0],  1'b0};
                readAddr17  = {readAddr[12:0],  1'b0};
                readAddr16  = {readAddr[12:0],  1'b0};
                readAddr15  = {readAddr[12:0],  1'b0};
                readAddr14  = {readAddr[12:0],  1'b0};
                readAddr13  = {readAddr[12:0],  1'b0};
                readAddr12  = {readAddr[12:0],  1'b0};
                readAddr11  = {readAddr[12:0],  1'b0};
                readAddr10  = {readAddr[12:0],  1'b0};
                readAddr9  = {readAddr[12:0],  1'b0};
                readAddr8  = {readAddr[12:0],  1'b0};
                readAddr7  = {readAddr[12:0],  1'b0};
                readAddr6  = {readAddr[12:0],  1'b0};
                readAddr5  = {readAddr[12:0],  1'b0};
                readAddr4  = {readAddr[12:0],  1'b0};
                readAddr3  = {readAddr[12:0],  1'b0};
                readAddr2  = {readAddr[9:0],  4'b0};
                readAddr1  = {readAddr[9:0],  4'b0};

                writeData50 = {17'b0, writeData[31]};
                writeData49 = {17'b0, writeData[30]};
                writeData48 = {17'b0, writeData[29]};
                writeData47 = {17'b0, writeData[28]};
                writeData46 = {17'b0, writeData[27]};
                writeData45 = {17'b0, writeData[26]};
                writeData44 = {17'b0, writeData[25]};
                writeData43 = {17'b0, writeData[24]};
                writeData42 = {17'b0, writeData[23]};
                writeData41 = {17'b0, writeData[22]};
                writeData40 = {17'b0, writeData[21]};
                writeData39 = {17'b0, writeData[20]};
                writeData38 = {17'b0, writeData[19]};
                writeData37 = {17'b0, writeData[18]};
                writeData36 = {17'b0, writeData[17]};
                writeData35 = {17'b0, writeData[16]};
                writeData34 = {17'b0, writeData[15]};
                writeData33 = {17'b0, writeData[14]};
                writeData32 = {17'b0, writeData[13]};
                writeData31 = {17'b0, writeData[12]};
                writeData30 = {17'b0, writeData[11]};
                writeData29 = {17'b0, writeData[10]};
                writeData28 = {17'b0, writeData[9]};
                writeData27 = {17'b0, writeData[8]};
                writeData26 = {17'b0, writeData[7]};
                writeData25 = {17'b0, writeData[6]};
                writeData24 = {17'b0, writeData[5]};
                writeData23 = {17'b0, writeData[4]};
                writeData22 = {17'b0, writeData[3]};
                writeData21 = {17'b0, writeData[2]};
                writeData20 = {17'b0, writeData[1]};
                writeData19 = {17'b0, writeData[0]};
                writeData18 = {16'b0, writeData[31:30]};
                writeData17 = {16'b0, writeData[29:28]};
                writeData16 = {16'b0, writeData[27:26]};
                writeData15 = {16'b0, writeData[25:24]};
                writeData14 = {16'b0, writeData[23:22]};
                writeData13 = {16'b0, writeData[21:20]};
                writeData12 = {16'b0, writeData[19:18]};
                writeData11 = {16'b0, writeData[17:16]};
                writeData10 = {16'b0, writeData[15:14]};
                writeData9 = {16'b0, writeData[13:12]};
                writeData8 = {16'b0, writeData[11:10]};
                writeData7 = {16'b0, writeData[9:8]};
                writeData6 = {16'b0, writeData[7:6]};
                writeData5 = {16'b0, writeData[5:4]};
                writeData4 = {16'b0, writeData[3:2]};
                writeData3 = {16'b0, writeData[1:0]};
                writeData2 = {1'b0, writeData[31:24], 1'b0, writeData[23:16]};
                writeData1 = {1'b0, writeData[15:8], 1'b0, writeData[7:0]};

                case (writeAddr[14:9])
                    6'b000000, 6'b000001, 6'b000010, 6'b000011,
                    6'b000100, 6'b000101, 6'b000110, 6'b000111,
                    6'b001000, 6'b001001, 6'b001010, 6'b001011,
                    6'b001100, 6'b001101, 6'b001110, 6'b001111,
                    6'b010000, 6'b010001, 6'b010010, 6'b010011,
                    6'b010100, 6'b010101, 6'b010110, 6'b010111,
                    6'b011000, 6'b011001, 6'b011010, 6'b011011,
                    6'b011100, 6'b011101, 6'b011110, 6'b011111 : begin
                        wen_a50 = {1'b0, wen};
                        wen_a49 = {1'b0, wen};
                        wen_a48 = {1'b0, wen};
                        wen_a47 = {1'b0, wen};
                        wen_a46 = {1'b0, wen};
                        wen_a45 = {1'b0, wen};
                        wen_a44 = {1'b0, wen};
                        wen_a43 = {1'b0, wen};
                        wen_a42 = {1'b0, wen};
                        wen_a41 = {1'b0, wen};
                        wen_a40 = {1'b0, wen};
                        wen_a39 = {1'b0, wen};
                        wen_a38 = {1'b0, wen};
                        wen_a37 = {1'b0, wen};
                        wen_a36 = {1'b0, wen};
                        wen_a35 = {1'b0, wen};
                        wen_a34 = {1'b0, wen};
                        wen_a33 = {1'b0, wen};
                        wen_a32 = {1'b0, wen};
                        wen_a31 = {1'b0, wen};
                        wen_a30 = {1'b0, wen};
                        wen_a29 = {1'b0, wen};
                        wen_a28 = {1'b0, wen};
                        wen_a27 = {1'b0, wen};
                        wen_a26 = {1'b0, wen};
                        wen_a25 = {1'b0, wen};
                        wen_a24 = {1'b0, wen};
                        wen_a23 = {1'b0, wen};
                        wen_a22 = {1'b0, wen};
                        wen_a21 = {1'b0, wen};
                        wen_a20 = {1'b0, wen};
                        wen_a19 = {1'b0, wen};
                        wen_a18 = {1'b0, 1'b0};
                        wen_a17 = {1'b0, 1'b0};
                        wen_a16 = {1'b0, 1'b0};
                        wen_a15 = {1'b0, 1'b0};
                        wen_a14 = {1'b0, 1'b0};
                        wen_a13 = {1'b0, 1'b0};
                        wen_a12 = {1'b0, 1'b0};
                        wen_a11 = {1'b0, 1'b0};
                        wen_a10 = {1'b0, 1'b0};
                        wen_a9 = {1'b0, 1'b0};
                        wen_a8 = {1'b0, 1'b0};
                        wen_a7 = {1'b0, 1'b0};
                        wen_a6 = {1'b0, 1'b0};
                        wen_a5 = {1'b0, 1'b0};
                        wen_a4 = {1'b0, 1'b0};
                        wen_a3 = {1'b0, 1'b0};
                        wen_a2 = {1'b0, 1'b0};
                        wen_a1 = {1'b0, 1'b0};
                    end
                    6'b100000, 6'b100001, 6'b100010, 6'b100011,
                    6'b100100, 6'b100101, 6'b100110, 6'b100111,
                    6'b101000, 6'b101001, 6'b101010, 6'b101011,
                    6'b101100, 6'b101101, 6'b101110, 6'b101111 : begin
                        wen_a50 = {1'b0, 1'b0};
                        wen_a49 = {1'b0, 1'b0};
                        wen_a48 = {1'b0, 1'b0};
                        wen_a47 = {1'b0, 1'b0};
                        wen_a46 = {1'b0, 1'b0};
                        wen_a45 = {1'b0, 1'b0};
                        wen_a44 = {1'b0, 1'b0};
                        wen_a43 = {1'b0, 1'b0};
                        wen_a42 = {1'b0, 1'b0};
                        wen_a41 = {1'b0, 1'b0};
                        wen_a40 = {1'b0, 1'b0};
                        wen_a39 = {1'b0, 1'b0};
                        wen_a38 = {1'b0, 1'b0};
                        wen_a37 = {1'b0, 1'b0};
                        wen_a36 = {1'b0, 1'b0};
                        wen_a35 = {1'b0, 1'b0};
                        wen_a34 = {1'b0, 1'b0};
                        wen_a33 = {1'b0, 1'b0};
                        wen_a32 = {1'b0, 1'b0};
                        wen_a31 = {1'b0, 1'b0};
                        wen_a30 = {1'b0, 1'b0};
                        wen_a29 = {1'b0, 1'b0};
                        wen_a28 = {1'b0, 1'b0};
                        wen_a27 = {1'b0, 1'b0};
                        wen_a26 = {1'b0, 1'b0};
                        wen_a25 = {1'b0, 1'b0};
                        wen_a24 = {1'b0, 1'b0};
                        wen_a23 = {1'b0, 1'b0};
                        wen_a22 = {1'b0, 1'b0};
                        wen_a21 = {1'b0, 1'b0};
                        wen_a20 = {1'b0, 1'b0};
                        wen_a19 = {1'b0, 1'b0};
                        wen_a18 = {1'b0, wen};
                        wen_a17 = {1'b0, wen};
                        wen_a16 = {1'b0, wen};
                        wen_a15 = {1'b0, wen};
                        wen_a14 = {1'b0, wen};
                        wen_a13 = {1'b0, wen};
                        wen_a12 = {1'b0, wen};
                        wen_a11 = {1'b0, wen};
                        wen_a10 = {1'b0, wen};
                        wen_a9 = {1'b0, wen};
                        wen_a8 = {1'b0, wen};
                        wen_a7 = {1'b0, wen};
                        wen_a6 = {1'b0, wen};
                        wen_a5 = {1'b0, wen};
                        wen_a4 = {1'b0, wen};
                        wen_a3 = {1'b0, wen};
                        wen_a2 = {1'b0, 1'b0};
                        wen_a1 = {1'b0, 1'b0};
                    end
                    6'b110000, 6'b110001 : begin
                        wen_a50 = {1'b0, 1'b0};
                        wen_a49 = {1'b0, 1'b0};
                        wen_a48 = {1'b0, 1'b0};
                        wen_a47 = {1'b0, 1'b0};
                        wen_a46 = {1'b0, 1'b0};
                        wen_a45 = {1'b0, 1'b0};
                        wen_a44 = {1'b0, 1'b0};
                        wen_a43 = {1'b0, 1'b0};
                        wen_a42 = {1'b0, 1'b0};
                        wen_a41 = {1'b0, 1'b0};
                        wen_a40 = {1'b0, 1'b0};
                        wen_a39 = {1'b0, 1'b0};
                        wen_a38 = {1'b0, 1'b0};
                        wen_a37 = {1'b0, 1'b0};
                        wen_a36 = {1'b0, 1'b0};
                        wen_a35 = {1'b0, 1'b0};
                        wen_a34 = {1'b0, 1'b0};
                        wen_a33 = {1'b0, 1'b0};
                        wen_a32 = {1'b0, 1'b0};
                        wen_a31 = {1'b0, 1'b0};
                        wen_a30 = {1'b0, 1'b0};
                        wen_a29 = {1'b0, 1'b0};
                        wen_a28 = {1'b0, 1'b0};
                        wen_a27 = {1'b0, 1'b0};
                        wen_a26 = {1'b0, 1'b0};
                        wen_a25 = {1'b0, 1'b0};
                        wen_a24 = {1'b0, 1'b0};
                        wen_a23 = {1'b0, 1'b0};
                        wen_a22 = {1'b0, 1'b0};
                        wen_a21 = {1'b0, 1'b0};
                        wen_a20 = {1'b0, 1'b0};
                        wen_a19 = {1'b0, 1'b0};
                        wen_a18 = {1'b0, 1'b0};
                        wen_a17 = {1'b0, 1'b0};
                        wen_a16 = {1'b0, 1'b0};
                        wen_a15 = {1'b0, 1'b0};
                        wen_a14 = {1'b0, 1'b0};
                        wen_a13 = {1'b0, 1'b0};
                        wen_a12 = {1'b0, 1'b0};
                        wen_a11 = {1'b0, 1'b0};
                        wen_a10 = {1'b0, 1'b0};
                        wen_a9 = {1'b0, 1'b0};
                        wen_a8 = {1'b0, 1'b0};
                        wen_a7 = {1'b0, 1'b0};
                        wen_a6 = {1'b0, 1'b0};
                        wen_a5 = {1'b0, 1'b0};
                        wen_a4 = {1'b0, 1'b0};
                        wen_a3 = {1'b0, 1'b0};
                        wen_a2 = {wen, wen};
                        wen_a1 = {wen, wen};
                    end
                    default : begin
                        wen_a50 = {1'b0, 1'b0};
                        wen_a49 = {1'b0, 1'b0};
                        wen_a48 = {1'b0, 1'b0};
                        wen_a47 = {1'b0, 1'b0};
                        wen_a46 = {1'b0, 1'b0};
                        wen_a45 = {1'b0, 1'b0};
                        wen_a44 = {1'b0, 1'b0};
                        wen_a43 = {1'b0, 1'b0};
                        wen_a42 = {1'b0, 1'b0};
                        wen_a41 = {1'b0, 1'b0};
                        wen_a40 = {1'b0, 1'b0};
                        wen_a39 = {1'b0, 1'b0};
                        wen_a38 = {1'b0, 1'b0};
                        wen_a37 = {1'b0, 1'b0};
                        wen_a36 = {1'b0, 1'b0};
                        wen_a35 = {1'b0, 1'b0};
                        wen_a34 = {1'b0, 1'b0};
                        wen_a33 = {1'b0, 1'b0};
                        wen_a32 = {1'b0, 1'b0};
                        wen_a31 = {1'b0, 1'b0};
                        wen_a30 = {1'b0, 1'b0};
                        wen_a29 = {1'b0, 1'b0};
                        wen_a28 = {1'b0, 1'b0};
                        wen_a27 = {1'b0, 1'b0};
                        wen_a26 = {1'b0, 1'b0};
                        wen_a25 = {1'b0, 1'b0};
                        wen_a24 = {1'b0, 1'b0};
                        wen_a23 = {1'b0, 1'b0};
                        wen_a22 = {1'b0, 1'b0};
                        wen_a21 = {1'b0, 1'b0};
                        wen_a20 = {1'b0, 1'b0};
                        wen_a19 = {1'b0, 1'b0};
                        wen_a18 = {1'b0, 1'b0};
                        wen_a17 = {1'b0, 1'b0};
                        wen_a16 = {1'b0, 1'b0};
                        wen_a15 = {1'b0, 1'b0};
                        wen_a14 = {1'b0, 1'b0};
                        wen_a13 = {1'b0, 1'b0};
                        wen_a12 = {1'b0, 1'b0};
                        wen_a11 = {1'b0, 1'b0};
                        wen_a10 = {1'b0, 1'b0};
                        wen_a9 = {1'b0, 1'b0};
                        wen_a8 = {1'b0, 1'b0};
                        wen_a7 = {1'b0, 1'b0};
                        wen_a6 = {1'b0, 1'b0};
                        wen_a5 = {1'b0, 1'b0};
                        wen_a4 = {1'b0, 1'b0};
                        wen_a3 = {1'b0, 1'b0};
                        wen_a2 = {1'b0, 1'b0};
                        wen_a1 = {1'b0, 1'b0};
                    end
                endcase

                case (ckRdAddr[14:9])
                    6'b000000, 6'b000001, 6'b000010, 6'b000011,
                    6'b000100, 6'b000101, 6'b000110, 6'b000111,
                    6'b001000, 6'b001001, 6'b001010, 6'b001011,
                    6'b001100, 6'b001101, 6'b001110, 6'b001111,
                    6'b010000, 6'b010001, 6'b010010, 6'b010011,
                    6'b010100, 6'b010101, 6'b010110, 6'b010111,
                    6'b011000, 6'b011001, 6'b011010, 6'b011011,
                    6'b011100, 6'b011101, 6'b011110, 6'b011111 : begin
                        readData = {
                                        readData50[0],
                                        readData49[0],
                                        readData48[0],
                                        readData47[0],
                                        readData46[0],
                                        readData45[0],
                                        readData44[0],
                                        readData43[0],
                                        readData42[0],
                                        readData41[0],
                                        readData40[0],
                                        readData39[0],
                                        readData38[0],
                                        readData37[0],
                                        readData36[0],
                                        readData35[0],
                                        readData34[0],
                                        readData33[0],
                                        readData32[0],
                                        readData31[0],
                                        readData30[0],
                                        readData29[0],
                                        readData28[0],
                                        readData27[0],
                                        readData26[0],
                                        readData25[0],
                                        readData24[0],
                                        readData23[0],
                                        readData22[0],
                                        readData21[0],
                                        readData20[0],
                                        readData19[0]
                        };
                    end
                    6'b100000, 6'b100001, 6'b100010, 6'b100011,
                    6'b100100, 6'b100101, 6'b100110, 6'b100111,
                    6'b101000, 6'b101001, 6'b101010, 6'b101011,
                    6'b101100, 6'b101101, 6'b101110, 6'b101111 : begin
                        readData = {
                                        readData18[1:0],
                                        readData17[1:0],
                                        readData16[1:0],
                                        readData15[1:0],
                                        readData14[1:0],
                                        readData13[1:0],
                                        readData12[1:0],
                                        readData11[1:0],
                                        readData10[1:0],
                                        readData9[1:0],
                                        readData8[1:0],
                                        readData7[1:0],
                                        readData6[1:0],
                                        readData5[1:0],
                                        readData4[1:0],
                                        readData3[1:0]
                        };
                    end
                    6'b110000, 6'b110001 : begin
                        readData = {readData2[16:9],readData2[7:0],readData1[16:9],readData1[7:0]};
                    end
                    default : begin
                        readData = 32'b0;
                    end
                endcase
            end        
            26112: begin
                width50 = 3'b000;
                width49 = 3'b000;
                width48 = 3'b000;
                width47 = 3'b000;
                width46 = 3'b000;
                width45 = 3'b000;
                width44 = 3'b000;
                width43 = 3'b000;
                width42 = 3'b000;
                width41 = 3'b000;
                width40 = 3'b000;
                width39 = 3'b000;
                width38 = 3'b000;
                width37 = 3'b000;
                width36 = 3'b000;
                width35 = 3'b000;
                width34 = 3'b000;
                width33 = 3'b000;
                width32 = 3'b000;
                width31 = 3'b000;
                width30 = 3'b000;
                width29 = 3'b000;
                width28 = 3'b000;
                width27 = 3'b000;
                width26 = 3'b000;
                width25 = 3'b000;
                width24 = 3'b000;
                width23 = 3'b000;
                width22 = 3'b000;
                width21 = 3'b000;
                width20 = 3'b000;
                width19 = 3'b000;
                width18 = 3'b001;
                width17 = 3'b001;
                width16 = 3'b001;
                width15 = 3'b001;
                width14 = 3'b001;
                width13 = 3'b001;
                width12 = 3'b001;
                width11 = 3'b001;
                width10 = 3'b001;
                width9 = 3'b001;
                width8 = 3'b001;
                width7 = 3'b001;
                width6 = 3'b001;
                width5 = 3'b001;
                width4 = 3'b001;
                width3 = 3'b001;
                width2 = 3'b100;
                width1 = 3'b100;
                width0 = 3'b101;

                writeAddr50 = {writeAddr[13:0]};
                writeAddr49 = {writeAddr[13:0]};
                writeAddr48 = {writeAddr[13:0]};
                writeAddr47 = {writeAddr[13:0]};
                writeAddr46 = {writeAddr[13:0]};
                writeAddr45 = {writeAddr[13:0]};
                writeAddr44 = {writeAddr[13:0]};
                writeAddr43 = {writeAddr[13:0]};
                writeAddr42 = {writeAddr[13:0]};
                writeAddr41 = {writeAddr[13:0]};
                writeAddr40 = {writeAddr[13:0]};
                writeAddr39 = {writeAddr[13:0]};
                writeAddr38 = {writeAddr[13:0]};
                writeAddr37 = {writeAddr[13:0]};
                writeAddr36 = {writeAddr[13:0]};
                writeAddr35 = {writeAddr[13:0]};
                writeAddr34 = {writeAddr[13:0]};
                writeAddr33 = {writeAddr[13:0]};
                writeAddr32 = {writeAddr[13:0]};
                writeAddr31 = {writeAddr[13:0]};
                writeAddr30 = {writeAddr[13:0]};
                writeAddr29 = {writeAddr[13:0]};
                writeAddr28 = {writeAddr[13:0]};
                writeAddr27 = {writeAddr[13:0]};
                writeAddr26 = {writeAddr[13:0]};
                writeAddr25 = {writeAddr[13:0]};
                writeAddr24 = {writeAddr[13:0]};
                writeAddr23 = {writeAddr[13:0]};
                writeAddr22 = {writeAddr[13:0]};
                writeAddr21 = {writeAddr[13:0]};
                writeAddr20 = {writeAddr[13:0]};
                writeAddr19 = {writeAddr[13:0]};
                writeAddr18 = {writeAddr[12:0], 1'b0};
                writeAddr17 = {writeAddr[12:0], 1'b0};
                writeAddr16 = {writeAddr[12:0], 1'b0};
                writeAddr15 = {writeAddr[12:0], 1'b0};
                writeAddr14 = {writeAddr[12:0], 1'b0};
                writeAddr13 = {writeAddr[12:0], 1'b0};
                writeAddr12 = {writeAddr[12:0], 1'b0};
                writeAddr11 = {writeAddr[12:0], 1'b0};
                writeAddr10 = {writeAddr[12:0], 1'b0};
                writeAddr9 = {writeAddr[12:0], 1'b0};
                writeAddr8 = {writeAddr[12:0], 1'b0};
                writeAddr7 = {writeAddr[12:0], 1'b0};
                writeAddr6 = {writeAddr[12:0], 1'b0};
                writeAddr5 = {writeAddr[12:0], 1'b0};
                writeAddr4 = {writeAddr[12:0], 1'b0};
                writeAddr3 = {writeAddr[12:0], 1'b0};
                writeAddr2 = {writeAddr[9:0], 4'b0};
                writeAddr1 = {writeAddr[9:0], 4'b0};
                writeAddr0 = {writeAddr[8:0], 5'b0};

                readAddr50 = {writeAddr[13:0]};
                readAddr49 = {writeAddr[13:0]};
                readAddr48 = {writeAddr[13:0]};
                readAddr47 = {writeAddr[13:0]};
                readAddr46 = {writeAddr[13:0]};
                readAddr45 = {writeAddr[13:0]};
                readAddr44 = {writeAddr[13:0]};
                readAddr43 = {writeAddr[13:0]};
                readAddr42 = {writeAddr[13:0]};
                readAddr41 = {writeAddr[13:0]};
                readAddr40 = {writeAddr[13:0]};
                readAddr39 = {writeAddr[13:0]};
                readAddr38 = {writeAddr[13:0]};
                readAddr37 = {writeAddr[13:0]};
                readAddr36 = {writeAddr[13:0]};
                readAddr35 = {writeAddr[13:0]};
                readAddr34 = {writeAddr[13:0]};
                readAddr33 = {writeAddr[13:0]};
                readAddr32 = {writeAddr[13:0]};
                readAddr31 = {writeAddr[13:0]};
                readAddr30 = {writeAddr[13:0]};
                readAddr29 = {writeAddr[13:0]};
                readAddr28 = {writeAddr[13:0]};
                readAddr27 = {writeAddr[13:0]};
                readAddr26 = {writeAddr[13:0]};
                readAddr25 = {writeAddr[13:0]};
                readAddr24 = {writeAddr[13:0]};
                readAddr23 = {writeAddr[13:0]};
                readAddr22 = {writeAddr[13:0]};
                readAddr21 = {writeAddr[13:0]};
                readAddr20 = {writeAddr[13:0]};
                readAddr19 = {writeAddr[13:0]};
                readAddr18  = {readAddr[12:0],  1'b0};
                readAddr17  = {readAddr[12:0],  1'b0};
                readAddr16  = {readAddr[12:0],  1'b0};
                readAddr15  = {readAddr[12:0],  1'b0};
                readAddr14  = {readAddr[12:0],  1'b0};
                readAddr13  = {readAddr[12:0],  1'b0};
                readAddr12  = {readAddr[12:0],  1'b0};
                readAddr11  = {readAddr[12:0],  1'b0};
                readAddr10  = {readAddr[12:0],  1'b0};
                readAddr9  = {readAddr[12:0],  1'b0};
                readAddr8  = {readAddr[12:0],  1'b0};
                readAddr7  = {readAddr[12:0],  1'b0};
                readAddr6  = {readAddr[12:0],  1'b0};
                readAddr5  = {readAddr[12:0],  1'b0};
                readAddr4  = {readAddr[12:0],  1'b0};
                readAddr3  = {readAddr[12:0],  1'b0};
                readAddr2  = {readAddr[9:0],  4'b0};
                readAddr1  = {readAddr[9:0],  4'b0};
                readAddr0  = {readAddr[8:0],  5'b0};

                writeData50 = {17'b0, writeData[31]};
                writeData49 = {17'b0, writeData[30]};
                writeData48 = {17'b0, writeData[29]};
                writeData47 = {17'b0, writeData[28]};
                writeData46 = {17'b0, writeData[27]};
                writeData45 = {17'b0, writeData[26]};
                writeData44 = {17'b0, writeData[25]};
                writeData43 = {17'b0, writeData[24]};
                writeData42 = {17'b0, writeData[23]};
                writeData41 = {17'b0, writeData[22]};
                writeData40 = {17'b0, writeData[21]};
                writeData39 = {17'b0, writeData[20]};
                writeData38 = {17'b0, writeData[19]};
                writeData37 = {17'b0, writeData[18]};
                writeData36 = {17'b0, writeData[17]};
                writeData35 = {17'b0, writeData[16]};
                writeData34 = {17'b0, writeData[15]};
                writeData33 = {17'b0, writeData[14]};
                writeData32 = {17'b0, writeData[13]};
                writeData31 = {17'b0, writeData[12]};
                writeData30 = {17'b0, writeData[11]};
                writeData29 = {17'b0, writeData[10]};
                writeData28 = {17'b0, writeData[9]};
                writeData27 = {17'b0, writeData[8]};
                writeData26 = {17'b0, writeData[7]};
                writeData25 = {17'b0, writeData[6]};
                writeData24 = {17'b0, writeData[5]};
                writeData23 = {17'b0, writeData[4]};
                writeData22 = {17'b0, writeData[3]};
                writeData21 = {17'b0, writeData[2]};
                writeData20 = {17'b0, writeData[1]};
                writeData19 = {17'b0, writeData[0]};
                writeData18 = {16'b0, writeData[31:30]};
                writeData17 = {16'b0, writeData[29:28]};
                writeData16 = {16'b0, writeData[27:26]};
                writeData15 = {16'b0, writeData[25:24]};
                writeData14 = {16'b0, writeData[23:22]};
                writeData13 = {16'b0, writeData[21:20]};
                writeData12 = {16'b0, writeData[19:18]};
                writeData11 = {16'b0, writeData[17:16]};
                writeData10 = {16'b0, writeData[15:14]};
                writeData9 = {16'b0, writeData[13:12]};
                writeData8 = {16'b0, writeData[11:10]};
                writeData7 = {16'b0, writeData[9:8]};
                writeData6 = {16'b0, writeData[7:6]};
                writeData5 = {16'b0, writeData[5:4]};
                writeData4 = {16'b0, writeData[3:2]};
                writeData3 = {16'b0, writeData[1:0]};
                writeData2 = {1'b0, writeData[31:24], 1'b0, writeData[23:16]};
                writeData1 = {1'b0, writeData[15:8], 1'b0, writeData[7:0]};
                writeData0 = {1'b0, writeData[31:24], 1'b0, writeData[23:16], 1'b0, writeData[15:8], 1'b0, writeData[7:0]};

                case (writeAddr[14:9])
                    6'b000000, 6'b000001, 6'b000010, 6'b000011,
                    6'b000100, 6'b000101, 6'b000110, 6'b000111,
                    6'b001000, 6'b001001, 6'b001010, 6'b001011,
                    6'b001100, 6'b001101, 6'b001110, 6'b001111,
                    6'b010000, 6'b010001, 6'b010010, 6'b010011,
                    6'b010100, 6'b010101, 6'b010110, 6'b010111,
                    6'b011000, 6'b011001, 6'b011010, 6'b011011,
                    6'b011100, 6'b011101, 6'b011110, 6'b011111 : begin
                        wen_a50 = {1'b0, wen};
                        wen_a49 = {1'b0, wen};
                        wen_a48 = {1'b0, wen};
                        wen_a47 = {1'b0, wen};
                        wen_a46 = {1'b0, wen};
                        wen_a45 = {1'b0, wen};
                        wen_a44 = {1'b0, wen};
                        wen_a43 = {1'b0, wen};
                        wen_a42 = {1'b0, wen};
                        wen_a41 = {1'b0, wen};
                        wen_a40 = {1'b0, wen};
                        wen_a39 = {1'b0, wen};
                        wen_a38 = {1'b0, wen};
                        wen_a37 = {1'b0, wen};
                        wen_a36 = {1'b0, wen};
                        wen_a35 = {1'b0, wen};
                        wen_a34 = {1'b0, wen};
                        wen_a33 = {1'b0, wen};
                        wen_a32 = {1'b0, wen};
                        wen_a31 = {1'b0, wen};
                        wen_a30 = {1'b0, wen};
                        wen_a29 = {1'b0, wen};
                        wen_a28 = {1'b0, wen};
                        wen_a27 = {1'b0, wen};
                        wen_a26 = {1'b0, wen};
                        wen_a25 = {1'b0, wen};
                        wen_a24 = {1'b0, wen};
                        wen_a23 = {1'b0, wen};
                        wen_a22 = {1'b0, wen};
                        wen_a21 = {1'b0, wen};
                        wen_a20 = {1'b0, wen};
                        wen_a19 = {1'b0, wen};
                        wen_a18 = {1'b0, 1'b0};
                        wen_a17 = {1'b0, 1'b0};
                        wen_a16 = {1'b0, 1'b0};
                        wen_a15 = {1'b0, 1'b0};
                        wen_a14 = {1'b0, 1'b0};
                        wen_a13 = {1'b0, 1'b0};
                        wen_a12 = {1'b0, 1'b0};
                        wen_a11 = {1'b0, 1'b0};
                        wen_a10 = {1'b0, 1'b0};
                        wen_a9 = {1'b0, 1'b0};
                        wen_a8 = {1'b0, 1'b0};
                        wen_a7 = {1'b0, 1'b0};
                        wen_a6 = {1'b0, 1'b0};
                        wen_a5 = {1'b0, 1'b0};
                        wen_a4 = {1'b0, 1'b0};
                        wen_a3 = {1'b0, 1'b0};
                        wen_a2 = {1'b0, 1'b0};
                        wen_a1 = {1'b0, 1'b0};
                        wen_a0 = {1'b0, 1'b0};
                        wen_b0 = {1'b0, 1'b0};
                    end
                    6'b100000, 6'b100001, 6'b100010, 6'b100011,
                    6'b100100, 6'b100101, 6'b100110, 6'b100111,
                    6'b101000, 6'b101001, 6'b101010, 6'b101011,
                    6'b101100, 6'b101101, 6'b101110, 6'b101111 : begin
                        wen_a50 = {1'b0, 1'b0};
                        wen_a49 = {1'b0, 1'b0};
                        wen_a48 = {1'b0, 1'b0};
                        wen_a47 = {1'b0, 1'b0};
                        wen_a46 = {1'b0, 1'b0};
                        wen_a45 = {1'b0, 1'b0};
                        wen_a44 = {1'b0, 1'b0};
                        wen_a43 = {1'b0, 1'b0};
                        wen_a42 = {1'b0, 1'b0};
                        wen_a41 = {1'b0, 1'b0};
                        wen_a40 = {1'b0, 1'b0};
                        wen_a39 = {1'b0, 1'b0};
                        wen_a38 = {1'b0, 1'b0};
                        wen_a37 = {1'b0, 1'b0};
                        wen_a36 = {1'b0, 1'b0};
                        wen_a35 = {1'b0, 1'b0};
                        wen_a34 = {1'b0, 1'b0};
                        wen_a33 = {1'b0, 1'b0};
                        wen_a32 = {1'b0, 1'b0};
                        wen_a31 = {1'b0, 1'b0};
                        wen_a30 = {1'b0, 1'b0};
                        wen_a29 = {1'b0, 1'b0};
                        wen_a28 = {1'b0, 1'b0};
                        wen_a27 = {1'b0, 1'b0};
                        wen_a26 = {1'b0, 1'b0};
                        wen_a25 = {1'b0, 1'b0};
                        wen_a24 = {1'b0, 1'b0};
                        wen_a23 = {1'b0, 1'b0};
                        wen_a22 = {1'b0, 1'b0};
                        wen_a21 = {1'b0, 1'b0};
                        wen_a20 = {1'b0, 1'b0};
                        wen_a19 = {1'b0, 1'b0};
                        wen_a18 = {1'b0, wen};
                        wen_a17 = {1'b0, wen};
                        wen_a16 = {1'b0, wen};
                        wen_a15 = {1'b0, wen};
                        wen_a14 = {1'b0, wen};
                        wen_a13 = {1'b0, wen};
                        wen_a12 = {1'b0, wen};
                        wen_a11 = {1'b0, wen};
                        wen_a10 = {1'b0, wen};
                        wen_a9 = {1'b0, wen};
                        wen_a8 = {1'b0, wen};
                        wen_a7 = {1'b0, wen};
                        wen_a6 = {1'b0, wen};
                        wen_a5 = {1'b0, wen};
                        wen_a4 = {1'b0, wen};
                        wen_a3 = {1'b0, wen};
                        wen_a2 = {1'b0, 1'b0};
                        wen_a1 = {1'b0, 1'b0};
                        wen_a0 = {1'b0, 1'b0};
                        wen_b0 = {1'b0, 1'b0};
                    end
                    6'b110000, 6'b110001 : begin
                        wen_a50 = {1'b0, 1'b0};
                        wen_a49 = {1'b0, 1'b0};
                        wen_a48 = {1'b0, 1'b0};
                        wen_a47 = {1'b0, 1'b0};
                        wen_a46 = {1'b0, 1'b0};
                        wen_a45 = {1'b0, 1'b0};
                        wen_a44 = {1'b0, 1'b0};
                        wen_a43 = {1'b0, 1'b0};
                        wen_a42 = {1'b0, 1'b0};
                        wen_a41 = {1'b0, 1'b0};
                        wen_a40 = {1'b0, 1'b0};
                        wen_a39 = {1'b0, 1'b0};
                        wen_a38 = {1'b0, 1'b0};
                        wen_a37 = {1'b0, 1'b0};
                        wen_a36 = {1'b0, 1'b0};
                        wen_a35 = {1'b0, 1'b0};
                        wen_a34 = {1'b0, 1'b0};
                        wen_a33 = {1'b0, 1'b0};
                        wen_a32 = {1'b0, 1'b0};
                        wen_a31 = {1'b0, 1'b0};
                        wen_a30 = {1'b0, 1'b0};
                        wen_a29 = {1'b0, 1'b0};
                        wen_a28 = {1'b0, 1'b0};
                        wen_a27 = {1'b0, 1'b0};
                        wen_a26 = {1'b0, 1'b0};
                        wen_a25 = {1'b0, 1'b0};
                        wen_a24 = {1'b0, 1'b0};
                        wen_a23 = {1'b0, 1'b0};
                        wen_a22 = {1'b0, 1'b0};
                        wen_a21 = {1'b0, 1'b0};
                        wen_a20 = {1'b0, 1'b0};
                        wen_a19 = {1'b0, 1'b0};
                        wen_a18 = {1'b0, 1'b0};
                        wen_a17 = {1'b0, 1'b0};
                        wen_a16 = {1'b0, 1'b0};
                        wen_a15 = {1'b0, 1'b0};
                        wen_a14 = {1'b0, 1'b0};
                        wen_a13 = {1'b0, 1'b0};
                        wen_a12 = {1'b0, 1'b0};
                        wen_a11 = {1'b0, 1'b0};
                        wen_a10 = {1'b0, 1'b0};
                        wen_a9 = {1'b0, 1'b0};
                        wen_a8 = {1'b0, 1'b0};
                        wen_a7 = {1'b0, 1'b0};
                        wen_a6 = {1'b0, 1'b0};
                        wen_a5 = {1'b0, 1'b0};
                        wen_a4 = {1'b0, 1'b0};
                        wen_a3 = {1'b0, 1'b0};
                        wen_a2 = {wen, wen};
                        wen_a1 = {wen, wen};
                        wen_a0 = {1'b0, 1'b0};
                        wen_b0 = {1'b0, 1'b0};
                    end
                    6'b110010 : begin
                        wen_a50 = {1'b0, 1'b0};
                        wen_a49 = {1'b0, 1'b0};
                        wen_a48 = {1'b0, 1'b0};
                        wen_a47 = {1'b0, 1'b0};
                        wen_a46 = {1'b0, 1'b0};
                        wen_a45 = {1'b0, 1'b0};
                        wen_a44 = {1'b0, 1'b0};
                        wen_a43 = {1'b0, 1'b0};
                        wen_a42 = {1'b0, 1'b0};
                        wen_a41 = {1'b0, 1'b0};
                        wen_a40 = {1'b0, 1'b0};
                        wen_a39 = {1'b0, 1'b0};
                        wen_a38 = {1'b0, 1'b0};
                        wen_a37 = {1'b0, 1'b0};
                        wen_a36 = {1'b0, 1'b0};
                        wen_a35 = {1'b0, 1'b0};
                        wen_a34 = {1'b0, 1'b0};
                        wen_a33 = {1'b0, 1'b0};
                        wen_a32 = {1'b0, 1'b0};
                        wen_a31 = {1'b0, 1'b0};
                        wen_a30 = {1'b0, 1'b0};
                        wen_a29 = {1'b0, 1'b0};
                        wen_a28 = {1'b0, 1'b0};
                        wen_a27 = {1'b0, 1'b0};
                        wen_a26 = {1'b0, 1'b0};
                        wen_a25 = {1'b0, 1'b0};
                        wen_a24 = {1'b0, 1'b0};
                        wen_a23 = {1'b0, 1'b0};
                        wen_a22 = {1'b0, 1'b0};
                        wen_a21 = {1'b0, 1'b0};
                        wen_a20 = {1'b0, 1'b0};
                        wen_a19 = {1'b0, 1'b0};
                        wen_a18 = {1'b0, 1'b0};
                        wen_a17 = {1'b0, 1'b0};
                        wen_a16 = {1'b0, 1'b0};
                        wen_a15 = {1'b0, 1'b0};
                        wen_a14 = {1'b0, 1'b0};
                        wen_a13 = {1'b0, 1'b0};
                        wen_a12 = {1'b0, 1'b0};
                        wen_a11 = {1'b0, 1'b0};
                        wen_a10 = {1'b0, 1'b0};
                        wen_a9 = {1'b0, 1'b0};
                        wen_a8 = {1'b0, 1'b0};
                        wen_a7 = {1'b0, 1'b0};
                        wen_a6 = {1'b0, 1'b0};
                        wen_a5 = {1'b0, 1'b0};
                        wen_a4 = {1'b0, 1'b0};
                        wen_a3 = {1'b0, 1'b0};
                        wen_a2 = {1'b0, 1'b0};
                        wen_a1 = {1'b0, 1'b0};
                        wen_a0 = {wen, wen};
                        wen_b0 = {wen, wen};
                    end
                    default : begin
                        wen_a50 = {1'b0, 1'b0};
                        wen_a49 = {1'b0, 1'b0};
                        wen_a48 = {1'b0, 1'b0};
                        wen_a47 = {1'b0, 1'b0};
                        wen_a46 = {1'b0, 1'b0};
                        wen_a45 = {1'b0, 1'b0};
                        wen_a44 = {1'b0, 1'b0};
                        wen_a43 = {1'b0, 1'b0};
                        wen_a42 = {1'b0, 1'b0};
                        wen_a41 = {1'b0, 1'b0};
                        wen_a40 = {1'b0, 1'b0};
                        wen_a39 = {1'b0, 1'b0};
                        wen_a38 = {1'b0, 1'b0};
                        wen_a37 = {1'b0, 1'b0};
                        wen_a36 = {1'b0, 1'b0};
                        wen_a35 = {1'b0, 1'b0};
                        wen_a34 = {1'b0, 1'b0};
                        wen_a33 = {1'b0, 1'b0};
                        wen_a32 = {1'b0, 1'b0};
                        wen_a31 = {1'b0, 1'b0};
                        wen_a30 = {1'b0, 1'b0};
                        wen_a29 = {1'b0, 1'b0};
                        wen_a28 = {1'b0, 1'b0};
                        wen_a27 = {1'b0, 1'b0};
                        wen_a26 = {1'b0, 1'b0};
                        wen_a25 = {1'b0, 1'b0};
                        wen_a24 = {1'b0, 1'b0};
                        wen_a23 = {1'b0, 1'b0};
                        wen_a22 = {1'b0, 1'b0};
                        wen_a21 = {1'b0, 1'b0};
                        wen_a20 = {1'b0, 1'b0};
                        wen_a19 = {1'b0, 1'b0};
                        wen_a18 = {1'b0, 1'b0};
                        wen_a17 = {1'b0, 1'b0};
                        wen_a16 = {1'b0, 1'b0};
                        wen_a15 = {1'b0, 1'b0};
                        wen_a14 = {1'b0, 1'b0};
                        wen_a13 = {1'b0, 1'b0};
                        wen_a12 = {1'b0, 1'b0};
                        wen_a11 = {1'b0, 1'b0};
                        wen_a10 = {1'b0, 1'b0};
                        wen_a9 = {1'b0, 1'b0};
                        wen_a8 = {1'b0, 1'b0};
                        wen_a7 = {1'b0, 1'b0};
                        wen_a6 = {1'b0, 1'b0};
                        wen_a5 = {1'b0, 1'b0};
                        wen_a4 = {1'b0, 1'b0};
                        wen_a3 = {1'b0, 1'b0};
                        wen_a2 = {1'b0, 1'b0};
                        wen_a1 = {1'b0, 1'b0};
                        wen_a0 = {1'b0, 1'b0};
                        wen_b0 = {1'b0, 1'b0};
                    end
                endcase

                case (ckRdAddr[14:9])
                    6'b000000, 6'b000001, 6'b000010, 6'b000011,
                    6'b000100, 6'b000101, 6'b000110, 6'b000111,
                    6'b001000, 6'b001001, 6'b001010, 6'b001011,
                    6'b001100, 6'b001101, 6'b001110, 6'b001111,
                    6'b010000, 6'b010001, 6'b010010, 6'b010011,
                    6'b010100, 6'b010101, 6'b010110, 6'b010111,
                    6'b011000, 6'b011001, 6'b011010, 6'b011011,
                    6'b011100, 6'b011101, 6'b011110, 6'b011111 : begin
                        readData = {
                                        readData50[0],
                                        readData49[0],
                                        readData48[0],
                                        readData47[0],
                                        readData46[0],
                                        readData45[0],
                                        readData44[0],
                                        readData43[0],
                                        readData42[0],
                                        readData41[0],
                                        readData40[0],
                                        readData39[0],
                                        readData38[0],
                                        readData37[0],
                                        readData36[0],
                                        readData35[0],
                                        readData34[0],
                                        readData33[0],
                                        readData32[0],
                                        readData31[0],
                                        readData30[0],
                                        readData29[0],
                                        readData28[0],
                                        readData27[0],
                                        readData26[0],
                                        readData25[0],
                                        readData24[0],
                                        readData23[0],
                                        readData22[0],
                                        readData21[0],
                                        readData20[0],
                                        readData19[0]
                        };
                    end
                    6'b100000, 6'b100001, 6'b100010, 6'b100011,
                    6'b100100, 6'b100101, 6'b100110, 6'b100111,
                    6'b101000, 6'b101001, 6'b101010, 6'b101011,
                    6'b101100, 6'b101101, 6'b101110, 6'b101111 : begin
                        readData = {
                                        readData18[1:0],
                                        readData17[1:0],
                                        readData16[1:0],
                                        readData15[1:0],
                                        readData14[1:0],
                                        readData13[1:0],
                                        readData12[1:0],
                                        readData11[1:0],
                                        readData10[1:0],
                                        readData9[1:0],
                                        readData8[1:0],
                                        readData7[1:0],
                                        readData6[1:0],
                                        readData5[1:0],
                                        readData4[1:0],
                                        readData3[1:0]
                        };
                    end
                    6'b110000, 6'b110001 : begin
                        readData = {readData2[16:9],readData2[7:0],readData1[16:9],readData1[7:0]};
                    end
                    6'b110010 : begin
                        readData = {readData0[34:27],readData0[25:18],readData0[16:9],readData0[7:0]};
                    end
                    default : begin
                        readData = 32'b0;
                    end
                endcase
            end        
            26624: begin
                width52 = 3'b000;
                width51 = 3'b000;
                width50 = 3'b000;
                width49 = 3'b000;
                width48 = 3'b000;
                width47 = 3'b000;
                width46 = 3'b000;
                width45 = 3'b000;
                width44 = 3'b000;
                width43 = 3'b000;
                width42 = 3'b000;
                width41 = 3'b000;
                width40 = 3'b000;
                width39 = 3'b000;
                width38 = 3'b000;
                width37 = 3'b000;
                width36 = 3'b000;
                width35 = 3'b000;
                width34 = 3'b000;
                width33 = 3'b000;
                width32 = 3'b000;
                width31 = 3'b000;
                width30 = 3'b000;
                width29 = 3'b000;
                width28 = 3'b000;
                width27 = 3'b000;
                width26 = 3'b000;
                width25 = 3'b000;
                width24 = 3'b000;
                width23 = 3'b000;
                width22 = 3'b000;
                width21 = 3'b000;
                width20 = 3'b001;
                width19 = 3'b001;
                width18 = 3'b001;
                width17 = 3'b001;
                width16 = 3'b001;
                width15 = 3'b001;
                width14 = 3'b001;
                width13 = 3'b001;
                width12 = 3'b001;
                width11 = 3'b001;
                width10 = 3'b001;
                width9 = 3'b001;
                width8 = 3'b001;
                width7 = 3'b001;
                width6 = 3'b001;
                width5 = 3'b001;
                width4 = 3'b011;
                width3 = 3'b011;
                width2 = 3'b011;
                width1 = 3'b011;

                writeAddr52 = {writeAddr[13:0]};
                writeAddr51 = {writeAddr[13:0]};
                writeAddr50 = {writeAddr[13:0]};
                writeAddr49 = {writeAddr[13:0]};
                writeAddr48 = {writeAddr[13:0]};
                writeAddr47 = {writeAddr[13:0]};
                writeAddr46 = {writeAddr[13:0]};
                writeAddr45 = {writeAddr[13:0]};
                writeAddr44 = {writeAddr[13:0]};
                writeAddr43 = {writeAddr[13:0]};
                writeAddr42 = {writeAddr[13:0]};
                writeAddr41 = {writeAddr[13:0]};
                writeAddr40 = {writeAddr[13:0]};
                writeAddr39 = {writeAddr[13:0]};
                writeAddr38 = {writeAddr[13:0]};
                writeAddr37 = {writeAddr[13:0]};
                writeAddr36 = {writeAddr[13:0]};
                writeAddr35 = {writeAddr[13:0]};
                writeAddr34 = {writeAddr[13:0]};
                writeAddr33 = {writeAddr[13:0]};
                writeAddr32 = {writeAddr[13:0]};
                writeAddr31 = {writeAddr[13:0]};
                writeAddr30 = {writeAddr[13:0]};
                writeAddr29 = {writeAddr[13:0]};
                writeAddr28 = {writeAddr[13:0]};
                writeAddr27 = {writeAddr[13:0]};
                writeAddr26 = {writeAddr[13:0]};
                writeAddr25 = {writeAddr[13:0]};
                writeAddr24 = {writeAddr[13:0]};
                writeAddr23 = {writeAddr[13:0]};
                writeAddr22 = {writeAddr[13:0]};
                writeAddr21 = {writeAddr[13:0]};
                writeAddr20 = {writeAddr[12:0], 1'b0};
                writeAddr19 = {writeAddr[12:0], 1'b0};
                writeAddr18 = {writeAddr[12:0], 1'b0};
                writeAddr17 = {writeAddr[12:0], 1'b0};
                writeAddr16 = {writeAddr[12:0], 1'b0};
                writeAddr15 = {writeAddr[12:0], 1'b0};
                writeAddr14 = {writeAddr[12:0], 1'b0};
                writeAddr13 = {writeAddr[12:0], 1'b0};
                writeAddr12 = {writeAddr[12:0], 1'b0};
                writeAddr11 = {writeAddr[12:0], 1'b0};
                writeAddr10 = {writeAddr[12:0], 1'b0};
                writeAddr9 = {writeAddr[12:0], 1'b0};
                writeAddr8 = {writeAddr[12:0], 1'b0};
                writeAddr7 = {writeAddr[12:0], 1'b0};
                writeAddr6 = {writeAddr[12:0], 1'b0};
                writeAddr5 = {writeAddr[12:0], 1'b0};
                writeAddr4 = {writeAddr[10:0], 3'b0};
                writeAddr3 = {writeAddr[10:0], 3'b0};
                writeAddr2 = {writeAddr[10:0], 3'b0};
                writeAddr1 = {writeAddr[10:0], 3'b0};

                readAddr52 = {writeAddr[13:0]};
                readAddr51 = {writeAddr[13:0]};
                readAddr50 = {writeAddr[13:0]};
                readAddr49 = {writeAddr[13:0]};
                readAddr48 = {writeAddr[13:0]};
                readAddr47 = {writeAddr[13:0]};
                readAddr46 = {writeAddr[13:0]};
                readAddr45 = {writeAddr[13:0]};
                readAddr44 = {writeAddr[13:0]};
                readAddr43 = {writeAddr[13:0]};
                readAddr42 = {writeAddr[13:0]};
                readAddr41 = {writeAddr[13:0]};
                readAddr40 = {writeAddr[13:0]};
                readAddr39 = {writeAddr[13:0]};
                readAddr38 = {writeAddr[13:0]};
                readAddr37 = {writeAddr[13:0]};
                readAddr36 = {writeAddr[13:0]};
                readAddr35 = {writeAddr[13:0]};
                readAddr34 = {writeAddr[13:0]};
                readAddr33 = {writeAddr[13:0]};
                readAddr32 = {writeAddr[13:0]};
                readAddr31 = {writeAddr[13:0]};
                readAddr30 = {writeAddr[13:0]};
                readAddr29 = {writeAddr[13:0]};
                readAddr28 = {writeAddr[13:0]};
                readAddr27 = {writeAddr[13:0]};
                readAddr26 = {writeAddr[13:0]};
                readAddr25 = {writeAddr[13:0]};
                readAddr24 = {writeAddr[13:0]};
                readAddr23 = {writeAddr[13:0]};
                readAddr22 = {writeAddr[13:0]};
                readAddr21 = {writeAddr[13:0]};
                readAddr20  = {readAddr[12:0],  1'b0};
                readAddr19  = {readAddr[12:0],  1'b0};
                readAddr18  = {readAddr[12:0],  1'b0};
                readAddr17  = {readAddr[12:0],  1'b0};
                readAddr16  = {readAddr[12:0],  1'b0};
                readAddr15  = {readAddr[12:0],  1'b0};
                readAddr14  = {readAddr[12:0],  1'b0};
                readAddr13  = {readAddr[12:0],  1'b0};
                readAddr12  = {readAddr[12:0],  1'b0};
                readAddr11  = {readAddr[12:0],  1'b0};
                readAddr10  = {readAddr[12:0],  1'b0};
                readAddr9  = {readAddr[12:0],  1'b0};
                readAddr8  = {readAddr[12:0],  1'b0};
                readAddr7  = {readAddr[12:0],  1'b0};
                readAddr6  = {readAddr[12:0],  1'b0};
                readAddr5  = {readAddr[12:0],  1'b0};
                readAddr4  = {readAddr[10:0],  3'b0};
                readAddr3  = {readAddr[10:0],  3'b0};
                readAddr2  = {readAddr[10:0],  3'b0};
                readAddr1  = {readAddr[10:0],  3'b0};

                writeData52 = {17'b0, writeData[31]};
                writeData51 = {17'b0, writeData[30]};
                writeData50 = {17'b0, writeData[29]};
                writeData49 = {17'b0, writeData[28]};
                writeData48 = {17'b0, writeData[27]};
                writeData47 = {17'b0, writeData[26]};
                writeData46 = {17'b0, writeData[25]};
                writeData45 = {17'b0, writeData[24]};
                writeData44 = {17'b0, writeData[23]};
                writeData43 = {17'b0, writeData[22]};
                writeData42 = {17'b0, writeData[21]};
                writeData41 = {17'b0, writeData[20]};
                writeData40 = {17'b0, writeData[19]};
                writeData39 = {17'b0, writeData[18]};
                writeData38 = {17'b0, writeData[17]};
                writeData37 = {17'b0, writeData[16]};
                writeData36 = {17'b0, writeData[15]};
                writeData35 = {17'b0, writeData[14]};
                writeData34 = {17'b0, writeData[13]};
                writeData33 = {17'b0, writeData[12]};
                writeData32 = {17'b0, writeData[11]};
                writeData31 = {17'b0, writeData[10]};
                writeData30 = {17'b0, writeData[9]};
                writeData29 = {17'b0, writeData[8]};
                writeData28 = {17'b0, writeData[7]};
                writeData27 = {17'b0, writeData[6]};
                writeData26 = {17'b0, writeData[5]};
                writeData25 = {17'b0, writeData[4]};
                writeData24 = {17'b0, writeData[3]};
                writeData23 = {17'b0, writeData[2]};
                writeData22 = {17'b0, writeData[1]};
                writeData21 = {17'b0, writeData[0]};
                writeData20 = {16'b0, writeData[31:30]};
                writeData19 = {16'b0, writeData[29:28]};
                writeData18 = {16'b0, writeData[27:26]};
                writeData17 = {16'b0, writeData[25:24]};
                writeData16 = {16'b0, writeData[23:22]};
                writeData15 = {16'b0, writeData[21:20]};
                writeData14 = {16'b0, writeData[19:18]};
                writeData13 = {16'b0, writeData[17:16]};
                writeData12 = {16'b0, writeData[15:14]};
                writeData11 = {16'b0, writeData[13:12]};
                writeData10 = {16'b0, writeData[11:10]};
                writeData9 = {16'b0, writeData[9:8]};
                writeData8 = {16'b0, writeData[7:6]};
                writeData7 = {16'b0, writeData[5:4]};
                writeData6 = {16'b0, writeData[3:2]};
                writeData5 = {16'b0, writeData[1:0]};
                writeData4 = {10'b0, writeData[31:24]};
                writeData3 = {10'b0, writeData[23:16]};
                writeData2 = {10'b0, writeData[15:8]};
                writeData1 = {10'b0, writeData[7:0]};

                case (writeAddr[14:9])
                    6'b000000, 6'b000001, 6'b000010, 6'b000011,
                    6'b000100, 6'b000101, 6'b000110, 6'b000111,
                    6'b001000, 6'b001001, 6'b001010, 6'b001011,
                    6'b001100, 6'b001101, 6'b001110, 6'b001111,
                    6'b010000, 6'b010001, 6'b010010, 6'b010011,
                    6'b010100, 6'b010101, 6'b010110, 6'b010111,
                    6'b011000, 6'b011001, 6'b011010, 6'b011011,
                    6'b011100, 6'b011101, 6'b011110, 6'b011111 : begin
                        wen_a52 = {1'b0, wen};
                        wen_a51 = {1'b0, wen};
                        wen_a50 = {1'b0, wen};
                        wen_a49 = {1'b0, wen};
                        wen_a48 = {1'b0, wen};
                        wen_a47 = {1'b0, wen};
                        wen_a46 = {1'b0, wen};
                        wen_a45 = {1'b0, wen};
                        wen_a44 = {1'b0, wen};
                        wen_a43 = {1'b0, wen};
                        wen_a42 = {1'b0, wen};
                        wen_a41 = {1'b0, wen};
                        wen_a40 = {1'b0, wen};
                        wen_a39 = {1'b0, wen};
                        wen_a38 = {1'b0, wen};
                        wen_a37 = {1'b0, wen};
                        wen_a36 = {1'b0, wen};
                        wen_a35 = {1'b0, wen};
                        wen_a34 = {1'b0, wen};
                        wen_a33 = {1'b0, wen};
                        wen_a32 = {1'b0, wen};
                        wen_a31 = {1'b0, wen};
                        wen_a30 = {1'b0, wen};
                        wen_a29 = {1'b0, wen};
                        wen_a28 = {1'b0, wen};
                        wen_a27 = {1'b0, wen};
                        wen_a26 = {1'b0, wen};
                        wen_a25 = {1'b0, wen};
                        wen_a24 = {1'b0, wen};
                        wen_a23 = {1'b0, wen};
                        wen_a22 = {1'b0, wen};
                        wen_a21 = {1'b0, wen};
                        wen_a20 = {1'b0, 1'b0};
                        wen_a19 = {1'b0, 1'b0};
                        wen_a18 = {1'b0, 1'b0};
                        wen_a17 = {1'b0, 1'b0};
                        wen_a16 = {1'b0, 1'b0};
                        wen_a15 = {1'b0, 1'b0};
                        wen_a14 = {1'b0, 1'b0};
                        wen_a13 = {1'b0, 1'b0};
                        wen_a12 = {1'b0, 1'b0};
                        wen_a11 = {1'b0, 1'b0};
                        wen_a10 = {1'b0, 1'b0};
                        wen_a9 = {1'b0, 1'b0};
                        wen_a8 = {1'b0, 1'b0};
                        wen_a7 = {1'b0, 1'b0};
                        wen_a6 = {1'b0, 1'b0};
                        wen_a5 = {1'b0, 1'b0};
                        wen_a4 = {1'b0, 1'b0};
                        wen_a3 = {1'b0, 1'b0};
                        wen_a2 = {1'b0, 1'b0};
                        wen_a1 = {1'b0, 1'b0};
                    end
                    6'b100000, 6'b100001, 6'b100010, 6'b100011,
                    6'b100100, 6'b100101, 6'b100110, 6'b100111,
                    6'b101000, 6'b101001, 6'b101010, 6'b101011,
                    6'b101100, 6'b101101, 6'b101110, 6'b101111 : begin
                        wen_a52 = {1'b0, 1'b0};
                        wen_a51 = {1'b0, 1'b0};
                        wen_a50 = {1'b0, 1'b0};
                        wen_a49 = {1'b0, 1'b0};
                        wen_a48 = {1'b0, 1'b0};
                        wen_a47 = {1'b0, 1'b0};
                        wen_a46 = {1'b0, 1'b0};
                        wen_a45 = {1'b0, 1'b0};
                        wen_a44 = {1'b0, 1'b0};
                        wen_a43 = {1'b0, 1'b0};
                        wen_a42 = {1'b0, 1'b0};
                        wen_a41 = {1'b0, 1'b0};
                        wen_a40 = {1'b0, 1'b0};
                        wen_a39 = {1'b0, 1'b0};
                        wen_a38 = {1'b0, 1'b0};
                        wen_a37 = {1'b0, 1'b0};
                        wen_a36 = {1'b0, 1'b0};
                        wen_a35 = {1'b0, 1'b0};
                        wen_a34 = {1'b0, 1'b0};
                        wen_a33 = {1'b0, 1'b0};
                        wen_a32 = {1'b0, 1'b0};
                        wen_a31 = {1'b0, 1'b0};
                        wen_a30 = {1'b0, 1'b0};
                        wen_a29 = {1'b0, 1'b0};
                        wen_a28 = {1'b0, 1'b0};
                        wen_a27 = {1'b0, 1'b0};
                        wen_a26 = {1'b0, 1'b0};
                        wen_a25 = {1'b0, 1'b0};
                        wen_a24 = {1'b0, 1'b0};
                        wen_a23 = {1'b0, 1'b0};
                        wen_a22 = {1'b0, 1'b0};
                        wen_a21 = {1'b0, 1'b0};
                        wen_a20 = {1'b0, wen};
                        wen_a19 = {1'b0, wen};
                        wen_a18 = {1'b0, wen};
                        wen_a17 = {1'b0, wen};
                        wen_a16 = {1'b0, wen};
                        wen_a15 = {1'b0, wen};
                        wen_a14 = {1'b0, wen};
                        wen_a13 = {1'b0, wen};
                        wen_a12 = {1'b0, wen};
                        wen_a11 = {1'b0, wen};
                        wen_a10 = {1'b0, wen};
                        wen_a9 = {1'b0, wen};
                        wen_a8 = {1'b0, wen};
                        wen_a7 = {1'b0, wen};
                        wen_a6 = {1'b0, wen};
                        wen_a5 = {1'b0, wen};
                        wen_a4 = {1'b0, 1'b0};
                        wen_a3 = {1'b0, 1'b0};
                        wen_a2 = {1'b0, 1'b0};
                        wen_a1 = {1'b0, 1'b0};
                    end
                    6'b110000, 6'b110001, 6'b110010, 6'b110011 : begin
                        wen_a52 = {1'b0, 1'b0};
                        wen_a51 = {1'b0, 1'b0};
                        wen_a50 = {1'b0, 1'b0};
                        wen_a49 = {1'b0, 1'b0};
                        wen_a48 = {1'b0, 1'b0};
                        wen_a47 = {1'b0, 1'b0};
                        wen_a46 = {1'b0, 1'b0};
                        wen_a45 = {1'b0, 1'b0};
                        wen_a44 = {1'b0, 1'b0};
                        wen_a43 = {1'b0, 1'b0};
                        wen_a42 = {1'b0, 1'b0};
                        wen_a41 = {1'b0, 1'b0};
                        wen_a40 = {1'b0, 1'b0};
                        wen_a39 = {1'b0, 1'b0};
                        wen_a38 = {1'b0, 1'b0};
                        wen_a37 = {1'b0, 1'b0};
                        wen_a36 = {1'b0, 1'b0};
                        wen_a35 = {1'b0, 1'b0};
                        wen_a34 = {1'b0, 1'b0};
                        wen_a33 = {1'b0, 1'b0};
                        wen_a32 = {1'b0, 1'b0};
                        wen_a31 = {1'b0, 1'b0};
                        wen_a30 = {1'b0, 1'b0};
                        wen_a29 = {1'b0, 1'b0};
                        wen_a28 = {1'b0, 1'b0};
                        wen_a27 = {1'b0, 1'b0};
                        wen_a26 = {1'b0, 1'b0};
                        wen_a25 = {1'b0, 1'b0};
                        wen_a24 = {1'b0, 1'b0};
                        wen_a23 = {1'b0, 1'b0};
                        wen_a22 = {1'b0, 1'b0};
                        wen_a21 = {1'b0, 1'b0};
                        wen_a20 = {1'b0, 1'b0};
                        wen_a19 = {1'b0, 1'b0};
                        wen_a18 = {1'b0, 1'b0};
                        wen_a17 = {1'b0, 1'b0};
                        wen_a16 = {1'b0, 1'b0};
                        wen_a15 = {1'b0, 1'b0};
                        wen_a14 = {1'b0, 1'b0};
                        wen_a13 = {1'b0, 1'b0};
                        wen_a12 = {1'b0, 1'b0};
                        wen_a11 = {1'b0, 1'b0};
                        wen_a10 = {1'b0, 1'b0};
                        wen_a9 = {1'b0, 1'b0};
                        wen_a8 = {1'b0, 1'b0};
                        wen_a7 = {1'b0, 1'b0};
                        wen_a6 = {1'b0, 1'b0};
                        wen_a5 = {1'b0, 1'b0};
                        wen_a4 = {1'b0, wen};
                        wen_a3 = {1'b0, wen};
                        wen_a2 = {1'b0, wen};
                        wen_a1 = {1'b0, wen};
                    end
                    default : begin
                        wen_a52 = {1'b0, 1'b0};
                        wen_a51 = {1'b0, 1'b0};
                        wen_a50 = {1'b0, 1'b0};
                        wen_a49 = {1'b0, 1'b0};
                        wen_a48 = {1'b0, 1'b0};
                        wen_a47 = {1'b0, 1'b0};
                        wen_a46 = {1'b0, 1'b0};
                        wen_a45 = {1'b0, 1'b0};
                        wen_a44 = {1'b0, 1'b0};
                        wen_a43 = {1'b0, 1'b0};
                        wen_a42 = {1'b0, 1'b0};
                        wen_a41 = {1'b0, 1'b0};
                        wen_a40 = {1'b0, 1'b0};
                        wen_a39 = {1'b0, 1'b0};
                        wen_a38 = {1'b0, 1'b0};
                        wen_a37 = {1'b0, 1'b0};
                        wen_a36 = {1'b0, 1'b0};
                        wen_a35 = {1'b0, 1'b0};
                        wen_a34 = {1'b0, 1'b0};
                        wen_a33 = {1'b0, 1'b0};
                        wen_a32 = {1'b0, 1'b0};
                        wen_a31 = {1'b0, 1'b0};
                        wen_a30 = {1'b0, 1'b0};
                        wen_a29 = {1'b0, 1'b0};
                        wen_a28 = {1'b0, 1'b0};
                        wen_a27 = {1'b0, 1'b0};
                        wen_a26 = {1'b0, 1'b0};
                        wen_a25 = {1'b0, 1'b0};
                        wen_a24 = {1'b0, 1'b0};
                        wen_a23 = {1'b0, 1'b0};
                        wen_a22 = {1'b0, 1'b0};
                        wen_a21 = {1'b0, 1'b0};
                        wen_a20 = {1'b0, 1'b0};
                        wen_a19 = {1'b0, 1'b0};
                        wen_a18 = {1'b0, 1'b0};
                        wen_a17 = {1'b0, 1'b0};
                        wen_a16 = {1'b0, 1'b0};
                        wen_a15 = {1'b0, 1'b0};
                        wen_a14 = {1'b0, 1'b0};
                        wen_a13 = {1'b0, 1'b0};
                        wen_a12 = {1'b0, 1'b0};
                        wen_a11 = {1'b0, 1'b0};
                        wen_a10 = {1'b0, 1'b0};
                        wen_a9 = {1'b0, 1'b0};
                        wen_a8 = {1'b0, 1'b0};
                        wen_a7 = {1'b0, 1'b0};
                        wen_a6 = {1'b0, 1'b0};
                        wen_a5 = {1'b0, 1'b0};
                        wen_a4 = {1'b0, 1'b0};
                        wen_a3 = {1'b0, 1'b0};
                        wen_a2 = {1'b0, 1'b0};
                        wen_a1 = {1'b0, 1'b0};
                    end
                endcase

                case (ckRdAddr[14:9])
                    6'b000000, 6'b000001, 6'b000010, 6'b000011,
                    6'b000100, 6'b000101, 6'b000110, 6'b000111,
                    6'b001000, 6'b001001, 6'b001010, 6'b001011,
                    6'b001100, 6'b001101, 6'b001110, 6'b001111,
                    6'b010000, 6'b010001, 6'b010010, 6'b010011,
                    6'b010100, 6'b010101, 6'b010110, 6'b010111,
                    6'b011000, 6'b011001, 6'b011010, 6'b011011,
                    6'b011100, 6'b011101, 6'b011110, 6'b011111 : begin
                        readData = {
                                        readData52[0],
                                        readData51[0],
                                        readData50[0],
                                        readData49[0],
                                        readData48[0],
                                        readData47[0],
                                        readData46[0],
                                        readData45[0],
                                        readData44[0],
                                        readData43[0],
                                        readData42[0],
                                        readData41[0],
                                        readData40[0],
                                        readData39[0],
                                        readData38[0],
                                        readData37[0],
                                        readData36[0],
                                        readData35[0],
                                        readData34[0],
                                        readData33[0],
                                        readData32[0],
                                        readData31[0],
                                        readData30[0],
                                        readData29[0],
                                        readData28[0],
                                        readData27[0],
                                        readData26[0],
                                        readData25[0],
                                        readData24[0],
                                        readData23[0],
                                        readData22[0],
                                        readData21[0]
                        };
                    end
                    6'b100000, 6'b100001, 6'b100010, 6'b100011,
                    6'b100100, 6'b100101, 6'b100110, 6'b100111,
                    6'b101000, 6'b101001, 6'b101010, 6'b101011,
                    6'b101100, 6'b101101, 6'b101110, 6'b101111 : begin
                        readData = {
                                        readData20[1:0],
                                        readData19[1:0],
                                        readData18[1:0],
                                        readData17[1:0],
                                        readData16[1:0],
                                        readData15[1:0],
                                        readData14[1:0],
                                        readData13[1:0],
                                        readData12[1:0],
                                        readData11[1:0],
                                        readData10[1:0],
                                        readData9[1:0],
                                        readData8[1:0],
                                        readData7[1:0],
                                        readData6[1:0],
                                        readData5[1:0]
                        };
                    end
                    6'b110000, 6'b110001, 6'b110010, 6'b110011 : begin
                        readData = {readData4[7:0],readData3[7:0],readData2[7:0],readData1[7:0]};
                    end
                    default : begin
                        readData = 32'b0;
                    end
                endcase
            end        
            27136: begin
                width52 = 3'b000;
                width51 = 3'b000;
                width50 = 3'b000;
                width49 = 3'b000;
                width48 = 3'b000;
                width47 = 3'b000;
                width46 = 3'b000;
                width45 = 3'b000;
                width44 = 3'b000;
                width43 = 3'b000;
                width42 = 3'b000;
                width41 = 3'b000;
                width40 = 3'b000;
                width39 = 3'b000;
                width38 = 3'b000;
                width37 = 3'b000;
                width36 = 3'b000;
                width35 = 3'b000;
                width34 = 3'b000;
                width33 = 3'b000;
                width32 = 3'b000;
                width31 = 3'b000;
                width30 = 3'b000;
                width29 = 3'b000;
                width28 = 3'b000;
                width27 = 3'b000;
                width26 = 3'b000;
                width25 = 3'b000;
                width24 = 3'b000;
                width23 = 3'b000;
                width22 = 3'b000;
                width21 = 3'b000;
                width20 = 3'b001;
                width19 = 3'b001;
                width18 = 3'b001;
                width17 = 3'b001;
                width16 = 3'b001;
                width15 = 3'b001;
                width14 = 3'b001;
                width13 = 3'b001;
                width12 = 3'b001;
                width11 = 3'b001;
                width10 = 3'b001;
                width9 = 3'b001;
                width8 = 3'b001;
                width7 = 3'b001;
                width6 = 3'b001;
                width5 = 3'b001;
                width4 = 3'b011;
                width3 = 3'b011;
                width2 = 3'b011;
                width1 = 3'b011;
                width0 = 3'b101;

                writeAddr52 = {writeAddr[13:0]};
                writeAddr51 = {writeAddr[13:0]};
                writeAddr50 = {writeAddr[13:0]};
                writeAddr49 = {writeAddr[13:0]};
                writeAddr48 = {writeAddr[13:0]};
                writeAddr47 = {writeAddr[13:0]};
                writeAddr46 = {writeAddr[13:0]};
                writeAddr45 = {writeAddr[13:0]};
                writeAddr44 = {writeAddr[13:0]};
                writeAddr43 = {writeAddr[13:0]};
                writeAddr42 = {writeAddr[13:0]};
                writeAddr41 = {writeAddr[13:0]};
                writeAddr40 = {writeAddr[13:0]};
                writeAddr39 = {writeAddr[13:0]};
                writeAddr38 = {writeAddr[13:0]};
                writeAddr37 = {writeAddr[13:0]};
                writeAddr36 = {writeAddr[13:0]};
                writeAddr35 = {writeAddr[13:0]};
                writeAddr34 = {writeAddr[13:0]};
                writeAddr33 = {writeAddr[13:0]};
                writeAddr32 = {writeAddr[13:0]};
                writeAddr31 = {writeAddr[13:0]};
                writeAddr30 = {writeAddr[13:0]};
                writeAddr29 = {writeAddr[13:0]};
                writeAddr28 = {writeAddr[13:0]};
                writeAddr27 = {writeAddr[13:0]};
                writeAddr26 = {writeAddr[13:0]};
                writeAddr25 = {writeAddr[13:0]};
                writeAddr24 = {writeAddr[13:0]};
                writeAddr23 = {writeAddr[13:0]};
                writeAddr22 = {writeAddr[13:0]};
                writeAddr21 = {writeAddr[13:0]};
                writeAddr20 = {writeAddr[12:0], 1'b0};
                writeAddr19 = {writeAddr[12:0], 1'b0};
                writeAddr18 = {writeAddr[12:0], 1'b0};
                writeAddr17 = {writeAddr[12:0], 1'b0};
                writeAddr16 = {writeAddr[12:0], 1'b0};
                writeAddr15 = {writeAddr[12:0], 1'b0};
                writeAddr14 = {writeAddr[12:0], 1'b0};
                writeAddr13 = {writeAddr[12:0], 1'b0};
                writeAddr12 = {writeAddr[12:0], 1'b0};
                writeAddr11 = {writeAddr[12:0], 1'b0};
                writeAddr10 = {writeAddr[12:0], 1'b0};
                writeAddr9 = {writeAddr[12:0], 1'b0};
                writeAddr8 = {writeAddr[12:0], 1'b0};
                writeAddr7 = {writeAddr[12:0], 1'b0};
                writeAddr6 = {writeAddr[12:0], 1'b0};
                writeAddr5 = {writeAddr[12:0], 1'b0};
                writeAddr4 = {writeAddr[10:0], 3'b0};
                writeAddr3 = {writeAddr[10:0], 3'b0};
                writeAddr2 = {writeAddr[10:0], 3'b0};
                writeAddr1 = {writeAddr[10:0], 3'b0};
                writeAddr0 = {writeAddr[8:0], 5'b0};

                readAddr52 = {writeAddr[13:0]};
                readAddr51 = {writeAddr[13:0]};
                readAddr50 = {writeAddr[13:0]};
                readAddr49 = {writeAddr[13:0]};
                readAddr48 = {writeAddr[13:0]};
                readAddr47 = {writeAddr[13:0]};
                readAddr46 = {writeAddr[13:0]};
                readAddr45 = {writeAddr[13:0]};
                readAddr44 = {writeAddr[13:0]};
                readAddr43 = {writeAddr[13:0]};
                readAddr42 = {writeAddr[13:0]};
                readAddr41 = {writeAddr[13:0]};
                readAddr40 = {writeAddr[13:0]};
                readAddr39 = {writeAddr[13:0]};
                readAddr38 = {writeAddr[13:0]};
                readAddr37 = {writeAddr[13:0]};
                readAddr36 = {writeAddr[13:0]};
                readAddr35 = {writeAddr[13:0]};
                readAddr34 = {writeAddr[13:0]};
                readAddr33 = {writeAddr[13:0]};
                readAddr32 = {writeAddr[13:0]};
                readAddr31 = {writeAddr[13:0]};
                readAddr30 = {writeAddr[13:0]};
                readAddr29 = {writeAddr[13:0]};
                readAddr28 = {writeAddr[13:0]};
                readAddr27 = {writeAddr[13:0]};
                readAddr26 = {writeAddr[13:0]};
                readAddr25 = {writeAddr[13:0]};
                readAddr24 = {writeAddr[13:0]};
                readAddr23 = {writeAddr[13:0]};
                readAddr22 = {writeAddr[13:0]};
                readAddr21 = {writeAddr[13:0]};
                readAddr20  = {readAddr[12:0],  1'b0};
                readAddr19  = {readAddr[12:0],  1'b0};
                readAddr18  = {readAddr[12:0],  1'b0};
                readAddr17  = {readAddr[12:0],  1'b0};
                readAddr16  = {readAddr[12:0],  1'b0};
                readAddr15  = {readAddr[12:0],  1'b0};
                readAddr14  = {readAddr[12:0],  1'b0};
                readAddr13  = {readAddr[12:0],  1'b0};
                readAddr12  = {readAddr[12:0],  1'b0};
                readAddr11  = {readAddr[12:0],  1'b0};
                readAddr10  = {readAddr[12:0],  1'b0};
                readAddr9  = {readAddr[12:0],  1'b0};
                readAddr8  = {readAddr[12:0],  1'b0};
                readAddr7  = {readAddr[12:0],  1'b0};
                readAddr6  = {readAddr[12:0],  1'b0};
                readAddr5  = {readAddr[12:0],  1'b0};
                readAddr4  = {readAddr[10:0],  3'b0};
                readAddr3  = {readAddr[10:0],  3'b0};
                readAddr2  = {readAddr[10:0],  3'b0};
                readAddr1  = {readAddr[10:0],  3'b0};
                readAddr0  = {readAddr[8:0],  5'b0};

                writeData52 = {17'b0, writeData[31]};
                writeData51 = {17'b0, writeData[30]};
                writeData50 = {17'b0, writeData[29]};
                writeData49 = {17'b0, writeData[28]};
                writeData48 = {17'b0, writeData[27]};
                writeData47 = {17'b0, writeData[26]};
                writeData46 = {17'b0, writeData[25]};
                writeData45 = {17'b0, writeData[24]};
                writeData44 = {17'b0, writeData[23]};
                writeData43 = {17'b0, writeData[22]};
                writeData42 = {17'b0, writeData[21]};
                writeData41 = {17'b0, writeData[20]};
                writeData40 = {17'b0, writeData[19]};
                writeData39 = {17'b0, writeData[18]};
                writeData38 = {17'b0, writeData[17]};
                writeData37 = {17'b0, writeData[16]};
                writeData36 = {17'b0, writeData[15]};
                writeData35 = {17'b0, writeData[14]};
                writeData34 = {17'b0, writeData[13]};
                writeData33 = {17'b0, writeData[12]};
                writeData32 = {17'b0, writeData[11]};
                writeData31 = {17'b0, writeData[10]};
                writeData30 = {17'b0, writeData[9]};
                writeData29 = {17'b0, writeData[8]};
                writeData28 = {17'b0, writeData[7]};
                writeData27 = {17'b0, writeData[6]};
                writeData26 = {17'b0, writeData[5]};
                writeData25 = {17'b0, writeData[4]};
                writeData24 = {17'b0, writeData[3]};
                writeData23 = {17'b0, writeData[2]};
                writeData22 = {17'b0, writeData[1]};
                writeData21 = {17'b0, writeData[0]};
                writeData20 = {16'b0, writeData[31:30]};
                writeData19 = {16'b0, writeData[29:28]};
                writeData18 = {16'b0, writeData[27:26]};
                writeData17 = {16'b0, writeData[25:24]};
                writeData16 = {16'b0, writeData[23:22]};
                writeData15 = {16'b0, writeData[21:20]};
                writeData14 = {16'b0, writeData[19:18]};
                writeData13 = {16'b0, writeData[17:16]};
                writeData12 = {16'b0, writeData[15:14]};
                writeData11 = {16'b0, writeData[13:12]};
                writeData10 = {16'b0, writeData[11:10]};
                writeData9 = {16'b0, writeData[9:8]};
                writeData8 = {16'b0, writeData[7:6]};
                writeData7 = {16'b0, writeData[5:4]};
                writeData6 = {16'b0, writeData[3:2]};
                writeData5 = {16'b0, writeData[1:0]};
                writeData4 = {10'b0, writeData[31:24]};
                writeData3 = {10'b0, writeData[23:16]};
                writeData2 = {10'b0, writeData[15:8]};
                writeData1 = {10'b0, writeData[7:0]};
                writeData0 = {1'b0, writeData[31:24], 1'b0, writeData[23:16], 1'b0, writeData[15:8], 1'b0, writeData[7:0]};

                case (writeAddr[14:9])
                    6'b000000, 6'b000001, 6'b000010, 6'b000011,
                    6'b000100, 6'b000101, 6'b000110, 6'b000111,
                    6'b001000, 6'b001001, 6'b001010, 6'b001011,
                    6'b001100, 6'b001101, 6'b001110, 6'b001111,
                    6'b010000, 6'b010001, 6'b010010, 6'b010011,
                    6'b010100, 6'b010101, 6'b010110, 6'b010111,
                    6'b011000, 6'b011001, 6'b011010, 6'b011011,
                    6'b011100, 6'b011101, 6'b011110, 6'b011111 : begin
                        wen_a52 = {1'b0, wen};
                        wen_a51 = {1'b0, wen};
                        wen_a50 = {1'b0, wen};
                        wen_a49 = {1'b0, wen};
                        wen_a48 = {1'b0, wen};
                        wen_a47 = {1'b0, wen};
                        wen_a46 = {1'b0, wen};
                        wen_a45 = {1'b0, wen};
                        wen_a44 = {1'b0, wen};
                        wen_a43 = {1'b0, wen};
                        wen_a42 = {1'b0, wen};
                        wen_a41 = {1'b0, wen};
                        wen_a40 = {1'b0, wen};
                        wen_a39 = {1'b0, wen};
                        wen_a38 = {1'b0, wen};
                        wen_a37 = {1'b0, wen};
                        wen_a36 = {1'b0, wen};
                        wen_a35 = {1'b0, wen};
                        wen_a34 = {1'b0, wen};
                        wen_a33 = {1'b0, wen};
                        wen_a32 = {1'b0, wen};
                        wen_a31 = {1'b0, wen};
                        wen_a30 = {1'b0, wen};
                        wen_a29 = {1'b0, wen};
                        wen_a28 = {1'b0, wen};
                        wen_a27 = {1'b0, wen};
                        wen_a26 = {1'b0, wen};
                        wen_a25 = {1'b0, wen};
                        wen_a24 = {1'b0, wen};
                        wen_a23 = {1'b0, wen};
                        wen_a22 = {1'b0, wen};
                        wen_a21 = {1'b0, wen};
                        wen_a20 = {1'b0, 1'b0};
                        wen_a19 = {1'b0, 1'b0};
                        wen_a18 = {1'b0, 1'b0};
                        wen_a17 = {1'b0, 1'b0};
                        wen_a16 = {1'b0, 1'b0};
                        wen_a15 = {1'b0, 1'b0};
                        wen_a14 = {1'b0, 1'b0};
                        wen_a13 = {1'b0, 1'b0};
                        wen_a12 = {1'b0, 1'b0};
                        wen_a11 = {1'b0, 1'b0};
                        wen_a10 = {1'b0, 1'b0};
                        wen_a9 = {1'b0, 1'b0};
                        wen_a8 = {1'b0, 1'b0};
                        wen_a7 = {1'b0, 1'b0};
                        wen_a6 = {1'b0, 1'b0};
                        wen_a5 = {1'b0, 1'b0};
                        wen_a4 = {1'b0, 1'b0};
                        wen_a3 = {1'b0, 1'b0};
                        wen_a2 = {1'b0, 1'b0};
                        wen_a1 = {1'b0, 1'b0};
                        wen_a0 = {1'b0, 1'b0};
                        wen_b0 = {1'b0, 1'b0};
                    end
                    6'b100000, 6'b100001, 6'b100010, 6'b100011,
                    6'b100100, 6'b100101, 6'b100110, 6'b100111,
                    6'b101000, 6'b101001, 6'b101010, 6'b101011,
                    6'b101100, 6'b101101, 6'b101110, 6'b101111 : begin
                        wen_a52 = {1'b0, 1'b0};
                        wen_a51 = {1'b0, 1'b0};
                        wen_a50 = {1'b0, 1'b0};
                        wen_a49 = {1'b0, 1'b0};
                        wen_a48 = {1'b0, 1'b0};
                        wen_a47 = {1'b0, 1'b0};
                        wen_a46 = {1'b0, 1'b0};
                        wen_a45 = {1'b0, 1'b0};
                        wen_a44 = {1'b0, 1'b0};
                        wen_a43 = {1'b0, 1'b0};
                        wen_a42 = {1'b0, 1'b0};
                        wen_a41 = {1'b0, 1'b0};
                        wen_a40 = {1'b0, 1'b0};
                        wen_a39 = {1'b0, 1'b0};
                        wen_a38 = {1'b0, 1'b0};
                        wen_a37 = {1'b0, 1'b0};
                        wen_a36 = {1'b0, 1'b0};
                        wen_a35 = {1'b0, 1'b0};
                        wen_a34 = {1'b0, 1'b0};
                        wen_a33 = {1'b0, 1'b0};
                        wen_a32 = {1'b0, 1'b0};
                        wen_a31 = {1'b0, 1'b0};
                        wen_a30 = {1'b0, 1'b0};
                        wen_a29 = {1'b0, 1'b0};
                        wen_a28 = {1'b0, 1'b0};
                        wen_a27 = {1'b0, 1'b0};
                        wen_a26 = {1'b0, 1'b0};
                        wen_a25 = {1'b0, 1'b0};
                        wen_a24 = {1'b0, 1'b0};
                        wen_a23 = {1'b0, 1'b0};
                        wen_a22 = {1'b0, 1'b0};
                        wen_a21 = {1'b0, 1'b0};
                        wen_a20 = {1'b0, wen};
                        wen_a19 = {1'b0, wen};
                        wen_a18 = {1'b0, wen};
                        wen_a17 = {1'b0, wen};
                        wen_a16 = {1'b0, wen};
                        wen_a15 = {1'b0, wen};
                        wen_a14 = {1'b0, wen};
                        wen_a13 = {1'b0, wen};
                        wen_a12 = {1'b0, wen};
                        wen_a11 = {1'b0, wen};
                        wen_a10 = {1'b0, wen};
                        wen_a9 = {1'b0, wen};
                        wen_a8 = {1'b0, wen};
                        wen_a7 = {1'b0, wen};
                        wen_a6 = {1'b0, wen};
                        wen_a5 = {1'b0, wen};
                        wen_a4 = {1'b0, 1'b0};
                        wen_a3 = {1'b0, 1'b0};
                        wen_a2 = {1'b0, 1'b0};
                        wen_a1 = {1'b0, 1'b0};
                        wen_a0 = {1'b0, 1'b0};
                        wen_b0 = {1'b0, 1'b0};
                    end
                    6'b110000, 6'b110001, 6'b110010, 6'b110011 : begin
                        wen_a52 = {1'b0, 1'b0};
                        wen_a51 = {1'b0, 1'b0};
                        wen_a50 = {1'b0, 1'b0};
                        wen_a49 = {1'b0, 1'b0};
                        wen_a48 = {1'b0, 1'b0};
                        wen_a47 = {1'b0, 1'b0};
                        wen_a46 = {1'b0, 1'b0};
                        wen_a45 = {1'b0, 1'b0};
                        wen_a44 = {1'b0, 1'b0};
                        wen_a43 = {1'b0, 1'b0};
                        wen_a42 = {1'b0, 1'b0};
                        wen_a41 = {1'b0, 1'b0};
                        wen_a40 = {1'b0, 1'b0};
                        wen_a39 = {1'b0, 1'b0};
                        wen_a38 = {1'b0, 1'b0};
                        wen_a37 = {1'b0, 1'b0};
                        wen_a36 = {1'b0, 1'b0};
                        wen_a35 = {1'b0, 1'b0};
                        wen_a34 = {1'b0, 1'b0};
                        wen_a33 = {1'b0, 1'b0};
                        wen_a32 = {1'b0, 1'b0};
                        wen_a31 = {1'b0, 1'b0};
                        wen_a30 = {1'b0, 1'b0};
                        wen_a29 = {1'b0, 1'b0};
                        wen_a28 = {1'b0, 1'b0};
                        wen_a27 = {1'b0, 1'b0};
                        wen_a26 = {1'b0, 1'b0};
                        wen_a25 = {1'b0, 1'b0};
                        wen_a24 = {1'b0, 1'b0};
                        wen_a23 = {1'b0, 1'b0};
                        wen_a22 = {1'b0, 1'b0};
                        wen_a21 = {1'b0, 1'b0};
                        wen_a20 = {1'b0, 1'b0};
                        wen_a19 = {1'b0, 1'b0};
                        wen_a18 = {1'b0, 1'b0};
                        wen_a17 = {1'b0, 1'b0};
                        wen_a16 = {1'b0, 1'b0};
                        wen_a15 = {1'b0, 1'b0};
                        wen_a14 = {1'b0, 1'b0};
                        wen_a13 = {1'b0, 1'b0};
                        wen_a12 = {1'b0, 1'b0};
                        wen_a11 = {1'b0, 1'b0};
                        wen_a10 = {1'b0, 1'b0};
                        wen_a9 = {1'b0, 1'b0};
                        wen_a8 = {1'b0, 1'b0};
                        wen_a7 = {1'b0, 1'b0};
                        wen_a6 = {1'b0, 1'b0};
                        wen_a5 = {1'b0, 1'b0};
                        wen_a4 = {1'b0, wen};
                        wen_a3 = {1'b0, wen};
                        wen_a2 = {1'b0, wen};
                        wen_a1 = {1'b0, wen};
                        wen_a0 = {1'b0, 1'b0};
                        wen_b0 = {1'b0, 1'b0};
                    end
                    6'b110100 : begin
                        wen_a52 = {1'b0, 1'b0};
                        wen_a51 = {1'b0, 1'b0};
                        wen_a50 = {1'b0, 1'b0};
                        wen_a49 = {1'b0, 1'b0};
                        wen_a48 = {1'b0, 1'b0};
                        wen_a47 = {1'b0, 1'b0};
                        wen_a46 = {1'b0, 1'b0};
                        wen_a45 = {1'b0, 1'b0};
                        wen_a44 = {1'b0, 1'b0};
                        wen_a43 = {1'b0, 1'b0};
                        wen_a42 = {1'b0, 1'b0};
                        wen_a41 = {1'b0, 1'b0};
                        wen_a40 = {1'b0, 1'b0};
                        wen_a39 = {1'b0, 1'b0};
                        wen_a38 = {1'b0, 1'b0};
                        wen_a37 = {1'b0, 1'b0};
                        wen_a36 = {1'b0, 1'b0};
                        wen_a35 = {1'b0, 1'b0};
                        wen_a34 = {1'b0, 1'b0};
                        wen_a33 = {1'b0, 1'b0};
                        wen_a32 = {1'b0, 1'b0};
                        wen_a31 = {1'b0, 1'b0};
                        wen_a30 = {1'b0, 1'b0};
                        wen_a29 = {1'b0, 1'b0};
                        wen_a28 = {1'b0, 1'b0};
                        wen_a27 = {1'b0, 1'b0};
                        wen_a26 = {1'b0, 1'b0};
                        wen_a25 = {1'b0, 1'b0};
                        wen_a24 = {1'b0, 1'b0};
                        wen_a23 = {1'b0, 1'b0};
                        wen_a22 = {1'b0, 1'b0};
                        wen_a21 = {1'b0, 1'b0};
                        wen_a20 = {1'b0, 1'b0};
                        wen_a19 = {1'b0, 1'b0};
                        wen_a18 = {1'b0, 1'b0};
                        wen_a17 = {1'b0, 1'b0};
                        wen_a16 = {1'b0, 1'b0};
                        wen_a15 = {1'b0, 1'b0};
                        wen_a14 = {1'b0, 1'b0};
                        wen_a13 = {1'b0, 1'b0};
                        wen_a12 = {1'b0, 1'b0};
                        wen_a11 = {1'b0, 1'b0};
                        wen_a10 = {1'b0, 1'b0};
                        wen_a9 = {1'b0, 1'b0};
                        wen_a8 = {1'b0, 1'b0};
                        wen_a7 = {1'b0, 1'b0};
                        wen_a6 = {1'b0, 1'b0};
                        wen_a5 = {1'b0, 1'b0};
                        wen_a4 = {1'b0, 1'b0};
                        wen_a3 = {1'b0, 1'b0};
                        wen_a2 = {1'b0, 1'b0};
                        wen_a1 = {1'b0, 1'b0};
                        wen_a0 = {wen, wen};
                        wen_b0 = {wen, wen};
                    end
                    default : begin
                        wen_a52 = {1'b0, 1'b0};
                        wen_a51 = {1'b0, 1'b0};
                        wen_a50 = {1'b0, 1'b0};
                        wen_a49 = {1'b0, 1'b0};
                        wen_a48 = {1'b0, 1'b0};
                        wen_a47 = {1'b0, 1'b0};
                        wen_a46 = {1'b0, 1'b0};
                        wen_a45 = {1'b0, 1'b0};
                        wen_a44 = {1'b0, 1'b0};
                        wen_a43 = {1'b0, 1'b0};
                        wen_a42 = {1'b0, 1'b0};
                        wen_a41 = {1'b0, 1'b0};
                        wen_a40 = {1'b0, 1'b0};
                        wen_a39 = {1'b0, 1'b0};
                        wen_a38 = {1'b0, 1'b0};
                        wen_a37 = {1'b0, 1'b0};
                        wen_a36 = {1'b0, 1'b0};
                        wen_a35 = {1'b0, 1'b0};
                        wen_a34 = {1'b0, 1'b0};
                        wen_a33 = {1'b0, 1'b0};
                        wen_a32 = {1'b0, 1'b0};
                        wen_a31 = {1'b0, 1'b0};
                        wen_a30 = {1'b0, 1'b0};
                        wen_a29 = {1'b0, 1'b0};
                        wen_a28 = {1'b0, 1'b0};
                        wen_a27 = {1'b0, 1'b0};
                        wen_a26 = {1'b0, 1'b0};
                        wen_a25 = {1'b0, 1'b0};
                        wen_a24 = {1'b0, 1'b0};
                        wen_a23 = {1'b0, 1'b0};
                        wen_a22 = {1'b0, 1'b0};
                        wen_a21 = {1'b0, 1'b0};
                        wen_a20 = {1'b0, 1'b0};
                        wen_a19 = {1'b0, 1'b0};
                        wen_a18 = {1'b0, 1'b0};
                        wen_a17 = {1'b0, 1'b0};
                        wen_a16 = {1'b0, 1'b0};
                        wen_a15 = {1'b0, 1'b0};
                        wen_a14 = {1'b0, 1'b0};
                        wen_a13 = {1'b0, 1'b0};
                        wen_a12 = {1'b0, 1'b0};
                        wen_a11 = {1'b0, 1'b0};
                        wen_a10 = {1'b0, 1'b0};
                        wen_a9 = {1'b0, 1'b0};
                        wen_a8 = {1'b0, 1'b0};
                        wen_a7 = {1'b0, 1'b0};
                        wen_a6 = {1'b0, 1'b0};
                        wen_a5 = {1'b0, 1'b0};
                        wen_a4 = {1'b0, 1'b0};
                        wen_a3 = {1'b0, 1'b0};
                        wen_a2 = {1'b0, 1'b0};
                        wen_a1 = {1'b0, 1'b0};
                        wen_a0 = {1'b0, 1'b0};
                        wen_b0 = {1'b0, 1'b0};
                    end
                endcase

                case (ckRdAddr[14:9])
                    6'b000000, 6'b000001, 6'b000010, 6'b000011,
                    6'b000100, 6'b000101, 6'b000110, 6'b000111,
                    6'b001000, 6'b001001, 6'b001010, 6'b001011,
                    6'b001100, 6'b001101, 6'b001110, 6'b001111,
                    6'b010000, 6'b010001, 6'b010010, 6'b010011,
                    6'b010100, 6'b010101, 6'b010110, 6'b010111,
                    6'b011000, 6'b011001, 6'b011010, 6'b011011,
                    6'b011100, 6'b011101, 6'b011110, 6'b011111 : begin
                        readData = {
                                        readData52[0],
                                        readData51[0],
                                        readData50[0],
                                        readData49[0],
                                        readData48[0],
                                        readData47[0],
                                        readData46[0],
                                        readData45[0],
                                        readData44[0],
                                        readData43[0],
                                        readData42[0],
                                        readData41[0],
                                        readData40[0],
                                        readData39[0],
                                        readData38[0],
                                        readData37[0],
                                        readData36[0],
                                        readData35[0],
                                        readData34[0],
                                        readData33[0],
                                        readData32[0],
                                        readData31[0],
                                        readData30[0],
                                        readData29[0],
                                        readData28[0],
                                        readData27[0],
                                        readData26[0],
                                        readData25[0],
                                        readData24[0],
                                        readData23[0],
                                        readData22[0],
                                        readData21[0]
                        };
                    end
                    6'b100000, 6'b100001, 6'b100010, 6'b100011,
                    6'b100100, 6'b100101, 6'b100110, 6'b100111,
                    6'b101000, 6'b101001, 6'b101010, 6'b101011,
                    6'b101100, 6'b101101, 6'b101110, 6'b101111 : begin
                        readData = {
                                        readData20[1:0],
                                        readData19[1:0],
                                        readData18[1:0],
                                        readData17[1:0],
                                        readData16[1:0],
                                        readData15[1:0],
                                        readData14[1:0],
                                        readData13[1:0],
                                        readData12[1:0],
                                        readData11[1:0],
                                        readData10[1:0],
                                        readData9[1:0],
                                        readData8[1:0],
                                        readData7[1:0],
                                        readData6[1:0],
                                        readData5[1:0]
                        };
                    end
                    6'b110000, 6'b110001, 6'b110010, 6'b110011 : begin
                        readData = {readData4[7:0],readData3[7:0],readData2[7:0],readData1[7:0]};
                    end
                    6'b110100 : begin
                        readData = {readData0[34:27],readData0[25:18],readData0[16:9],readData0[7:0]};
                    end
                    default : begin
                        readData = 32'b0;
                    end
                endcase
            end        
            27648: begin
                width54 = 3'b000;
                width53 = 3'b000;
                width52 = 3'b000;
                width51 = 3'b000;
                width50 = 3'b000;
                width49 = 3'b000;
                width48 = 3'b000;
                width47 = 3'b000;
                width46 = 3'b000;
                width45 = 3'b000;
                width44 = 3'b000;
                width43 = 3'b000;
                width42 = 3'b000;
                width41 = 3'b000;
                width40 = 3'b000;
                width39 = 3'b000;
                width38 = 3'b000;
                width37 = 3'b000;
                width36 = 3'b000;
                width35 = 3'b000;
                width34 = 3'b000;
                width33 = 3'b000;
                width32 = 3'b000;
                width31 = 3'b000;
                width30 = 3'b000;
                width29 = 3'b000;
                width28 = 3'b000;
                width27 = 3'b000;
                width26 = 3'b000;
                width25 = 3'b000;
                width24 = 3'b000;
                width23 = 3'b000;
                width22 = 3'b001;
                width21 = 3'b001;
                width20 = 3'b001;
                width19 = 3'b001;
                width18 = 3'b001;
                width17 = 3'b001;
                width16 = 3'b001;
                width15 = 3'b001;
                width14 = 3'b001;
                width13 = 3'b001;
                width12 = 3'b001;
                width11 = 3'b001;
                width10 = 3'b001;
                width9 = 3'b001;
                width8 = 3'b001;
                width7 = 3'b001;
                width6 = 3'b011;
                width5 = 3'b011;
                width4 = 3'b011;
                width3 = 3'b011;
                width2 = 3'b100;
                width1 = 3'b100;

                writeAddr54 = {writeAddr[13:0]};
                writeAddr53 = {writeAddr[13:0]};
                writeAddr52 = {writeAddr[13:0]};
                writeAddr51 = {writeAddr[13:0]};
                writeAddr50 = {writeAddr[13:0]};
                writeAddr49 = {writeAddr[13:0]};
                writeAddr48 = {writeAddr[13:0]};
                writeAddr47 = {writeAddr[13:0]};
                writeAddr46 = {writeAddr[13:0]};
                writeAddr45 = {writeAddr[13:0]};
                writeAddr44 = {writeAddr[13:0]};
                writeAddr43 = {writeAddr[13:0]};
                writeAddr42 = {writeAddr[13:0]};
                writeAddr41 = {writeAddr[13:0]};
                writeAddr40 = {writeAddr[13:0]};
                writeAddr39 = {writeAddr[13:0]};
                writeAddr38 = {writeAddr[13:0]};
                writeAddr37 = {writeAddr[13:0]};
                writeAddr36 = {writeAddr[13:0]};
                writeAddr35 = {writeAddr[13:0]};
                writeAddr34 = {writeAddr[13:0]};
                writeAddr33 = {writeAddr[13:0]};
                writeAddr32 = {writeAddr[13:0]};
                writeAddr31 = {writeAddr[13:0]};
                writeAddr30 = {writeAddr[13:0]};
                writeAddr29 = {writeAddr[13:0]};
                writeAddr28 = {writeAddr[13:0]};
                writeAddr27 = {writeAddr[13:0]};
                writeAddr26 = {writeAddr[13:0]};
                writeAddr25 = {writeAddr[13:0]};
                writeAddr24 = {writeAddr[13:0]};
                writeAddr23 = {writeAddr[13:0]};
                writeAddr22 = {writeAddr[12:0], 1'b0};
                writeAddr21 = {writeAddr[12:0], 1'b0};
                writeAddr20 = {writeAddr[12:0], 1'b0};
                writeAddr19 = {writeAddr[12:0], 1'b0};
                writeAddr18 = {writeAddr[12:0], 1'b0};
                writeAddr17 = {writeAddr[12:0], 1'b0};
                writeAddr16 = {writeAddr[12:0], 1'b0};
                writeAddr15 = {writeAddr[12:0], 1'b0};
                writeAddr14 = {writeAddr[12:0], 1'b0};
                writeAddr13 = {writeAddr[12:0], 1'b0};
                writeAddr12 = {writeAddr[12:0], 1'b0};
                writeAddr11 = {writeAddr[12:0], 1'b0};
                writeAddr10 = {writeAddr[12:0], 1'b0};
                writeAddr9 = {writeAddr[12:0], 1'b0};
                writeAddr8 = {writeAddr[12:0], 1'b0};
                writeAddr7 = {writeAddr[12:0], 1'b0};
                writeAddr6 = {writeAddr[10:0], 3'b0};
                writeAddr5 = {writeAddr[10:0], 3'b0};
                writeAddr4 = {writeAddr[10:0], 3'b0};
                writeAddr3 = {writeAddr[10:0], 3'b0};
                writeAddr2 = {writeAddr[9:0], 4'b0};
                writeAddr1 = {writeAddr[9:0], 4'b0};

                readAddr54 = {writeAddr[13:0]};
                readAddr53 = {writeAddr[13:0]};
                readAddr52 = {writeAddr[13:0]};
                readAddr51 = {writeAddr[13:0]};
                readAddr50 = {writeAddr[13:0]};
                readAddr49 = {writeAddr[13:0]};
                readAddr48 = {writeAddr[13:0]};
                readAddr47 = {writeAddr[13:0]};
                readAddr46 = {writeAddr[13:0]};
                readAddr45 = {writeAddr[13:0]};
                readAddr44 = {writeAddr[13:0]};
                readAddr43 = {writeAddr[13:0]};
                readAddr42 = {writeAddr[13:0]};
                readAddr41 = {writeAddr[13:0]};
                readAddr40 = {writeAddr[13:0]};
                readAddr39 = {writeAddr[13:0]};
                readAddr38 = {writeAddr[13:0]};
                readAddr37 = {writeAddr[13:0]};
                readAddr36 = {writeAddr[13:0]};
                readAddr35 = {writeAddr[13:0]};
                readAddr34 = {writeAddr[13:0]};
                readAddr33 = {writeAddr[13:0]};
                readAddr32 = {writeAddr[13:0]};
                readAddr31 = {writeAddr[13:0]};
                readAddr30 = {writeAddr[13:0]};
                readAddr29 = {writeAddr[13:0]};
                readAddr28 = {writeAddr[13:0]};
                readAddr27 = {writeAddr[13:0]};
                readAddr26 = {writeAddr[13:0]};
                readAddr25 = {writeAddr[13:0]};
                readAddr24 = {writeAddr[13:0]};
                readAddr23 = {writeAddr[13:0]};
                readAddr22  = {readAddr[12:0],  1'b0};
                readAddr21  = {readAddr[12:0],  1'b0};
                readAddr20  = {readAddr[12:0],  1'b0};
                readAddr19  = {readAddr[12:0],  1'b0};
                readAddr18  = {readAddr[12:0],  1'b0};
                readAddr17  = {readAddr[12:0],  1'b0};
                readAddr16  = {readAddr[12:0],  1'b0};
                readAddr15  = {readAddr[12:0],  1'b0};
                readAddr14  = {readAddr[12:0],  1'b0};
                readAddr13  = {readAddr[12:0],  1'b0};
                readAddr12  = {readAddr[12:0],  1'b0};
                readAddr11  = {readAddr[12:0],  1'b0};
                readAddr10  = {readAddr[12:0],  1'b0};
                readAddr9  = {readAddr[12:0],  1'b0};
                readAddr8  = {readAddr[12:0],  1'b0};
                readAddr7  = {readAddr[12:0],  1'b0};
                readAddr6  = {readAddr[10:0],  3'b0};
                readAddr5  = {readAddr[10:0],  3'b0};
                readAddr4  = {readAddr[10:0],  3'b0};
                readAddr3  = {readAddr[10:0],  3'b0};
                readAddr2  = {readAddr[9:0],  4'b0};
                readAddr1  = {readAddr[9:0],  4'b0};

                writeData54 = {17'b0, writeData[31]};
                writeData53 = {17'b0, writeData[30]};
                writeData52 = {17'b0, writeData[29]};
                writeData51 = {17'b0, writeData[28]};
                writeData50 = {17'b0, writeData[27]};
                writeData49 = {17'b0, writeData[26]};
                writeData48 = {17'b0, writeData[25]};
                writeData47 = {17'b0, writeData[24]};
                writeData46 = {17'b0, writeData[23]};
                writeData45 = {17'b0, writeData[22]};
                writeData44 = {17'b0, writeData[21]};
                writeData43 = {17'b0, writeData[20]};
                writeData42 = {17'b0, writeData[19]};
                writeData41 = {17'b0, writeData[18]};
                writeData40 = {17'b0, writeData[17]};
                writeData39 = {17'b0, writeData[16]};
                writeData38 = {17'b0, writeData[15]};
                writeData37 = {17'b0, writeData[14]};
                writeData36 = {17'b0, writeData[13]};
                writeData35 = {17'b0, writeData[12]};
                writeData34 = {17'b0, writeData[11]};
                writeData33 = {17'b0, writeData[10]};
                writeData32 = {17'b0, writeData[9]};
                writeData31 = {17'b0, writeData[8]};
                writeData30 = {17'b0, writeData[7]};
                writeData29 = {17'b0, writeData[6]};
                writeData28 = {17'b0, writeData[5]};
                writeData27 = {17'b0, writeData[4]};
                writeData26 = {17'b0, writeData[3]};
                writeData25 = {17'b0, writeData[2]};
                writeData24 = {17'b0, writeData[1]};
                writeData23 = {17'b0, writeData[0]};
                writeData22 = {16'b0, writeData[31:30]};
                writeData21 = {16'b0, writeData[29:28]};
                writeData20 = {16'b0, writeData[27:26]};
                writeData19 = {16'b0, writeData[25:24]};
                writeData18 = {16'b0, writeData[23:22]};
                writeData17 = {16'b0, writeData[21:20]};
                writeData16 = {16'b0, writeData[19:18]};
                writeData15 = {16'b0, writeData[17:16]};
                writeData14 = {16'b0, writeData[15:14]};
                writeData13 = {16'b0, writeData[13:12]};
                writeData12 = {16'b0, writeData[11:10]};
                writeData11 = {16'b0, writeData[9:8]};
                writeData10 = {16'b0, writeData[7:6]};
                writeData9 = {16'b0, writeData[5:4]};
                writeData8 = {16'b0, writeData[3:2]};
                writeData7 = {16'b0, writeData[1:0]};
                writeData6 = {10'b0, writeData[31:24]};
                writeData5 = {10'b0, writeData[23:16]};
                writeData4 = {10'b0, writeData[15:8]};
                writeData3 = {10'b0, writeData[7:0]};
                writeData2 = {1'b0, writeData[31:24], 1'b0, writeData[23:16]};
                writeData1 = {1'b0, writeData[15:8], 1'b0, writeData[7:0]};

                case (writeAddr[14:9])
                    6'b000000, 6'b000001, 6'b000010, 6'b000011,
                    6'b000100, 6'b000101, 6'b000110, 6'b000111,
                    6'b001000, 6'b001001, 6'b001010, 6'b001011,
                    6'b001100, 6'b001101, 6'b001110, 6'b001111,
                    6'b010000, 6'b010001, 6'b010010, 6'b010011,
                    6'b010100, 6'b010101, 6'b010110, 6'b010111,
                    6'b011000, 6'b011001, 6'b011010, 6'b011011,
                    6'b011100, 6'b011101, 6'b011110, 6'b011111 : begin
                        wen_a54 = {1'b0, wen};
                        wen_a53 = {1'b0, wen};
                        wen_a52 = {1'b0, wen};
                        wen_a51 = {1'b0, wen};
                        wen_a50 = {1'b0, wen};
                        wen_a49 = {1'b0, wen};
                        wen_a48 = {1'b0, wen};
                        wen_a47 = {1'b0, wen};
                        wen_a46 = {1'b0, wen};
                        wen_a45 = {1'b0, wen};
                        wen_a44 = {1'b0, wen};
                        wen_a43 = {1'b0, wen};
                        wen_a42 = {1'b0, wen};
                        wen_a41 = {1'b0, wen};
                        wen_a40 = {1'b0, wen};
                        wen_a39 = {1'b0, wen};
                        wen_a38 = {1'b0, wen};
                        wen_a37 = {1'b0, wen};
                        wen_a36 = {1'b0, wen};
                        wen_a35 = {1'b0, wen};
                        wen_a34 = {1'b0, wen};
                        wen_a33 = {1'b0, wen};
                        wen_a32 = {1'b0, wen};
                        wen_a31 = {1'b0, wen};
                        wen_a30 = {1'b0, wen};
                        wen_a29 = {1'b0, wen};
                        wen_a28 = {1'b0, wen};
                        wen_a27 = {1'b0, wen};
                        wen_a26 = {1'b0, wen};
                        wen_a25 = {1'b0, wen};
                        wen_a24 = {1'b0, wen};
                        wen_a23 = {1'b0, wen};
                        wen_a22 = {1'b0, 1'b0};
                        wen_a21 = {1'b0, 1'b0};
                        wen_a20 = {1'b0, 1'b0};
                        wen_a19 = {1'b0, 1'b0};
                        wen_a18 = {1'b0, 1'b0};
                        wen_a17 = {1'b0, 1'b0};
                        wen_a16 = {1'b0, 1'b0};
                        wen_a15 = {1'b0, 1'b0};
                        wen_a14 = {1'b0, 1'b0};
                        wen_a13 = {1'b0, 1'b0};
                        wen_a12 = {1'b0, 1'b0};
                        wen_a11 = {1'b0, 1'b0};
                        wen_a10 = {1'b0, 1'b0};
                        wen_a9 = {1'b0, 1'b0};
                        wen_a8 = {1'b0, 1'b0};
                        wen_a7 = {1'b0, 1'b0};
                        wen_a6 = {1'b0, 1'b0};
                        wen_a5 = {1'b0, 1'b0};
                        wen_a4 = {1'b0, 1'b0};
                        wen_a3 = {1'b0, 1'b0};
                        wen_a2 = {1'b0, 1'b0};
                        wen_a1 = {1'b0, 1'b0};
                    end
                    6'b100000, 6'b100001, 6'b100010, 6'b100011,
                    6'b100100, 6'b100101, 6'b100110, 6'b100111,
                    6'b101000, 6'b101001, 6'b101010, 6'b101011,
                    6'b101100, 6'b101101, 6'b101110, 6'b101111 : begin
                        wen_a54 = {1'b0, 1'b0};
                        wen_a53 = {1'b0, 1'b0};
                        wen_a52 = {1'b0, 1'b0};
                        wen_a51 = {1'b0, 1'b0};
                        wen_a50 = {1'b0, 1'b0};
                        wen_a49 = {1'b0, 1'b0};
                        wen_a48 = {1'b0, 1'b0};
                        wen_a47 = {1'b0, 1'b0};
                        wen_a46 = {1'b0, 1'b0};
                        wen_a45 = {1'b0, 1'b0};
                        wen_a44 = {1'b0, 1'b0};
                        wen_a43 = {1'b0, 1'b0};
                        wen_a42 = {1'b0, 1'b0};
                        wen_a41 = {1'b0, 1'b0};
                        wen_a40 = {1'b0, 1'b0};
                        wen_a39 = {1'b0, 1'b0};
                        wen_a38 = {1'b0, 1'b0};
                        wen_a37 = {1'b0, 1'b0};
                        wen_a36 = {1'b0, 1'b0};
                        wen_a35 = {1'b0, 1'b0};
                        wen_a34 = {1'b0, 1'b0};
                        wen_a33 = {1'b0, 1'b0};
                        wen_a32 = {1'b0, 1'b0};
                        wen_a31 = {1'b0, 1'b0};
                        wen_a30 = {1'b0, 1'b0};
                        wen_a29 = {1'b0, 1'b0};
                        wen_a28 = {1'b0, 1'b0};
                        wen_a27 = {1'b0, 1'b0};
                        wen_a26 = {1'b0, 1'b0};
                        wen_a25 = {1'b0, 1'b0};
                        wen_a24 = {1'b0, 1'b0};
                        wen_a23 = {1'b0, 1'b0};
                        wen_a22 = {1'b0, wen};
                        wen_a21 = {1'b0, wen};
                        wen_a20 = {1'b0, wen};
                        wen_a19 = {1'b0, wen};
                        wen_a18 = {1'b0, wen};
                        wen_a17 = {1'b0, wen};
                        wen_a16 = {1'b0, wen};
                        wen_a15 = {1'b0, wen};
                        wen_a14 = {1'b0, wen};
                        wen_a13 = {1'b0, wen};
                        wen_a12 = {1'b0, wen};
                        wen_a11 = {1'b0, wen};
                        wen_a10 = {1'b0, wen};
                        wen_a9 = {1'b0, wen};
                        wen_a8 = {1'b0, wen};
                        wen_a7 = {1'b0, wen};
                        wen_a6 = {1'b0, 1'b0};
                        wen_a5 = {1'b0, 1'b0};
                        wen_a4 = {1'b0, 1'b0};
                        wen_a3 = {1'b0, 1'b0};
                        wen_a2 = {1'b0, 1'b0};
                        wen_a1 = {1'b0, 1'b0};
                    end
                    6'b110000, 6'b110001, 6'b110010, 6'b110011 : begin
                        wen_a54 = {1'b0, 1'b0};
                        wen_a53 = {1'b0, 1'b0};
                        wen_a52 = {1'b0, 1'b0};
                        wen_a51 = {1'b0, 1'b0};
                        wen_a50 = {1'b0, 1'b0};
                        wen_a49 = {1'b0, 1'b0};
                        wen_a48 = {1'b0, 1'b0};
                        wen_a47 = {1'b0, 1'b0};
                        wen_a46 = {1'b0, 1'b0};
                        wen_a45 = {1'b0, 1'b0};
                        wen_a44 = {1'b0, 1'b0};
                        wen_a43 = {1'b0, 1'b0};
                        wen_a42 = {1'b0, 1'b0};
                        wen_a41 = {1'b0, 1'b0};
                        wen_a40 = {1'b0, 1'b0};
                        wen_a39 = {1'b0, 1'b0};
                        wen_a38 = {1'b0, 1'b0};
                        wen_a37 = {1'b0, 1'b0};
                        wen_a36 = {1'b0, 1'b0};
                        wen_a35 = {1'b0, 1'b0};
                        wen_a34 = {1'b0, 1'b0};
                        wen_a33 = {1'b0, 1'b0};
                        wen_a32 = {1'b0, 1'b0};
                        wen_a31 = {1'b0, 1'b0};
                        wen_a30 = {1'b0, 1'b0};
                        wen_a29 = {1'b0, 1'b0};
                        wen_a28 = {1'b0, 1'b0};
                        wen_a27 = {1'b0, 1'b0};
                        wen_a26 = {1'b0, 1'b0};
                        wen_a25 = {1'b0, 1'b0};
                        wen_a24 = {1'b0, 1'b0};
                        wen_a23 = {1'b0, 1'b0};
                        wen_a22 = {1'b0, 1'b0};
                        wen_a21 = {1'b0, 1'b0};
                        wen_a20 = {1'b0, 1'b0};
                        wen_a19 = {1'b0, 1'b0};
                        wen_a18 = {1'b0, 1'b0};
                        wen_a17 = {1'b0, 1'b0};
                        wen_a16 = {1'b0, 1'b0};
                        wen_a15 = {1'b0, 1'b0};
                        wen_a14 = {1'b0, 1'b0};
                        wen_a13 = {1'b0, 1'b0};
                        wen_a12 = {1'b0, 1'b0};
                        wen_a11 = {1'b0, 1'b0};
                        wen_a10 = {1'b0, 1'b0};
                        wen_a9 = {1'b0, 1'b0};
                        wen_a8 = {1'b0, 1'b0};
                        wen_a7 = {1'b0, 1'b0};
                        wen_a6 = {1'b0, wen};
                        wen_a5 = {1'b0, wen};
                        wen_a4 = {1'b0, wen};
                        wen_a3 = {1'b0, wen};
                        wen_a2 = {1'b0, 1'b0};
                        wen_a1 = {1'b0, 1'b0};
                    end
                    6'b110100, 6'b110101 : begin
                        wen_a54 = {1'b0, 1'b0};
                        wen_a53 = {1'b0, 1'b0};
                        wen_a52 = {1'b0, 1'b0};
                        wen_a51 = {1'b0, 1'b0};
                        wen_a50 = {1'b0, 1'b0};
                        wen_a49 = {1'b0, 1'b0};
                        wen_a48 = {1'b0, 1'b0};
                        wen_a47 = {1'b0, 1'b0};
                        wen_a46 = {1'b0, 1'b0};
                        wen_a45 = {1'b0, 1'b0};
                        wen_a44 = {1'b0, 1'b0};
                        wen_a43 = {1'b0, 1'b0};
                        wen_a42 = {1'b0, 1'b0};
                        wen_a41 = {1'b0, 1'b0};
                        wen_a40 = {1'b0, 1'b0};
                        wen_a39 = {1'b0, 1'b0};
                        wen_a38 = {1'b0, 1'b0};
                        wen_a37 = {1'b0, 1'b0};
                        wen_a36 = {1'b0, 1'b0};
                        wen_a35 = {1'b0, 1'b0};
                        wen_a34 = {1'b0, 1'b0};
                        wen_a33 = {1'b0, 1'b0};
                        wen_a32 = {1'b0, 1'b0};
                        wen_a31 = {1'b0, 1'b0};
                        wen_a30 = {1'b0, 1'b0};
                        wen_a29 = {1'b0, 1'b0};
                        wen_a28 = {1'b0, 1'b0};
                        wen_a27 = {1'b0, 1'b0};
                        wen_a26 = {1'b0, 1'b0};
                        wen_a25 = {1'b0, 1'b0};
                        wen_a24 = {1'b0, 1'b0};
                        wen_a23 = {1'b0, 1'b0};
                        wen_a22 = {1'b0, 1'b0};
                        wen_a21 = {1'b0, 1'b0};
                        wen_a20 = {1'b0, 1'b0};
                        wen_a19 = {1'b0, 1'b0};
                        wen_a18 = {1'b0, 1'b0};
                        wen_a17 = {1'b0, 1'b0};
                        wen_a16 = {1'b0, 1'b0};
                        wen_a15 = {1'b0, 1'b0};
                        wen_a14 = {1'b0, 1'b0};
                        wen_a13 = {1'b0, 1'b0};
                        wen_a12 = {1'b0, 1'b0};
                        wen_a11 = {1'b0, 1'b0};
                        wen_a10 = {1'b0, 1'b0};
                        wen_a9 = {1'b0, 1'b0};
                        wen_a8 = {1'b0, 1'b0};
                        wen_a7 = {1'b0, 1'b0};
                        wen_a6 = {1'b0, 1'b0};
                        wen_a5 = {1'b0, 1'b0};
                        wen_a4 = {1'b0, 1'b0};
                        wen_a3 = {1'b0, 1'b0};
                        wen_a2 = {wen, wen};
                        wen_a1 = {wen, wen};
                    end
                    default : begin
                        wen_a54 = {1'b0, 1'b0};
                        wen_a53 = {1'b0, 1'b0};
                        wen_a52 = {1'b0, 1'b0};
                        wen_a51 = {1'b0, 1'b0};
                        wen_a50 = {1'b0, 1'b0};
                        wen_a49 = {1'b0, 1'b0};
                        wen_a48 = {1'b0, 1'b0};
                        wen_a47 = {1'b0, 1'b0};
                        wen_a46 = {1'b0, 1'b0};
                        wen_a45 = {1'b0, 1'b0};
                        wen_a44 = {1'b0, 1'b0};
                        wen_a43 = {1'b0, 1'b0};
                        wen_a42 = {1'b0, 1'b0};
                        wen_a41 = {1'b0, 1'b0};
                        wen_a40 = {1'b0, 1'b0};
                        wen_a39 = {1'b0, 1'b0};
                        wen_a38 = {1'b0, 1'b0};
                        wen_a37 = {1'b0, 1'b0};
                        wen_a36 = {1'b0, 1'b0};
                        wen_a35 = {1'b0, 1'b0};
                        wen_a34 = {1'b0, 1'b0};
                        wen_a33 = {1'b0, 1'b0};
                        wen_a32 = {1'b0, 1'b0};
                        wen_a31 = {1'b0, 1'b0};
                        wen_a30 = {1'b0, 1'b0};
                        wen_a29 = {1'b0, 1'b0};
                        wen_a28 = {1'b0, 1'b0};
                        wen_a27 = {1'b0, 1'b0};
                        wen_a26 = {1'b0, 1'b0};
                        wen_a25 = {1'b0, 1'b0};
                        wen_a24 = {1'b0, 1'b0};
                        wen_a23 = {1'b0, 1'b0};
                        wen_a22 = {1'b0, 1'b0};
                        wen_a21 = {1'b0, 1'b0};
                        wen_a20 = {1'b0, 1'b0};
                        wen_a19 = {1'b0, 1'b0};
                        wen_a18 = {1'b0, 1'b0};
                        wen_a17 = {1'b0, 1'b0};
                        wen_a16 = {1'b0, 1'b0};
                        wen_a15 = {1'b0, 1'b0};
                        wen_a14 = {1'b0, 1'b0};
                        wen_a13 = {1'b0, 1'b0};
                        wen_a12 = {1'b0, 1'b0};
                        wen_a11 = {1'b0, 1'b0};
                        wen_a10 = {1'b0, 1'b0};
                        wen_a9 = {1'b0, 1'b0};
                        wen_a8 = {1'b0, 1'b0};
                        wen_a7 = {1'b0, 1'b0};
                        wen_a6 = {1'b0, 1'b0};
                        wen_a5 = {1'b0, 1'b0};
                        wen_a4 = {1'b0, 1'b0};
                        wen_a3 = {1'b0, 1'b0};
                        wen_a2 = {1'b0, 1'b0};
                        wen_a1 = {1'b0, 1'b0};
                    end
                endcase

                case (ckRdAddr[14:9])
                    6'b000000, 6'b000001, 6'b000010, 6'b000011,
                    6'b000100, 6'b000101, 6'b000110, 6'b000111,
                    6'b001000, 6'b001001, 6'b001010, 6'b001011,
                    6'b001100, 6'b001101, 6'b001110, 6'b001111,
                    6'b010000, 6'b010001, 6'b010010, 6'b010011,
                    6'b010100, 6'b010101, 6'b010110, 6'b010111,
                    6'b011000, 6'b011001, 6'b011010, 6'b011011,
                    6'b011100, 6'b011101, 6'b011110, 6'b011111 : begin
                        readData = {
                                        readData54[0],
                                        readData53[0],
                                        readData52[0],
                                        readData51[0],
                                        readData50[0],
                                        readData49[0],
                                        readData48[0],
                                        readData47[0],
                                        readData46[0],
                                        readData45[0],
                                        readData44[0],
                                        readData43[0],
                                        readData42[0],
                                        readData41[0],
                                        readData40[0],
                                        readData39[0],
                                        readData38[0],
                                        readData37[0],
                                        readData36[0],
                                        readData35[0],
                                        readData34[0],
                                        readData33[0],
                                        readData32[0],
                                        readData31[0],
                                        readData30[0],
                                        readData29[0],
                                        readData28[0],
                                        readData27[0],
                                        readData26[0],
                                        readData25[0],
                                        readData24[0],
                                        readData23[0]
                        };
                    end
                    6'b100000, 6'b100001, 6'b100010, 6'b100011,
                    6'b100100, 6'b100101, 6'b100110, 6'b100111,
                    6'b101000, 6'b101001, 6'b101010, 6'b101011,
                    6'b101100, 6'b101101, 6'b101110, 6'b101111 : begin
                        readData = {
                                        readData22[1:0],
                                        readData21[1:0],
                                        readData20[1:0],
                                        readData19[1:0],
                                        readData18[1:0],
                                        readData17[1:0],
                                        readData16[1:0],
                                        readData15[1:0],
                                        readData14[1:0],
                                        readData13[1:0],
                                        readData12[1:0],
                                        readData11[1:0],
                                        readData10[1:0],
                                        readData9[1:0],
                                        readData8[1:0],
                                        readData7[1:0]
                        };
                    end
                    6'b110000, 6'b110001, 6'b110010, 6'b110011 : begin
                        readData = {readData6[7:0],readData5[7:0],readData4[7:0],readData3[7:0]};
                    end
                    6'b110100, 6'b110101 : begin
                        readData = {readData2[16:9],readData2[7:0],readData1[16:9],readData1[7:0]};
                    end
                    default : begin
                        readData = 32'b0;
                    end
                endcase
            end        
            28160: begin
                width54 = 3'b000;
                width53 = 3'b000;
                width52 = 3'b000;
                width51 = 3'b000;
                width50 = 3'b000;
                width49 = 3'b000;
                width48 = 3'b000;
                width47 = 3'b000;
                width46 = 3'b000;
                width45 = 3'b000;
                width44 = 3'b000;
                width43 = 3'b000;
                width42 = 3'b000;
                width41 = 3'b000;
                width40 = 3'b000;
                width39 = 3'b000;
                width38 = 3'b000;
                width37 = 3'b000;
                width36 = 3'b000;
                width35 = 3'b000;
                width34 = 3'b000;
                width33 = 3'b000;
                width32 = 3'b000;
                width31 = 3'b000;
                width30 = 3'b000;
                width29 = 3'b000;
                width28 = 3'b000;
                width27 = 3'b000;
                width26 = 3'b000;
                width25 = 3'b000;
                width24 = 3'b000;
                width23 = 3'b000;
                width22 = 3'b001;
                width21 = 3'b001;
                width20 = 3'b001;
                width19 = 3'b001;
                width18 = 3'b001;
                width17 = 3'b001;
                width16 = 3'b001;
                width15 = 3'b001;
                width14 = 3'b001;
                width13 = 3'b001;
                width12 = 3'b001;
                width11 = 3'b001;
                width10 = 3'b001;
                width9 = 3'b001;
                width8 = 3'b001;
                width7 = 3'b001;
                width6 = 3'b011;
                width5 = 3'b011;
                width4 = 3'b011;
                width3 = 3'b011;
                width2 = 3'b100;
                width1 = 3'b100;
                width0 = 3'b101;

                writeAddr54 = {writeAddr[13:0]};
                writeAddr53 = {writeAddr[13:0]};
                writeAddr52 = {writeAddr[13:0]};
                writeAddr51 = {writeAddr[13:0]};
                writeAddr50 = {writeAddr[13:0]};
                writeAddr49 = {writeAddr[13:0]};
                writeAddr48 = {writeAddr[13:0]};
                writeAddr47 = {writeAddr[13:0]};
                writeAddr46 = {writeAddr[13:0]};
                writeAddr45 = {writeAddr[13:0]};
                writeAddr44 = {writeAddr[13:0]};
                writeAddr43 = {writeAddr[13:0]};
                writeAddr42 = {writeAddr[13:0]};
                writeAddr41 = {writeAddr[13:0]};
                writeAddr40 = {writeAddr[13:0]};
                writeAddr39 = {writeAddr[13:0]};
                writeAddr38 = {writeAddr[13:0]};
                writeAddr37 = {writeAddr[13:0]};
                writeAddr36 = {writeAddr[13:0]};
                writeAddr35 = {writeAddr[13:0]};
                writeAddr34 = {writeAddr[13:0]};
                writeAddr33 = {writeAddr[13:0]};
                writeAddr32 = {writeAddr[13:0]};
                writeAddr31 = {writeAddr[13:0]};
                writeAddr30 = {writeAddr[13:0]};
                writeAddr29 = {writeAddr[13:0]};
                writeAddr28 = {writeAddr[13:0]};
                writeAddr27 = {writeAddr[13:0]};
                writeAddr26 = {writeAddr[13:0]};
                writeAddr25 = {writeAddr[13:0]};
                writeAddr24 = {writeAddr[13:0]};
                writeAddr23 = {writeAddr[13:0]};
                writeAddr22 = {writeAddr[12:0], 1'b0};
                writeAddr21 = {writeAddr[12:0], 1'b0};
                writeAddr20 = {writeAddr[12:0], 1'b0};
                writeAddr19 = {writeAddr[12:0], 1'b0};
                writeAddr18 = {writeAddr[12:0], 1'b0};
                writeAddr17 = {writeAddr[12:0], 1'b0};
                writeAddr16 = {writeAddr[12:0], 1'b0};
                writeAddr15 = {writeAddr[12:0], 1'b0};
                writeAddr14 = {writeAddr[12:0], 1'b0};
                writeAddr13 = {writeAddr[12:0], 1'b0};
                writeAddr12 = {writeAddr[12:0], 1'b0};
                writeAddr11 = {writeAddr[12:0], 1'b0};
                writeAddr10 = {writeAddr[12:0], 1'b0};
                writeAddr9 = {writeAddr[12:0], 1'b0};
                writeAddr8 = {writeAddr[12:0], 1'b0};
                writeAddr7 = {writeAddr[12:0], 1'b0};
                writeAddr6 = {writeAddr[10:0], 3'b0};
                writeAddr5 = {writeAddr[10:0], 3'b0};
                writeAddr4 = {writeAddr[10:0], 3'b0};
                writeAddr3 = {writeAddr[10:0], 3'b0};
                writeAddr2 = {writeAddr[9:0], 4'b0};
                writeAddr1 = {writeAddr[9:0], 4'b0};
                writeAddr0 = {writeAddr[8:0], 5'b0};

                readAddr54 = {writeAddr[13:0]};
                readAddr53 = {writeAddr[13:0]};
                readAddr52 = {writeAddr[13:0]};
                readAddr51 = {writeAddr[13:0]};
                readAddr50 = {writeAddr[13:0]};
                readAddr49 = {writeAddr[13:0]};
                readAddr48 = {writeAddr[13:0]};
                readAddr47 = {writeAddr[13:0]};
                readAddr46 = {writeAddr[13:0]};
                readAddr45 = {writeAddr[13:0]};
                readAddr44 = {writeAddr[13:0]};
                readAddr43 = {writeAddr[13:0]};
                readAddr42 = {writeAddr[13:0]};
                readAddr41 = {writeAddr[13:0]};
                readAddr40 = {writeAddr[13:0]};
                readAddr39 = {writeAddr[13:0]};
                readAddr38 = {writeAddr[13:0]};
                readAddr37 = {writeAddr[13:0]};
                readAddr36 = {writeAddr[13:0]};
                readAddr35 = {writeAddr[13:0]};
                readAddr34 = {writeAddr[13:0]};
                readAddr33 = {writeAddr[13:0]};
                readAddr32 = {writeAddr[13:0]};
                readAddr31 = {writeAddr[13:0]};
                readAddr30 = {writeAddr[13:0]};
                readAddr29 = {writeAddr[13:0]};
                readAddr28 = {writeAddr[13:0]};
                readAddr27 = {writeAddr[13:0]};
                readAddr26 = {writeAddr[13:0]};
                readAddr25 = {writeAddr[13:0]};
                readAddr24 = {writeAddr[13:0]};
                readAddr23 = {writeAddr[13:0]};
                readAddr22  = {readAddr[12:0],  1'b0};
                readAddr21  = {readAddr[12:0],  1'b0};
                readAddr20  = {readAddr[12:0],  1'b0};
                readAddr19  = {readAddr[12:0],  1'b0};
                readAddr18  = {readAddr[12:0],  1'b0};
                readAddr17  = {readAddr[12:0],  1'b0};
                readAddr16  = {readAddr[12:0],  1'b0};
                readAddr15  = {readAddr[12:0],  1'b0};
                readAddr14  = {readAddr[12:0],  1'b0};
                readAddr13  = {readAddr[12:0],  1'b0};
                readAddr12  = {readAddr[12:0],  1'b0};
                readAddr11  = {readAddr[12:0],  1'b0};
                readAddr10  = {readAddr[12:0],  1'b0};
                readAddr9  = {readAddr[12:0],  1'b0};
                readAddr8  = {readAddr[12:0],  1'b0};
                readAddr7  = {readAddr[12:0],  1'b0};
                readAddr6  = {readAddr[10:0],  3'b0};
                readAddr5  = {readAddr[10:0],  3'b0};
                readAddr4  = {readAddr[10:0],  3'b0};
                readAddr3  = {readAddr[10:0],  3'b0};
                readAddr2  = {readAddr[9:0],  4'b0};
                readAddr1  = {readAddr[9:0],  4'b0};
                readAddr0  = {readAddr[8:0],  5'b0};

                writeData54 = {17'b0, writeData[31]};
                writeData53 = {17'b0, writeData[30]};
                writeData52 = {17'b0, writeData[29]};
                writeData51 = {17'b0, writeData[28]};
                writeData50 = {17'b0, writeData[27]};
                writeData49 = {17'b0, writeData[26]};
                writeData48 = {17'b0, writeData[25]};
                writeData47 = {17'b0, writeData[24]};
                writeData46 = {17'b0, writeData[23]};
                writeData45 = {17'b0, writeData[22]};
                writeData44 = {17'b0, writeData[21]};
                writeData43 = {17'b0, writeData[20]};
                writeData42 = {17'b0, writeData[19]};
                writeData41 = {17'b0, writeData[18]};
                writeData40 = {17'b0, writeData[17]};
                writeData39 = {17'b0, writeData[16]};
                writeData38 = {17'b0, writeData[15]};
                writeData37 = {17'b0, writeData[14]};
                writeData36 = {17'b0, writeData[13]};
                writeData35 = {17'b0, writeData[12]};
                writeData34 = {17'b0, writeData[11]};
                writeData33 = {17'b0, writeData[10]};
                writeData32 = {17'b0, writeData[9]};
                writeData31 = {17'b0, writeData[8]};
                writeData30 = {17'b0, writeData[7]};
                writeData29 = {17'b0, writeData[6]};
                writeData28 = {17'b0, writeData[5]};
                writeData27 = {17'b0, writeData[4]};
                writeData26 = {17'b0, writeData[3]};
                writeData25 = {17'b0, writeData[2]};
                writeData24 = {17'b0, writeData[1]};
                writeData23 = {17'b0, writeData[0]};
                writeData22 = {16'b0, writeData[31:30]};
                writeData21 = {16'b0, writeData[29:28]};
                writeData20 = {16'b0, writeData[27:26]};
                writeData19 = {16'b0, writeData[25:24]};
                writeData18 = {16'b0, writeData[23:22]};
                writeData17 = {16'b0, writeData[21:20]};
                writeData16 = {16'b0, writeData[19:18]};
                writeData15 = {16'b0, writeData[17:16]};
                writeData14 = {16'b0, writeData[15:14]};
                writeData13 = {16'b0, writeData[13:12]};
                writeData12 = {16'b0, writeData[11:10]};
                writeData11 = {16'b0, writeData[9:8]};
                writeData10 = {16'b0, writeData[7:6]};
                writeData9 = {16'b0, writeData[5:4]};
                writeData8 = {16'b0, writeData[3:2]};
                writeData7 = {16'b0, writeData[1:0]};
                writeData6 = {10'b0, writeData[31:24]};
                writeData5 = {10'b0, writeData[23:16]};
                writeData4 = {10'b0, writeData[15:8]};
                writeData3 = {10'b0, writeData[7:0]};
                writeData2 = {1'b0, writeData[31:24], 1'b0, writeData[23:16]};
                writeData1 = {1'b0, writeData[15:8], 1'b0, writeData[7:0]};
                writeData0 = {1'b0, writeData[31:24], 1'b0, writeData[23:16], 1'b0, writeData[15:8], 1'b0, writeData[7:0]};

                case (writeAddr[14:9])
                    6'b000000, 6'b000001, 6'b000010, 6'b000011,
                    6'b000100, 6'b000101, 6'b000110, 6'b000111,
                    6'b001000, 6'b001001, 6'b001010, 6'b001011,
                    6'b001100, 6'b001101, 6'b001110, 6'b001111,
                    6'b010000, 6'b010001, 6'b010010, 6'b010011,
                    6'b010100, 6'b010101, 6'b010110, 6'b010111,
                    6'b011000, 6'b011001, 6'b011010, 6'b011011,
                    6'b011100, 6'b011101, 6'b011110, 6'b011111 : begin
                        wen_a54 = {1'b0, wen};
                        wen_a53 = {1'b0, wen};
                        wen_a52 = {1'b0, wen};
                        wen_a51 = {1'b0, wen};
                        wen_a50 = {1'b0, wen};
                        wen_a49 = {1'b0, wen};
                        wen_a48 = {1'b0, wen};
                        wen_a47 = {1'b0, wen};
                        wen_a46 = {1'b0, wen};
                        wen_a45 = {1'b0, wen};
                        wen_a44 = {1'b0, wen};
                        wen_a43 = {1'b0, wen};
                        wen_a42 = {1'b0, wen};
                        wen_a41 = {1'b0, wen};
                        wen_a40 = {1'b0, wen};
                        wen_a39 = {1'b0, wen};
                        wen_a38 = {1'b0, wen};
                        wen_a37 = {1'b0, wen};
                        wen_a36 = {1'b0, wen};
                        wen_a35 = {1'b0, wen};
                        wen_a34 = {1'b0, wen};
                        wen_a33 = {1'b0, wen};
                        wen_a32 = {1'b0, wen};
                        wen_a31 = {1'b0, wen};
                        wen_a30 = {1'b0, wen};
                        wen_a29 = {1'b0, wen};
                        wen_a28 = {1'b0, wen};
                        wen_a27 = {1'b0, wen};
                        wen_a26 = {1'b0, wen};
                        wen_a25 = {1'b0, wen};
                        wen_a24 = {1'b0, wen};
                        wen_a23 = {1'b0, wen};
                        wen_a22 = {1'b0, 1'b0};
                        wen_a21 = {1'b0, 1'b0};
                        wen_a20 = {1'b0, 1'b0};
                        wen_a19 = {1'b0, 1'b0};
                        wen_a18 = {1'b0, 1'b0};
                        wen_a17 = {1'b0, 1'b0};
                        wen_a16 = {1'b0, 1'b0};
                        wen_a15 = {1'b0, 1'b0};
                        wen_a14 = {1'b0, 1'b0};
                        wen_a13 = {1'b0, 1'b0};
                        wen_a12 = {1'b0, 1'b0};
                        wen_a11 = {1'b0, 1'b0};
                        wen_a10 = {1'b0, 1'b0};
                        wen_a9 = {1'b0, 1'b0};
                        wen_a8 = {1'b0, 1'b0};
                        wen_a7 = {1'b0, 1'b0};
                        wen_a6 = {1'b0, 1'b0};
                        wen_a5 = {1'b0, 1'b0};
                        wen_a4 = {1'b0, 1'b0};
                        wen_a3 = {1'b0, 1'b0};
                        wen_a2 = {1'b0, 1'b0};
                        wen_a1 = {1'b0, 1'b0};
                        wen_a0 = {1'b0, 1'b0};
                        wen_b0 = {1'b0, 1'b0};
                    end
                    6'b100000, 6'b100001, 6'b100010, 6'b100011,
                    6'b100100, 6'b100101, 6'b100110, 6'b100111,
                    6'b101000, 6'b101001, 6'b101010, 6'b101011,
                    6'b101100, 6'b101101, 6'b101110, 6'b101111 : begin
                        wen_a54 = {1'b0, 1'b0};
                        wen_a53 = {1'b0, 1'b0};
                        wen_a52 = {1'b0, 1'b0};
                        wen_a51 = {1'b0, 1'b0};
                        wen_a50 = {1'b0, 1'b0};
                        wen_a49 = {1'b0, 1'b0};
                        wen_a48 = {1'b0, 1'b0};
                        wen_a47 = {1'b0, 1'b0};
                        wen_a46 = {1'b0, 1'b0};
                        wen_a45 = {1'b0, 1'b0};
                        wen_a44 = {1'b0, 1'b0};
                        wen_a43 = {1'b0, 1'b0};
                        wen_a42 = {1'b0, 1'b0};
                        wen_a41 = {1'b0, 1'b0};
                        wen_a40 = {1'b0, 1'b0};
                        wen_a39 = {1'b0, 1'b0};
                        wen_a38 = {1'b0, 1'b0};
                        wen_a37 = {1'b0, 1'b0};
                        wen_a36 = {1'b0, 1'b0};
                        wen_a35 = {1'b0, 1'b0};
                        wen_a34 = {1'b0, 1'b0};
                        wen_a33 = {1'b0, 1'b0};
                        wen_a32 = {1'b0, 1'b0};
                        wen_a31 = {1'b0, 1'b0};
                        wen_a30 = {1'b0, 1'b0};
                        wen_a29 = {1'b0, 1'b0};
                        wen_a28 = {1'b0, 1'b0};
                        wen_a27 = {1'b0, 1'b0};
                        wen_a26 = {1'b0, 1'b0};
                        wen_a25 = {1'b0, 1'b0};
                        wen_a24 = {1'b0, 1'b0};
                        wen_a23 = {1'b0, 1'b0};
                        wen_a22 = {1'b0, wen};
                        wen_a21 = {1'b0, wen};
                        wen_a20 = {1'b0, wen};
                        wen_a19 = {1'b0, wen};
                        wen_a18 = {1'b0, wen};
                        wen_a17 = {1'b0, wen};
                        wen_a16 = {1'b0, wen};
                        wen_a15 = {1'b0, wen};
                        wen_a14 = {1'b0, wen};
                        wen_a13 = {1'b0, wen};
                        wen_a12 = {1'b0, wen};
                        wen_a11 = {1'b0, wen};
                        wen_a10 = {1'b0, wen};
                        wen_a9 = {1'b0, wen};
                        wen_a8 = {1'b0, wen};
                        wen_a7 = {1'b0, wen};
                        wen_a6 = {1'b0, 1'b0};
                        wen_a5 = {1'b0, 1'b0};
                        wen_a4 = {1'b0, 1'b0};
                        wen_a3 = {1'b0, 1'b0};
                        wen_a2 = {1'b0, 1'b0};
                        wen_a1 = {1'b0, 1'b0};
                        wen_a0 = {1'b0, 1'b0};
                        wen_b0 = {1'b0, 1'b0};
                    end
                    6'b110000, 6'b110001, 6'b110010, 6'b110011 : begin
                        wen_a54 = {1'b0, 1'b0};
                        wen_a53 = {1'b0, 1'b0};
                        wen_a52 = {1'b0, 1'b0};
                        wen_a51 = {1'b0, 1'b0};
                        wen_a50 = {1'b0, 1'b0};
                        wen_a49 = {1'b0, 1'b0};
                        wen_a48 = {1'b0, 1'b0};
                        wen_a47 = {1'b0, 1'b0};
                        wen_a46 = {1'b0, 1'b0};
                        wen_a45 = {1'b0, 1'b0};
                        wen_a44 = {1'b0, 1'b0};
                        wen_a43 = {1'b0, 1'b0};
                        wen_a42 = {1'b0, 1'b0};
                        wen_a41 = {1'b0, 1'b0};
                        wen_a40 = {1'b0, 1'b0};
                        wen_a39 = {1'b0, 1'b0};
                        wen_a38 = {1'b0, 1'b0};
                        wen_a37 = {1'b0, 1'b0};
                        wen_a36 = {1'b0, 1'b0};
                        wen_a35 = {1'b0, 1'b0};
                        wen_a34 = {1'b0, 1'b0};
                        wen_a33 = {1'b0, 1'b0};
                        wen_a32 = {1'b0, 1'b0};
                        wen_a31 = {1'b0, 1'b0};
                        wen_a30 = {1'b0, 1'b0};
                        wen_a29 = {1'b0, 1'b0};
                        wen_a28 = {1'b0, 1'b0};
                        wen_a27 = {1'b0, 1'b0};
                        wen_a26 = {1'b0, 1'b0};
                        wen_a25 = {1'b0, 1'b0};
                        wen_a24 = {1'b0, 1'b0};
                        wen_a23 = {1'b0, 1'b0};
                        wen_a22 = {1'b0, 1'b0};
                        wen_a21 = {1'b0, 1'b0};
                        wen_a20 = {1'b0, 1'b0};
                        wen_a19 = {1'b0, 1'b0};
                        wen_a18 = {1'b0, 1'b0};
                        wen_a17 = {1'b0, 1'b0};
                        wen_a16 = {1'b0, 1'b0};
                        wen_a15 = {1'b0, 1'b0};
                        wen_a14 = {1'b0, 1'b0};
                        wen_a13 = {1'b0, 1'b0};
                        wen_a12 = {1'b0, 1'b0};
                        wen_a11 = {1'b0, 1'b0};
                        wen_a10 = {1'b0, 1'b0};
                        wen_a9 = {1'b0, 1'b0};
                        wen_a8 = {1'b0, 1'b0};
                        wen_a7 = {1'b0, 1'b0};
                        wen_a6 = {1'b0, wen};
                        wen_a5 = {1'b0, wen};
                        wen_a4 = {1'b0, wen};
                        wen_a3 = {1'b0, wen};
                        wen_a2 = {1'b0, 1'b0};
                        wen_a1 = {1'b0, 1'b0};
                        wen_a0 = {1'b0, 1'b0};
                        wen_b0 = {1'b0, 1'b0};
                    end
                    6'b110100, 6'b110101 : begin
                        wen_a54 = {1'b0, 1'b0};
                        wen_a53 = {1'b0, 1'b0};
                        wen_a52 = {1'b0, 1'b0};
                        wen_a51 = {1'b0, 1'b0};
                        wen_a50 = {1'b0, 1'b0};
                        wen_a49 = {1'b0, 1'b0};
                        wen_a48 = {1'b0, 1'b0};
                        wen_a47 = {1'b0, 1'b0};
                        wen_a46 = {1'b0, 1'b0};
                        wen_a45 = {1'b0, 1'b0};
                        wen_a44 = {1'b0, 1'b0};
                        wen_a43 = {1'b0, 1'b0};
                        wen_a42 = {1'b0, 1'b0};
                        wen_a41 = {1'b0, 1'b0};
                        wen_a40 = {1'b0, 1'b0};
                        wen_a39 = {1'b0, 1'b0};
                        wen_a38 = {1'b0, 1'b0};
                        wen_a37 = {1'b0, 1'b0};
                        wen_a36 = {1'b0, 1'b0};
                        wen_a35 = {1'b0, 1'b0};
                        wen_a34 = {1'b0, 1'b0};
                        wen_a33 = {1'b0, 1'b0};
                        wen_a32 = {1'b0, 1'b0};
                        wen_a31 = {1'b0, 1'b0};
                        wen_a30 = {1'b0, 1'b0};
                        wen_a29 = {1'b0, 1'b0};
                        wen_a28 = {1'b0, 1'b0};
                        wen_a27 = {1'b0, 1'b0};
                        wen_a26 = {1'b0, 1'b0};
                        wen_a25 = {1'b0, 1'b0};
                        wen_a24 = {1'b0, 1'b0};
                        wen_a23 = {1'b0, 1'b0};
                        wen_a22 = {1'b0, 1'b0};
                        wen_a21 = {1'b0, 1'b0};
                        wen_a20 = {1'b0, 1'b0};
                        wen_a19 = {1'b0, 1'b0};
                        wen_a18 = {1'b0, 1'b0};
                        wen_a17 = {1'b0, 1'b0};
                        wen_a16 = {1'b0, 1'b0};
                        wen_a15 = {1'b0, 1'b0};
                        wen_a14 = {1'b0, 1'b0};
                        wen_a13 = {1'b0, 1'b0};
                        wen_a12 = {1'b0, 1'b0};
                        wen_a11 = {1'b0, 1'b0};
                        wen_a10 = {1'b0, 1'b0};
                        wen_a9 = {1'b0, 1'b0};
                        wen_a8 = {1'b0, 1'b0};
                        wen_a7 = {1'b0, 1'b0};
                        wen_a6 = {1'b0, 1'b0};
                        wen_a5 = {1'b0, 1'b0};
                        wen_a4 = {1'b0, 1'b0};
                        wen_a3 = {1'b0, 1'b0};
                        wen_a2 = {wen, wen};
                        wen_a1 = {wen, wen};
                        wen_a0 = {1'b0, 1'b0};
                        wen_b0 = {1'b0, 1'b0};
                    end
                    6'b110110 : begin
                        wen_a54 = {1'b0, 1'b0};
                        wen_a53 = {1'b0, 1'b0};
                        wen_a52 = {1'b0, 1'b0};
                        wen_a51 = {1'b0, 1'b0};
                        wen_a50 = {1'b0, 1'b0};
                        wen_a49 = {1'b0, 1'b0};
                        wen_a48 = {1'b0, 1'b0};
                        wen_a47 = {1'b0, 1'b0};
                        wen_a46 = {1'b0, 1'b0};
                        wen_a45 = {1'b0, 1'b0};
                        wen_a44 = {1'b0, 1'b0};
                        wen_a43 = {1'b0, 1'b0};
                        wen_a42 = {1'b0, 1'b0};
                        wen_a41 = {1'b0, 1'b0};
                        wen_a40 = {1'b0, 1'b0};
                        wen_a39 = {1'b0, 1'b0};
                        wen_a38 = {1'b0, 1'b0};
                        wen_a37 = {1'b0, 1'b0};
                        wen_a36 = {1'b0, 1'b0};
                        wen_a35 = {1'b0, 1'b0};
                        wen_a34 = {1'b0, 1'b0};
                        wen_a33 = {1'b0, 1'b0};
                        wen_a32 = {1'b0, 1'b0};
                        wen_a31 = {1'b0, 1'b0};
                        wen_a30 = {1'b0, 1'b0};
                        wen_a29 = {1'b0, 1'b0};
                        wen_a28 = {1'b0, 1'b0};
                        wen_a27 = {1'b0, 1'b0};
                        wen_a26 = {1'b0, 1'b0};
                        wen_a25 = {1'b0, 1'b0};
                        wen_a24 = {1'b0, 1'b0};
                        wen_a23 = {1'b0, 1'b0};
                        wen_a22 = {1'b0, 1'b0};
                        wen_a21 = {1'b0, 1'b0};
                        wen_a20 = {1'b0, 1'b0};
                        wen_a19 = {1'b0, 1'b0};
                        wen_a18 = {1'b0, 1'b0};
                        wen_a17 = {1'b0, 1'b0};
                        wen_a16 = {1'b0, 1'b0};
                        wen_a15 = {1'b0, 1'b0};
                        wen_a14 = {1'b0, 1'b0};
                        wen_a13 = {1'b0, 1'b0};
                        wen_a12 = {1'b0, 1'b0};
                        wen_a11 = {1'b0, 1'b0};
                        wen_a10 = {1'b0, 1'b0};
                        wen_a9 = {1'b0, 1'b0};
                        wen_a8 = {1'b0, 1'b0};
                        wen_a7 = {1'b0, 1'b0};
                        wen_a6 = {1'b0, 1'b0};
                        wen_a5 = {1'b0, 1'b0};
                        wen_a4 = {1'b0, 1'b0};
                        wen_a3 = {1'b0, 1'b0};
                        wen_a2 = {1'b0, 1'b0};
                        wen_a1 = {1'b0, 1'b0};
                        wen_a0 = {wen, wen};
                        wen_b0 = {wen, wen};
                    end
                    default : begin
                        wen_a54 = {1'b0, 1'b0};
                        wen_a53 = {1'b0, 1'b0};
                        wen_a52 = {1'b0, 1'b0};
                        wen_a51 = {1'b0, 1'b0};
                        wen_a50 = {1'b0, 1'b0};
                        wen_a49 = {1'b0, 1'b0};
                        wen_a48 = {1'b0, 1'b0};
                        wen_a47 = {1'b0, 1'b0};
                        wen_a46 = {1'b0, 1'b0};
                        wen_a45 = {1'b0, 1'b0};
                        wen_a44 = {1'b0, 1'b0};
                        wen_a43 = {1'b0, 1'b0};
                        wen_a42 = {1'b0, 1'b0};
                        wen_a41 = {1'b0, 1'b0};
                        wen_a40 = {1'b0, 1'b0};
                        wen_a39 = {1'b0, 1'b0};
                        wen_a38 = {1'b0, 1'b0};
                        wen_a37 = {1'b0, 1'b0};
                        wen_a36 = {1'b0, 1'b0};
                        wen_a35 = {1'b0, 1'b0};
                        wen_a34 = {1'b0, 1'b0};
                        wen_a33 = {1'b0, 1'b0};
                        wen_a32 = {1'b0, 1'b0};
                        wen_a31 = {1'b0, 1'b0};
                        wen_a30 = {1'b0, 1'b0};
                        wen_a29 = {1'b0, 1'b0};
                        wen_a28 = {1'b0, 1'b0};
                        wen_a27 = {1'b0, 1'b0};
                        wen_a26 = {1'b0, 1'b0};
                        wen_a25 = {1'b0, 1'b0};
                        wen_a24 = {1'b0, 1'b0};
                        wen_a23 = {1'b0, 1'b0};
                        wen_a22 = {1'b0, 1'b0};
                        wen_a21 = {1'b0, 1'b0};
                        wen_a20 = {1'b0, 1'b0};
                        wen_a19 = {1'b0, 1'b0};
                        wen_a18 = {1'b0, 1'b0};
                        wen_a17 = {1'b0, 1'b0};
                        wen_a16 = {1'b0, 1'b0};
                        wen_a15 = {1'b0, 1'b0};
                        wen_a14 = {1'b0, 1'b0};
                        wen_a13 = {1'b0, 1'b0};
                        wen_a12 = {1'b0, 1'b0};
                        wen_a11 = {1'b0, 1'b0};
                        wen_a10 = {1'b0, 1'b0};
                        wen_a9 = {1'b0, 1'b0};
                        wen_a8 = {1'b0, 1'b0};
                        wen_a7 = {1'b0, 1'b0};
                        wen_a6 = {1'b0, 1'b0};
                        wen_a5 = {1'b0, 1'b0};
                        wen_a4 = {1'b0, 1'b0};
                        wen_a3 = {1'b0, 1'b0};
                        wen_a2 = {1'b0, 1'b0};
                        wen_a1 = {1'b0, 1'b0};
                        wen_a0 = {1'b0, 1'b0};
                        wen_b0 = {1'b0, 1'b0};
                    end
                endcase

                case (ckRdAddr[14:9])
                    6'b000000, 6'b000001, 6'b000010, 6'b000011,
                    6'b000100, 6'b000101, 6'b000110, 6'b000111,
                    6'b001000, 6'b001001, 6'b001010, 6'b001011,
                    6'b001100, 6'b001101, 6'b001110, 6'b001111,
                    6'b010000, 6'b010001, 6'b010010, 6'b010011,
                    6'b010100, 6'b010101, 6'b010110, 6'b010111,
                    6'b011000, 6'b011001, 6'b011010, 6'b011011,
                    6'b011100, 6'b011101, 6'b011110, 6'b011111 : begin
                        readData = {
                                        readData54[0],
                                        readData53[0],
                                        readData52[0],
                                        readData51[0],
                                        readData50[0],
                                        readData49[0],
                                        readData48[0],
                                        readData47[0],
                                        readData46[0],
                                        readData45[0],
                                        readData44[0],
                                        readData43[0],
                                        readData42[0],
                                        readData41[0],
                                        readData40[0],
                                        readData39[0],
                                        readData38[0],
                                        readData37[0],
                                        readData36[0],
                                        readData35[0],
                                        readData34[0],
                                        readData33[0],
                                        readData32[0],
                                        readData31[0],
                                        readData30[0],
                                        readData29[0],
                                        readData28[0],
                                        readData27[0],
                                        readData26[0],
                                        readData25[0],
                                        readData24[0],
                                        readData23[0]
                        };
                    end
                    6'b100000, 6'b100001, 6'b100010, 6'b100011,
                    6'b100100, 6'b100101, 6'b100110, 6'b100111,
                    6'b101000, 6'b101001, 6'b101010, 6'b101011,
                    6'b101100, 6'b101101, 6'b101110, 6'b101111 : begin
                        readData = {
                                        readData22[1:0],
                                        readData21[1:0],
                                        readData20[1:0],
                                        readData19[1:0],
                                        readData18[1:0],
                                        readData17[1:0],
                                        readData16[1:0],
                                        readData15[1:0],
                                        readData14[1:0],
                                        readData13[1:0],
                                        readData12[1:0],
                                        readData11[1:0],
                                        readData10[1:0],
                                        readData9[1:0],
                                        readData8[1:0],
                                        readData7[1:0]
                        };
                    end
                    6'b110000, 6'b110001, 6'b110010, 6'b110011 : begin
                        readData = {readData6[7:0],readData5[7:0],readData4[7:0],readData3[7:0]};
                    end
                    6'b110100, 6'b110101 : begin
                        readData = {readData2[16:9],readData2[7:0],readData1[16:9],readData1[7:0]};
                    end
                    6'b110110 : begin
                        readData = {readData0[34:27],readData0[25:18],readData0[16:9],readData0[7:0]};
                    end
                    default : begin
                        readData = 32'b0;
                    end
                endcase
            end        
            28672: begin
                width56 = 3'b000;
                width55 = 3'b000;
                width54 = 3'b000;
                width53 = 3'b000;
                width52 = 3'b000;
                width51 = 3'b000;
                width50 = 3'b000;
                width49 = 3'b000;
                width48 = 3'b000;
                width47 = 3'b000;
                width46 = 3'b000;
                width45 = 3'b000;
                width44 = 3'b000;
                width43 = 3'b000;
                width42 = 3'b000;
                width41 = 3'b000;
                width40 = 3'b000;
                width39 = 3'b000;
                width38 = 3'b000;
                width37 = 3'b000;
                width36 = 3'b000;
                width35 = 3'b000;
                width34 = 3'b000;
                width33 = 3'b000;
                width32 = 3'b000;
                width31 = 3'b000;
                width30 = 3'b000;
                width29 = 3'b000;
                width28 = 3'b000;
                width27 = 3'b000;
                width26 = 3'b000;
                width25 = 3'b000;
                width24 = 3'b001;
                width23 = 3'b001;
                width22 = 3'b001;
                width21 = 3'b001;
                width20 = 3'b001;
                width19 = 3'b001;
                width18 = 3'b001;
                width17 = 3'b001;
                width16 = 3'b001;
                width15 = 3'b001;
                width14 = 3'b001;
                width13 = 3'b001;
                width12 = 3'b001;
                width11 = 3'b001;
                width10 = 3'b001;
                width9 = 3'b001;
                width8 = 3'b010;
                width7 = 3'b010;
                width6 = 3'b010;
                width5 = 3'b010;
                width4 = 3'b010;
                width3 = 3'b010;
                width2 = 3'b010;
                width1 = 3'b010;

                writeAddr56 = {writeAddr[13:0]};
                writeAddr55 = {writeAddr[13:0]};
                writeAddr54 = {writeAddr[13:0]};
                writeAddr53 = {writeAddr[13:0]};
                writeAddr52 = {writeAddr[13:0]};
                writeAddr51 = {writeAddr[13:0]};
                writeAddr50 = {writeAddr[13:0]};
                writeAddr49 = {writeAddr[13:0]};
                writeAddr48 = {writeAddr[13:0]};
                writeAddr47 = {writeAddr[13:0]};
                writeAddr46 = {writeAddr[13:0]};
                writeAddr45 = {writeAddr[13:0]};
                writeAddr44 = {writeAddr[13:0]};
                writeAddr43 = {writeAddr[13:0]};
                writeAddr42 = {writeAddr[13:0]};
                writeAddr41 = {writeAddr[13:0]};
                writeAddr40 = {writeAddr[13:0]};
                writeAddr39 = {writeAddr[13:0]};
                writeAddr38 = {writeAddr[13:0]};
                writeAddr37 = {writeAddr[13:0]};
                writeAddr36 = {writeAddr[13:0]};
                writeAddr35 = {writeAddr[13:0]};
                writeAddr34 = {writeAddr[13:0]};
                writeAddr33 = {writeAddr[13:0]};
                writeAddr32 = {writeAddr[13:0]};
                writeAddr31 = {writeAddr[13:0]};
                writeAddr30 = {writeAddr[13:0]};
                writeAddr29 = {writeAddr[13:0]};
                writeAddr28 = {writeAddr[13:0]};
                writeAddr27 = {writeAddr[13:0]};
                writeAddr26 = {writeAddr[13:0]};
                writeAddr25 = {writeAddr[13:0]};
                writeAddr24 = {writeAddr[12:0], 1'b0};
                writeAddr23 = {writeAddr[12:0], 1'b0};
                writeAddr22 = {writeAddr[12:0], 1'b0};
                writeAddr21 = {writeAddr[12:0], 1'b0};
                writeAddr20 = {writeAddr[12:0], 1'b0};
                writeAddr19 = {writeAddr[12:0], 1'b0};
                writeAddr18 = {writeAddr[12:0], 1'b0};
                writeAddr17 = {writeAddr[12:0], 1'b0};
                writeAddr16 = {writeAddr[12:0], 1'b0};
                writeAddr15 = {writeAddr[12:0], 1'b0};
                writeAddr14 = {writeAddr[12:0], 1'b0};
                writeAddr13 = {writeAddr[12:0], 1'b0};
                writeAddr12 = {writeAddr[12:0], 1'b0};
                writeAddr11 = {writeAddr[12:0], 1'b0};
                writeAddr10 = {writeAddr[12:0], 1'b0};
                writeAddr9 = {writeAddr[12:0], 1'b0};
                writeAddr8 = {writeAddr[11:0], 2'b0};
                writeAddr7 = {writeAddr[11:0], 2'b0};
                writeAddr6 = {writeAddr[11:0], 2'b0};
                writeAddr5 = {writeAddr[11:0], 2'b0};
                writeAddr4 = {writeAddr[11:0], 2'b0};
                writeAddr3 = {writeAddr[11:0], 2'b0};
                writeAddr2 = {writeAddr[11:0], 2'b0};
                writeAddr1 = {writeAddr[11:0], 2'b0};

                readAddr56 = {writeAddr[13:0]};
                readAddr55 = {writeAddr[13:0]};
                readAddr54 = {writeAddr[13:0]};
                readAddr53 = {writeAddr[13:0]};
                readAddr52 = {writeAddr[13:0]};
                readAddr51 = {writeAddr[13:0]};
                readAddr50 = {writeAddr[13:0]};
                readAddr49 = {writeAddr[13:0]};
                readAddr48 = {writeAddr[13:0]};
                readAddr47 = {writeAddr[13:0]};
                readAddr46 = {writeAddr[13:0]};
                readAddr45 = {writeAddr[13:0]};
                readAddr44 = {writeAddr[13:0]};
                readAddr43 = {writeAddr[13:0]};
                readAddr42 = {writeAddr[13:0]};
                readAddr41 = {writeAddr[13:0]};
                readAddr40 = {writeAddr[13:0]};
                readAddr39 = {writeAddr[13:0]};
                readAddr38 = {writeAddr[13:0]};
                readAddr37 = {writeAddr[13:0]};
                readAddr36 = {writeAddr[13:0]};
                readAddr35 = {writeAddr[13:0]};
                readAddr34 = {writeAddr[13:0]};
                readAddr33 = {writeAddr[13:0]};
                readAddr32 = {writeAddr[13:0]};
                readAddr31 = {writeAddr[13:0]};
                readAddr30 = {writeAddr[13:0]};
                readAddr29 = {writeAddr[13:0]};
                readAddr28 = {writeAddr[13:0]};
                readAddr27 = {writeAddr[13:0]};
                readAddr26 = {writeAddr[13:0]};
                readAddr25 = {writeAddr[13:0]};
                readAddr24  = {readAddr[12:0],  1'b0};
                readAddr23  = {readAddr[12:0],  1'b0};
                readAddr22  = {readAddr[12:0],  1'b0};
                readAddr21  = {readAddr[12:0],  1'b0};
                readAddr20  = {readAddr[12:0],  1'b0};
                readAddr19  = {readAddr[12:0],  1'b0};
                readAddr18  = {readAddr[12:0],  1'b0};
                readAddr17  = {readAddr[12:0],  1'b0};
                readAddr16  = {readAddr[12:0],  1'b0};
                readAddr15  = {readAddr[12:0],  1'b0};
                readAddr14  = {readAddr[12:0],  1'b0};
                readAddr13  = {readAddr[12:0],  1'b0};
                readAddr12  = {readAddr[12:0],  1'b0};
                readAddr11  = {readAddr[12:0],  1'b0};
                readAddr10  = {readAddr[12:0],  1'b0};
                readAddr9  = {readAddr[12:0],  1'b0};
                readAddr8  = {readAddr[11:0],  2'b0};
                readAddr7  = {readAddr[11:0],  2'b0};
                readAddr6  = {readAddr[11:0],  2'b0};
                readAddr5  = {readAddr[11:0],  2'b0};
                readAddr4  = {readAddr[11:0],  2'b0};
                readAddr3  = {readAddr[11:0],  2'b0};
                readAddr2  = {readAddr[11:0],  2'b0};
                readAddr1  = {readAddr[11:0],  2'b0};

                writeData56 = {17'b0, writeData[31]};
                writeData55 = {17'b0, writeData[30]};
                writeData54 = {17'b0, writeData[29]};
                writeData53 = {17'b0, writeData[28]};
                writeData52 = {17'b0, writeData[27]};
                writeData51 = {17'b0, writeData[26]};
                writeData50 = {17'b0, writeData[25]};
                writeData49 = {17'b0, writeData[24]};
                writeData48 = {17'b0, writeData[23]};
                writeData47 = {17'b0, writeData[22]};
                writeData46 = {17'b0, writeData[21]};
                writeData45 = {17'b0, writeData[20]};
                writeData44 = {17'b0, writeData[19]};
                writeData43 = {17'b0, writeData[18]};
                writeData42 = {17'b0, writeData[17]};
                writeData41 = {17'b0, writeData[16]};
                writeData40 = {17'b0, writeData[15]};
                writeData39 = {17'b0, writeData[14]};
                writeData38 = {17'b0, writeData[13]};
                writeData37 = {17'b0, writeData[12]};
                writeData36 = {17'b0, writeData[11]};
                writeData35 = {17'b0, writeData[10]};
                writeData34 = {17'b0, writeData[9]};
                writeData33 = {17'b0, writeData[8]};
                writeData32 = {17'b0, writeData[7]};
                writeData31 = {17'b0, writeData[6]};
                writeData30 = {17'b0, writeData[5]};
                writeData29 = {17'b0, writeData[4]};
                writeData28 = {17'b0, writeData[3]};
                writeData27 = {17'b0, writeData[2]};
                writeData26 = {17'b0, writeData[1]};
                writeData25 = {17'b0, writeData[0]};
                writeData24 = {16'b0, writeData[31:30]};
                writeData23 = {16'b0, writeData[29:28]};
                writeData22 = {16'b0, writeData[27:26]};
                writeData21 = {16'b0, writeData[25:24]};
                writeData20 = {16'b0, writeData[23:22]};
                writeData19 = {16'b0, writeData[21:20]};
                writeData18 = {16'b0, writeData[19:18]};
                writeData17 = {16'b0, writeData[17:16]};
                writeData16 = {16'b0, writeData[15:14]};
                writeData15 = {16'b0, writeData[13:12]};
                writeData14 = {16'b0, writeData[11:10]};
                writeData13 = {16'b0, writeData[9:8]};
                writeData12 = {16'b0, writeData[7:6]};
                writeData11 = {16'b0, writeData[5:4]};
                writeData10 = {16'b0, writeData[3:2]};
                writeData9 = {16'b0, writeData[1:0]};
                writeData8 = {14'b0, writeData[31:28]};
                writeData7 = {14'b0, writeData[27:24]};
                writeData6 = {14'b0, writeData[23:20]};
                writeData5 = {14'b0, writeData[19:16]};
                writeData4 = {14'b0, writeData[15:12]};
                writeData3 = {14'b0, writeData[11:8]};
                writeData2 = {14'b0, writeData[7:4]};
                writeData1 = {14'b0, writeData[3:0]};

                case (writeAddr[14:9])
                    6'b000000, 6'b000001, 6'b000010, 6'b000011,
                    6'b000100, 6'b000101, 6'b000110, 6'b000111,
                    6'b001000, 6'b001001, 6'b001010, 6'b001011,
                    6'b001100, 6'b001101, 6'b001110, 6'b001111,
                    6'b010000, 6'b010001, 6'b010010, 6'b010011,
                    6'b010100, 6'b010101, 6'b010110, 6'b010111,
                    6'b011000, 6'b011001, 6'b011010, 6'b011011,
                    6'b011100, 6'b011101, 6'b011110, 6'b011111 : begin
                        wen_a56 = {1'b0, wen};
                        wen_a55 = {1'b0, wen};
                        wen_a54 = {1'b0, wen};
                        wen_a53 = {1'b0, wen};
                        wen_a52 = {1'b0, wen};
                        wen_a51 = {1'b0, wen};
                        wen_a50 = {1'b0, wen};
                        wen_a49 = {1'b0, wen};
                        wen_a48 = {1'b0, wen};
                        wen_a47 = {1'b0, wen};
                        wen_a46 = {1'b0, wen};
                        wen_a45 = {1'b0, wen};
                        wen_a44 = {1'b0, wen};
                        wen_a43 = {1'b0, wen};
                        wen_a42 = {1'b0, wen};
                        wen_a41 = {1'b0, wen};
                        wen_a40 = {1'b0, wen};
                        wen_a39 = {1'b0, wen};
                        wen_a38 = {1'b0, wen};
                        wen_a37 = {1'b0, wen};
                        wen_a36 = {1'b0, wen};
                        wen_a35 = {1'b0, wen};
                        wen_a34 = {1'b0, wen};
                        wen_a33 = {1'b0, wen};
                        wen_a32 = {1'b0, wen};
                        wen_a31 = {1'b0, wen};
                        wen_a30 = {1'b0, wen};
                        wen_a29 = {1'b0, wen};
                        wen_a28 = {1'b0, wen};
                        wen_a27 = {1'b0, wen};
                        wen_a26 = {1'b0, wen};
                        wen_a25 = {1'b0, wen};
                        wen_a24 = {1'b0, 1'b0};
                        wen_a23 = {1'b0, 1'b0};
                        wen_a22 = {1'b0, 1'b0};
                        wen_a21 = {1'b0, 1'b0};
                        wen_a20 = {1'b0, 1'b0};
                        wen_a19 = {1'b0, 1'b0};
                        wen_a18 = {1'b0, 1'b0};
                        wen_a17 = {1'b0, 1'b0};
                        wen_a16 = {1'b0, 1'b0};
                        wen_a15 = {1'b0, 1'b0};
                        wen_a14 = {1'b0, 1'b0};
                        wen_a13 = {1'b0, 1'b0};
                        wen_a12 = {1'b0, 1'b0};
                        wen_a11 = {1'b0, 1'b0};
                        wen_a10 = {1'b0, 1'b0};
                        wen_a9 = {1'b0, 1'b0};
                        wen_a8 = {1'b0, 1'b0};
                        wen_a7 = {1'b0, 1'b0};
                        wen_a6 = {1'b0, 1'b0};
                        wen_a5 = {1'b0, 1'b0};
                        wen_a4 = {1'b0, 1'b0};
                        wen_a3 = {1'b0, 1'b0};
                        wen_a2 = {1'b0, 1'b0};
                        wen_a1 = {1'b0, 1'b0};
                    end
                    6'b100000, 6'b100001, 6'b100010, 6'b100011,
                    6'b100100, 6'b100101, 6'b100110, 6'b100111,
                    6'b101000, 6'b101001, 6'b101010, 6'b101011,
                    6'b101100, 6'b101101, 6'b101110, 6'b101111 : begin
                        wen_a56 = {1'b0, 1'b0};
                        wen_a55 = {1'b0, 1'b0};
                        wen_a54 = {1'b0, 1'b0};
                        wen_a53 = {1'b0, 1'b0};
                        wen_a52 = {1'b0, 1'b0};
                        wen_a51 = {1'b0, 1'b0};
                        wen_a50 = {1'b0, 1'b0};
                        wen_a49 = {1'b0, 1'b0};
                        wen_a48 = {1'b0, 1'b0};
                        wen_a47 = {1'b0, 1'b0};
                        wen_a46 = {1'b0, 1'b0};
                        wen_a45 = {1'b0, 1'b0};
                        wen_a44 = {1'b0, 1'b0};
                        wen_a43 = {1'b0, 1'b0};
                        wen_a42 = {1'b0, 1'b0};
                        wen_a41 = {1'b0, 1'b0};
                        wen_a40 = {1'b0, 1'b0};
                        wen_a39 = {1'b0, 1'b0};
                        wen_a38 = {1'b0, 1'b0};
                        wen_a37 = {1'b0, 1'b0};
                        wen_a36 = {1'b0, 1'b0};
                        wen_a35 = {1'b0, 1'b0};
                        wen_a34 = {1'b0, 1'b0};
                        wen_a33 = {1'b0, 1'b0};
                        wen_a32 = {1'b0, 1'b0};
                        wen_a31 = {1'b0, 1'b0};
                        wen_a30 = {1'b0, 1'b0};
                        wen_a29 = {1'b0, 1'b0};
                        wen_a28 = {1'b0, 1'b0};
                        wen_a27 = {1'b0, 1'b0};
                        wen_a26 = {1'b0, 1'b0};
                        wen_a25 = {1'b0, 1'b0};
                        wen_a24 = {1'b0, wen};
                        wen_a23 = {1'b0, wen};
                        wen_a22 = {1'b0, wen};
                        wen_a21 = {1'b0, wen};
                        wen_a20 = {1'b0, wen};
                        wen_a19 = {1'b0, wen};
                        wen_a18 = {1'b0, wen};
                        wen_a17 = {1'b0, wen};
                        wen_a16 = {1'b0, wen};
                        wen_a15 = {1'b0, wen};
                        wen_a14 = {1'b0, wen};
                        wen_a13 = {1'b0, wen};
                        wen_a12 = {1'b0, wen};
                        wen_a11 = {1'b0, wen};
                        wen_a10 = {1'b0, wen};
                        wen_a9 = {1'b0, wen};
                        wen_a8 = {1'b0, 1'b0};
                        wen_a7 = {1'b0, 1'b0};
                        wen_a6 = {1'b0, 1'b0};
                        wen_a5 = {1'b0, 1'b0};
                        wen_a4 = {1'b0, 1'b0};
                        wen_a3 = {1'b0, 1'b0};
                        wen_a2 = {1'b0, 1'b0};
                        wen_a1 = {1'b0, 1'b0};
                    end
                    6'b110000, 6'b110001, 6'b110010, 6'b110011,
                    6'b110100, 6'b110101, 6'b110110, 6'b110111 : begin
                        wen_a56 = {1'b0, 1'b0};
                        wen_a55 = {1'b0, 1'b0};
                        wen_a54 = {1'b0, 1'b0};
                        wen_a53 = {1'b0, 1'b0};
                        wen_a52 = {1'b0, 1'b0};
                        wen_a51 = {1'b0, 1'b0};
                        wen_a50 = {1'b0, 1'b0};
                        wen_a49 = {1'b0, 1'b0};
                        wen_a48 = {1'b0, 1'b0};
                        wen_a47 = {1'b0, 1'b0};
                        wen_a46 = {1'b0, 1'b0};
                        wen_a45 = {1'b0, 1'b0};
                        wen_a44 = {1'b0, 1'b0};
                        wen_a43 = {1'b0, 1'b0};
                        wen_a42 = {1'b0, 1'b0};
                        wen_a41 = {1'b0, 1'b0};
                        wen_a40 = {1'b0, 1'b0};
                        wen_a39 = {1'b0, 1'b0};
                        wen_a38 = {1'b0, 1'b0};
                        wen_a37 = {1'b0, 1'b0};
                        wen_a36 = {1'b0, 1'b0};
                        wen_a35 = {1'b0, 1'b0};
                        wen_a34 = {1'b0, 1'b0};
                        wen_a33 = {1'b0, 1'b0};
                        wen_a32 = {1'b0, 1'b0};
                        wen_a31 = {1'b0, 1'b0};
                        wen_a30 = {1'b0, 1'b0};
                        wen_a29 = {1'b0, 1'b0};
                        wen_a28 = {1'b0, 1'b0};
                        wen_a27 = {1'b0, 1'b0};
                        wen_a26 = {1'b0, 1'b0};
                        wen_a25 = {1'b0, 1'b0};
                        wen_a24 = {1'b0, 1'b0};
                        wen_a23 = {1'b0, 1'b0};
                        wen_a22 = {1'b0, 1'b0};
                        wen_a21 = {1'b0, 1'b0};
                        wen_a20 = {1'b0, 1'b0};
                        wen_a19 = {1'b0, 1'b0};
                        wen_a18 = {1'b0, 1'b0};
                        wen_a17 = {1'b0, 1'b0};
                        wen_a16 = {1'b0, 1'b0};
                        wen_a15 = {1'b0, 1'b0};
                        wen_a14 = {1'b0, 1'b0};
                        wen_a13 = {1'b0, 1'b0};
                        wen_a12 = {1'b0, 1'b0};
                        wen_a11 = {1'b0, 1'b0};
                        wen_a10 = {1'b0, 1'b0};
                        wen_a9 = {1'b0, 1'b0};
                        wen_a8 = {1'b0, wen};
                        wen_a7 = {1'b0, wen};
                        wen_a6 = {1'b0, wen};
                        wen_a5 = {1'b0, wen};
                        wen_a4 = {1'b0, wen};
                        wen_a3 = {1'b0, wen};
                        wen_a2 = {1'b0, wen};
                        wen_a1 = {1'b0, wen};
                    end
                    default : begin
                        wen_a56 = {1'b0, 1'b0};
                        wen_a55 = {1'b0, 1'b0};
                        wen_a54 = {1'b0, 1'b0};
                        wen_a53 = {1'b0, 1'b0};
                        wen_a52 = {1'b0, 1'b0};
                        wen_a51 = {1'b0, 1'b0};
                        wen_a50 = {1'b0, 1'b0};
                        wen_a49 = {1'b0, 1'b0};
                        wen_a48 = {1'b0, 1'b0};
                        wen_a47 = {1'b0, 1'b0};
                        wen_a46 = {1'b0, 1'b0};
                        wen_a45 = {1'b0, 1'b0};
                        wen_a44 = {1'b0, 1'b0};
                        wen_a43 = {1'b0, 1'b0};
                        wen_a42 = {1'b0, 1'b0};
                        wen_a41 = {1'b0, 1'b0};
                        wen_a40 = {1'b0, 1'b0};
                        wen_a39 = {1'b0, 1'b0};
                        wen_a38 = {1'b0, 1'b0};
                        wen_a37 = {1'b0, 1'b0};
                        wen_a36 = {1'b0, 1'b0};
                        wen_a35 = {1'b0, 1'b0};
                        wen_a34 = {1'b0, 1'b0};
                        wen_a33 = {1'b0, 1'b0};
                        wen_a32 = {1'b0, 1'b0};
                        wen_a31 = {1'b0, 1'b0};
                        wen_a30 = {1'b0, 1'b0};
                        wen_a29 = {1'b0, 1'b0};
                        wen_a28 = {1'b0, 1'b0};
                        wen_a27 = {1'b0, 1'b0};
                        wen_a26 = {1'b0, 1'b0};
                        wen_a25 = {1'b0, 1'b0};
                        wen_a24 = {1'b0, 1'b0};
                        wen_a23 = {1'b0, 1'b0};
                        wen_a22 = {1'b0, 1'b0};
                        wen_a21 = {1'b0, 1'b0};
                        wen_a20 = {1'b0, 1'b0};
                        wen_a19 = {1'b0, 1'b0};
                        wen_a18 = {1'b0, 1'b0};
                        wen_a17 = {1'b0, 1'b0};
                        wen_a16 = {1'b0, 1'b0};
                        wen_a15 = {1'b0, 1'b0};
                        wen_a14 = {1'b0, 1'b0};
                        wen_a13 = {1'b0, 1'b0};
                        wen_a12 = {1'b0, 1'b0};
                        wen_a11 = {1'b0, 1'b0};
                        wen_a10 = {1'b0, 1'b0};
                        wen_a9 = {1'b0, 1'b0};
                        wen_a8 = {1'b0, 1'b0};
                        wen_a7 = {1'b0, 1'b0};
                        wen_a6 = {1'b0, 1'b0};
                        wen_a5 = {1'b0, 1'b0};
                        wen_a4 = {1'b0, 1'b0};
                        wen_a3 = {1'b0, 1'b0};
                        wen_a2 = {1'b0, 1'b0};
                        wen_a1 = {1'b0, 1'b0};
                    end
                endcase

                case (ckRdAddr[14:9])
                    6'b000000, 6'b000001, 6'b000010, 6'b000011,
                    6'b000100, 6'b000101, 6'b000110, 6'b000111,
                    6'b001000, 6'b001001, 6'b001010, 6'b001011,
                    6'b001100, 6'b001101, 6'b001110, 6'b001111,
                    6'b010000, 6'b010001, 6'b010010, 6'b010011,
                    6'b010100, 6'b010101, 6'b010110, 6'b010111,
                    6'b011000, 6'b011001, 6'b011010, 6'b011011,
                    6'b011100, 6'b011101, 6'b011110, 6'b011111 : begin
                        readData = {
                                        readData56[0],
                                        readData55[0],
                                        readData54[0],
                                        readData53[0],
                                        readData52[0],
                                        readData51[0],
                                        readData50[0],
                                        readData49[0],
                                        readData48[0],
                                        readData47[0],
                                        readData46[0],
                                        readData45[0],
                                        readData44[0],
                                        readData43[0],
                                        readData42[0],
                                        readData41[0],
                                        readData40[0],
                                        readData39[0],
                                        readData38[0],
                                        readData37[0],
                                        readData36[0],
                                        readData35[0],
                                        readData34[0],
                                        readData33[0],
                                        readData32[0],
                                        readData31[0],
                                        readData30[0],
                                        readData29[0],
                                        readData28[0],
                                        readData27[0],
                                        readData26[0],
                                        readData25[0]
                        };
                    end
                    6'b100000, 6'b100001, 6'b100010, 6'b100011,
                    6'b100100, 6'b100101, 6'b100110, 6'b100111,
                    6'b101000, 6'b101001, 6'b101010, 6'b101011,
                    6'b101100, 6'b101101, 6'b101110, 6'b101111 : begin
                        readData = {
                                        readData24[1:0],
                                        readData23[1:0],
                                        readData22[1:0],
                                        readData21[1:0],
                                        readData20[1:0],
                                        readData19[1:0],
                                        readData18[1:0],
                                        readData17[1:0],
                                        readData16[1:0],
                                        readData15[1:0],
                                        readData14[1:0],
                                        readData13[1:0],
                                        readData12[1:0],
                                        readData11[1:0],
                                        readData10[1:0],
                                        readData9[1:0]
                        };
                    end
                    6'b110000, 6'b110001, 6'b110010, 6'b110011,
                    6'b110100, 6'b110101, 6'b110110, 6'b110111 : begin
                        readData = {
                                        readData8[3:0],
                                        readData7[3:0],
                                        readData6[3:0],
                                        readData5[3:0],
                                        readData4[3:0],
                                        readData3[3:0],
                                        readData2[3:0],
                                        readData1[3:0]
                        };
                    end
                    default : begin
                        readData = 32'b0;
                    end
                endcase
            end        
            29184: begin
                width56 = 3'b000;
                width55 = 3'b000;
                width54 = 3'b000;
                width53 = 3'b000;
                width52 = 3'b000;
                width51 = 3'b000;
                width50 = 3'b000;
                width49 = 3'b000;
                width48 = 3'b000;
                width47 = 3'b000;
                width46 = 3'b000;
                width45 = 3'b000;
                width44 = 3'b000;
                width43 = 3'b000;
                width42 = 3'b000;
                width41 = 3'b000;
                width40 = 3'b000;
                width39 = 3'b000;
                width38 = 3'b000;
                width37 = 3'b000;
                width36 = 3'b000;
                width35 = 3'b000;
                width34 = 3'b000;
                width33 = 3'b000;
                width32 = 3'b000;
                width31 = 3'b000;
                width30 = 3'b000;
                width29 = 3'b000;
                width28 = 3'b000;
                width27 = 3'b000;
                width26 = 3'b000;
                width25 = 3'b000;
                width24 = 3'b001;
                width23 = 3'b001;
                width22 = 3'b001;
                width21 = 3'b001;
                width20 = 3'b001;
                width19 = 3'b001;
                width18 = 3'b001;
                width17 = 3'b001;
                width16 = 3'b001;
                width15 = 3'b001;
                width14 = 3'b001;
                width13 = 3'b001;
                width12 = 3'b001;
                width11 = 3'b001;
                width10 = 3'b001;
                width9 = 3'b001;
                width8 = 3'b010;
                width7 = 3'b010;
                width6 = 3'b010;
                width5 = 3'b010;
                width4 = 3'b010;
                width3 = 3'b010;
                width2 = 3'b010;
                width1 = 3'b010;
                width0 = 3'b101;

                writeAddr56 = {writeAddr[13:0]};
                writeAddr55 = {writeAddr[13:0]};
                writeAddr54 = {writeAddr[13:0]};
                writeAddr53 = {writeAddr[13:0]};
                writeAddr52 = {writeAddr[13:0]};
                writeAddr51 = {writeAddr[13:0]};
                writeAddr50 = {writeAddr[13:0]};
                writeAddr49 = {writeAddr[13:0]};
                writeAddr48 = {writeAddr[13:0]};
                writeAddr47 = {writeAddr[13:0]};
                writeAddr46 = {writeAddr[13:0]};
                writeAddr45 = {writeAddr[13:0]};
                writeAddr44 = {writeAddr[13:0]};
                writeAddr43 = {writeAddr[13:0]};
                writeAddr42 = {writeAddr[13:0]};
                writeAddr41 = {writeAddr[13:0]};
                writeAddr40 = {writeAddr[13:0]};
                writeAddr39 = {writeAddr[13:0]};
                writeAddr38 = {writeAddr[13:0]};
                writeAddr37 = {writeAddr[13:0]};
                writeAddr36 = {writeAddr[13:0]};
                writeAddr35 = {writeAddr[13:0]};
                writeAddr34 = {writeAddr[13:0]};
                writeAddr33 = {writeAddr[13:0]};
                writeAddr32 = {writeAddr[13:0]};
                writeAddr31 = {writeAddr[13:0]};
                writeAddr30 = {writeAddr[13:0]};
                writeAddr29 = {writeAddr[13:0]};
                writeAddr28 = {writeAddr[13:0]};
                writeAddr27 = {writeAddr[13:0]};
                writeAddr26 = {writeAddr[13:0]};
                writeAddr25 = {writeAddr[13:0]};
                writeAddr24 = {writeAddr[12:0], 1'b0};
                writeAddr23 = {writeAddr[12:0], 1'b0};
                writeAddr22 = {writeAddr[12:0], 1'b0};
                writeAddr21 = {writeAddr[12:0], 1'b0};
                writeAddr20 = {writeAddr[12:0], 1'b0};
                writeAddr19 = {writeAddr[12:0], 1'b0};
                writeAddr18 = {writeAddr[12:0], 1'b0};
                writeAddr17 = {writeAddr[12:0], 1'b0};
                writeAddr16 = {writeAddr[12:0], 1'b0};
                writeAddr15 = {writeAddr[12:0], 1'b0};
                writeAddr14 = {writeAddr[12:0], 1'b0};
                writeAddr13 = {writeAddr[12:0], 1'b0};
                writeAddr12 = {writeAddr[12:0], 1'b0};
                writeAddr11 = {writeAddr[12:0], 1'b0};
                writeAddr10 = {writeAddr[12:0], 1'b0};
                writeAddr9 = {writeAddr[12:0], 1'b0};
                writeAddr8 = {writeAddr[11:0], 2'b0};
                writeAddr7 = {writeAddr[11:0], 2'b0};
                writeAddr6 = {writeAddr[11:0], 2'b0};
                writeAddr5 = {writeAddr[11:0], 2'b0};
                writeAddr4 = {writeAddr[11:0], 2'b0};
                writeAddr3 = {writeAddr[11:0], 2'b0};
                writeAddr2 = {writeAddr[11:0], 2'b0};
                writeAddr1 = {writeAddr[11:0], 2'b0};
                writeAddr0 = {writeAddr[8:0], 5'b0};

                readAddr56 = {writeAddr[13:0]};
                readAddr55 = {writeAddr[13:0]};
                readAddr54 = {writeAddr[13:0]};
                readAddr53 = {writeAddr[13:0]};
                readAddr52 = {writeAddr[13:0]};
                readAddr51 = {writeAddr[13:0]};
                readAddr50 = {writeAddr[13:0]};
                readAddr49 = {writeAddr[13:0]};
                readAddr48 = {writeAddr[13:0]};
                readAddr47 = {writeAddr[13:0]};
                readAddr46 = {writeAddr[13:0]};
                readAddr45 = {writeAddr[13:0]};
                readAddr44 = {writeAddr[13:0]};
                readAddr43 = {writeAddr[13:0]};
                readAddr42 = {writeAddr[13:0]};
                readAddr41 = {writeAddr[13:0]};
                readAddr40 = {writeAddr[13:0]};
                readAddr39 = {writeAddr[13:0]};
                readAddr38 = {writeAddr[13:0]};
                readAddr37 = {writeAddr[13:0]};
                readAddr36 = {writeAddr[13:0]};
                readAddr35 = {writeAddr[13:0]};
                readAddr34 = {writeAddr[13:0]};
                readAddr33 = {writeAddr[13:0]};
                readAddr32 = {writeAddr[13:0]};
                readAddr31 = {writeAddr[13:0]};
                readAddr30 = {writeAddr[13:0]};
                readAddr29 = {writeAddr[13:0]};
                readAddr28 = {writeAddr[13:0]};
                readAddr27 = {writeAddr[13:0]};
                readAddr26 = {writeAddr[13:0]};
                readAddr25 = {writeAddr[13:0]};
                readAddr24  = {readAddr[12:0],  1'b0};
                readAddr23  = {readAddr[12:0],  1'b0};
                readAddr22  = {readAddr[12:0],  1'b0};
                readAddr21  = {readAddr[12:0],  1'b0};
                readAddr20  = {readAddr[12:0],  1'b0};
                readAddr19  = {readAddr[12:0],  1'b0};
                readAddr18  = {readAddr[12:0],  1'b0};
                readAddr17  = {readAddr[12:0],  1'b0};
                readAddr16  = {readAddr[12:0],  1'b0};
                readAddr15  = {readAddr[12:0],  1'b0};
                readAddr14  = {readAddr[12:0],  1'b0};
                readAddr13  = {readAddr[12:0],  1'b0};
                readAddr12  = {readAddr[12:0],  1'b0};
                readAddr11  = {readAddr[12:0],  1'b0};
                readAddr10  = {readAddr[12:0],  1'b0};
                readAddr9  = {readAddr[12:0],  1'b0};
                readAddr8  = {readAddr[11:0],  2'b0};
                readAddr7  = {readAddr[11:0],  2'b0};
                readAddr6  = {readAddr[11:0],  2'b0};
                readAddr5  = {readAddr[11:0],  2'b0};
                readAddr4  = {readAddr[11:0],  2'b0};
                readAddr3  = {readAddr[11:0],  2'b0};
                readAddr2  = {readAddr[11:0],  2'b0};
                readAddr1  = {readAddr[11:0],  2'b0};
                readAddr0  = {readAddr[8:0],  5'b0};

                writeData56 = {17'b0, writeData[31]};
                writeData55 = {17'b0, writeData[30]};
                writeData54 = {17'b0, writeData[29]};
                writeData53 = {17'b0, writeData[28]};
                writeData52 = {17'b0, writeData[27]};
                writeData51 = {17'b0, writeData[26]};
                writeData50 = {17'b0, writeData[25]};
                writeData49 = {17'b0, writeData[24]};
                writeData48 = {17'b0, writeData[23]};
                writeData47 = {17'b0, writeData[22]};
                writeData46 = {17'b0, writeData[21]};
                writeData45 = {17'b0, writeData[20]};
                writeData44 = {17'b0, writeData[19]};
                writeData43 = {17'b0, writeData[18]};
                writeData42 = {17'b0, writeData[17]};
                writeData41 = {17'b0, writeData[16]};
                writeData40 = {17'b0, writeData[15]};
                writeData39 = {17'b0, writeData[14]};
                writeData38 = {17'b0, writeData[13]};
                writeData37 = {17'b0, writeData[12]};
                writeData36 = {17'b0, writeData[11]};
                writeData35 = {17'b0, writeData[10]};
                writeData34 = {17'b0, writeData[9]};
                writeData33 = {17'b0, writeData[8]};
                writeData32 = {17'b0, writeData[7]};
                writeData31 = {17'b0, writeData[6]};
                writeData30 = {17'b0, writeData[5]};
                writeData29 = {17'b0, writeData[4]};
                writeData28 = {17'b0, writeData[3]};
                writeData27 = {17'b0, writeData[2]};
                writeData26 = {17'b0, writeData[1]};
                writeData25 = {17'b0, writeData[0]};
                writeData24 = {16'b0, writeData[31:30]};
                writeData23 = {16'b0, writeData[29:28]};
                writeData22 = {16'b0, writeData[27:26]};
                writeData21 = {16'b0, writeData[25:24]};
                writeData20 = {16'b0, writeData[23:22]};
                writeData19 = {16'b0, writeData[21:20]};
                writeData18 = {16'b0, writeData[19:18]};
                writeData17 = {16'b0, writeData[17:16]};
                writeData16 = {16'b0, writeData[15:14]};
                writeData15 = {16'b0, writeData[13:12]};
                writeData14 = {16'b0, writeData[11:10]};
                writeData13 = {16'b0, writeData[9:8]};
                writeData12 = {16'b0, writeData[7:6]};
                writeData11 = {16'b0, writeData[5:4]};
                writeData10 = {16'b0, writeData[3:2]};
                writeData9 = {16'b0, writeData[1:0]};
                writeData8 = {14'b0, writeData[31:28]};
                writeData7 = {14'b0, writeData[27:24]};
                writeData6 = {14'b0, writeData[23:20]};
                writeData5 = {14'b0, writeData[19:16]};
                writeData4 = {14'b0, writeData[15:12]};
                writeData3 = {14'b0, writeData[11:8]};
                writeData2 = {14'b0, writeData[7:4]};
                writeData1 = {14'b0, writeData[3:0]};
                writeData0 = {1'b0, writeData[31:24], 1'b0, writeData[23:16], 1'b0, writeData[15:8], 1'b0, writeData[7:0]};

                case (writeAddr[14:9])
                    6'b000000, 6'b000001, 6'b000010, 6'b000011,
                    6'b000100, 6'b000101, 6'b000110, 6'b000111,
                    6'b001000, 6'b001001, 6'b001010, 6'b001011,
                    6'b001100, 6'b001101, 6'b001110, 6'b001111,
                    6'b010000, 6'b010001, 6'b010010, 6'b010011,
                    6'b010100, 6'b010101, 6'b010110, 6'b010111,
                    6'b011000, 6'b011001, 6'b011010, 6'b011011,
                    6'b011100, 6'b011101, 6'b011110, 6'b011111 : begin
                        wen_a56 = {1'b0, wen};
                        wen_a55 = {1'b0, wen};
                        wen_a54 = {1'b0, wen};
                        wen_a53 = {1'b0, wen};
                        wen_a52 = {1'b0, wen};
                        wen_a51 = {1'b0, wen};
                        wen_a50 = {1'b0, wen};
                        wen_a49 = {1'b0, wen};
                        wen_a48 = {1'b0, wen};
                        wen_a47 = {1'b0, wen};
                        wen_a46 = {1'b0, wen};
                        wen_a45 = {1'b0, wen};
                        wen_a44 = {1'b0, wen};
                        wen_a43 = {1'b0, wen};
                        wen_a42 = {1'b0, wen};
                        wen_a41 = {1'b0, wen};
                        wen_a40 = {1'b0, wen};
                        wen_a39 = {1'b0, wen};
                        wen_a38 = {1'b0, wen};
                        wen_a37 = {1'b0, wen};
                        wen_a36 = {1'b0, wen};
                        wen_a35 = {1'b0, wen};
                        wen_a34 = {1'b0, wen};
                        wen_a33 = {1'b0, wen};
                        wen_a32 = {1'b0, wen};
                        wen_a31 = {1'b0, wen};
                        wen_a30 = {1'b0, wen};
                        wen_a29 = {1'b0, wen};
                        wen_a28 = {1'b0, wen};
                        wen_a27 = {1'b0, wen};
                        wen_a26 = {1'b0, wen};
                        wen_a25 = {1'b0, wen};
                        wen_a24 = {1'b0, 1'b0};
                        wen_a23 = {1'b0, 1'b0};
                        wen_a22 = {1'b0, 1'b0};
                        wen_a21 = {1'b0, 1'b0};
                        wen_a20 = {1'b0, 1'b0};
                        wen_a19 = {1'b0, 1'b0};
                        wen_a18 = {1'b0, 1'b0};
                        wen_a17 = {1'b0, 1'b0};
                        wen_a16 = {1'b0, 1'b0};
                        wen_a15 = {1'b0, 1'b0};
                        wen_a14 = {1'b0, 1'b0};
                        wen_a13 = {1'b0, 1'b0};
                        wen_a12 = {1'b0, 1'b0};
                        wen_a11 = {1'b0, 1'b0};
                        wen_a10 = {1'b0, 1'b0};
                        wen_a9 = {1'b0, 1'b0};
                        wen_a8 = {1'b0, 1'b0};
                        wen_a7 = {1'b0, 1'b0};
                        wen_a6 = {1'b0, 1'b0};
                        wen_a5 = {1'b0, 1'b0};
                        wen_a4 = {1'b0, 1'b0};
                        wen_a3 = {1'b0, 1'b0};
                        wen_a2 = {1'b0, 1'b0};
                        wen_a1 = {1'b0, 1'b0};
                        wen_a0 = {1'b0, 1'b0};
                        wen_b0 = {1'b0, 1'b0};
                    end
                    6'b100000, 6'b100001, 6'b100010, 6'b100011,
                    6'b100100, 6'b100101, 6'b100110, 6'b100111,
                    6'b101000, 6'b101001, 6'b101010, 6'b101011,
                    6'b101100, 6'b101101, 6'b101110, 6'b101111 : begin
                        wen_a56 = {1'b0, 1'b0};
                        wen_a55 = {1'b0, 1'b0};
                        wen_a54 = {1'b0, 1'b0};
                        wen_a53 = {1'b0, 1'b0};
                        wen_a52 = {1'b0, 1'b0};
                        wen_a51 = {1'b0, 1'b0};
                        wen_a50 = {1'b0, 1'b0};
                        wen_a49 = {1'b0, 1'b0};
                        wen_a48 = {1'b0, 1'b0};
                        wen_a47 = {1'b0, 1'b0};
                        wen_a46 = {1'b0, 1'b0};
                        wen_a45 = {1'b0, 1'b0};
                        wen_a44 = {1'b0, 1'b0};
                        wen_a43 = {1'b0, 1'b0};
                        wen_a42 = {1'b0, 1'b0};
                        wen_a41 = {1'b0, 1'b0};
                        wen_a40 = {1'b0, 1'b0};
                        wen_a39 = {1'b0, 1'b0};
                        wen_a38 = {1'b0, 1'b0};
                        wen_a37 = {1'b0, 1'b0};
                        wen_a36 = {1'b0, 1'b0};
                        wen_a35 = {1'b0, 1'b0};
                        wen_a34 = {1'b0, 1'b0};
                        wen_a33 = {1'b0, 1'b0};
                        wen_a32 = {1'b0, 1'b0};
                        wen_a31 = {1'b0, 1'b0};
                        wen_a30 = {1'b0, 1'b0};
                        wen_a29 = {1'b0, 1'b0};
                        wen_a28 = {1'b0, 1'b0};
                        wen_a27 = {1'b0, 1'b0};
                        wen_a26 = {1'b0, 1'b0};
                        wen_a25 = {1'b0, 1'b0};
                        wen_a24 = {1'b0, wen};
                        wen_a23 = {1'b0, wen};
                        wen_a22 = {1'b0, wen};
                        wen_a21 = {1'b0, wen};
                        wen_a20 = {1'b0, wen};
                        wen_a19 = {1'b0, wen};
                        wen_a18 = {1'b0, wen};
                        wen_a17 = {1'b0, wen};
                        wen_a16 = {1'b0, wen};
                        wen_a15 = {1'b0, wen};
                        wen_a14 = {1'b0, wen};
                        wen_a13 = {1'b0, wen};
                        wen_a12 = {1'b0, wen};
                        wen_a11 = {1'b0, wen};
                        wen_a10 = {1'b0, wen};
                        wen_a9 = {1'b0, wen};
                        wen_a8 = {1'b0, 1'b0};
                        wen_a7 = {1'b0, 1'b0};
                        wen_a6 = {1'b0, 1'b0};
                        wen_a5 = {1'b0, 1'b0};
                        wen_a4 = {1'b0, 1'b0};
                        wen_a3 = {1'b0, 1'b0};
                        wen_a2 = {1'b0, 1'b0};
                        wen_a1 = {1'b0, 1'b0};
                        wen_a0 = {1'b0, 1'b0};
                        wen_b0 = {1'b0, 1'b0};
                    end
                    6'b110000, 6'b110001, 6'b110010, 6'b110011,
                    6'b110100, 6'b110101, 6'b110110, 6'b110111 : begin
                        wen_a56 = {1'b0, 1'b0};
                        wen_a55 = {1'b0, 1'b0};
                        wen_a54 = {1'b0, 1'b0};
                        wen_a53 = {1'b0, 1'b0};
                        wen_a52 = {1'b0, 1'b0};
                        wen_a51 = {1'b0, 1'b0};
                        wen_a50 = {1'b0, 1'b0};
                        wen_a49 = {1'b0, 1'b0};
                        wen_a48 = {1'b0, 1'b0};
                        wen_a47 = {1'b0, 1'b0};
                        wen_a46 = {1'b0, 1'b0};
                        wen_a45 = {1'b0, 1'b0};
                        wen_a44 = {1'b0, 1'b0};
                        wen_a43 = {1'b0, 1'b0};
                        wen_a42 = {1'b0, 1'b0};
                        wen_a41 = {1'b0, 1'b0};
                        wen_a40 = {1'b0, 1'b0};
                        wen_a39 = {1'b0, 1'b0};
                        wen_a38 = {1'b0, 1'b0};
                        wen_a37 = {1'b0, 1'b0};
                        wen_a36 = {1'b0, 1'b0};
                        wen_a35 = {1'b0, 1'b0};
                        wen_a34 = {1'b0, 1'b0};
                        wen_a33 = {1'b0, 1'b0};
                        wen_a32 = {1'b0, 1'b0};
                        wen_a31 = {1'b0, 1'b0};
                        wen_a30 = {1'b0, 1'b0};
                        wen_a29 = {1'b0, 1'b0};
                        wen_a28 = {1'b0, 1'b0};
                        wen_a27 = {1'b0, 1'b0};
                        wen_a26 = {1'b0, 1'b0};
                        wen_a25 = {1'b0, 1'b0};
                        wen_a24 = {1'b0, 1'b0};
                        wen_a23 = {1'b0, 1'b0};
                        wen_a22 = {1'b0, 1'b0};
                        wen_a21 = {1'b0, 1'b0};
                        wen_a20 = {1'b0, 1'b0};
                        wen_a19 = {1'b0, 1'b0};
                        wen_a18 = {1'b0, 1'b0};
                        wen_a17 = {1'b0, 1'b0};
                        wen_a16 = {1'b0, 1'b0};
                        wen_a15 = {1'b0, 1'b0};
                        wen_a14 = {1'b0, 1'b0};
                        wen_a13 = {1'b0, 1'b0};
                        wen_a12 = {1'b0, 1'b0};
                        wen_a11 = {1'b0, 1'b0};
                        wen_a10 = {1'b0, 1'b0};
                        wen_a9 = {1'b0, 1'b0};
                        wen_a8 = {1'b0, wen};
                        wen_a7 = {1'b0, wen};
                        wen_a6 = {1'b0, wen};
                        wen_a5 = {1'b0, wen};
                        wen_a4 = {1'b0, wen};
                        wen_a3 = {1'b0, wen};
                        wen_a2 = {1'b0, wen};
                        wen_a1 = {1'b0, wen};
                        wen_a0 = {1'b0, 1'b0};
                        wen_b0 = {1'b0, 1'b0};
                    end
                    6'b111000 : begin
                        wen_a56 = {1'b0, 1'b0};
                        wen_a55 = {1'b0, 1'b0};
                        wen_a54 = {1'b0, 1'b0};
                        wen_a53 = {1'b0, 1'b0};
                        wen_a52 = {1'b0, 1'b0};
                        wen_a51 = {1'b0, 1'b0};
                        wen_a50 = {1'b0, 1'b0};
                        wen_a49 = {1'b0, 1'b0};
                        wen_a48 = {1'b0, 1'b0};
                        wen_a47 = {1'b0, 1'b0};
                        wen_a46 = {1'b0, 1'b0};
                        wen_a45 = {1'b0, 1'b0};
                        wen_a44 = {1'b0, 1'b0};
                        wen_a43 = {1'b0, 1'b0};
                        wen_a42 = {1'b0, 1'b0};
                        wen_a41 = {1'b0, 1'b0};
                        wen_a40 = {1'b0, 1'b0};
                        wen_a39 = {1'b0, 1'b0};
                        wen_a38 = {1'b0, 1'b0};
                        wen_a37 = {1'b0, 1'b0};
                        wen_a36 = {1'b0, 1'b0};
                        wen_a35 = {1'b0, 1'b0};
                        wen_a34 = {1'b0, 1'b0};
                        wen_a33 = {1'b0, 1'b0};
                        wen_a32 = {1'b0, 1'b0};
                        wen_a31 = {1'b0, 1'b0};
                        wen_a30 = {1'b0, 1'b0};
                        wen_a29 = {1'b0, 1'b0};
                        wen_a28 = {1'b0, 1'b0};
                        wen_a27 = {1'b0, 1'b0};
                        wen_a26 = {1'b0, 1'b0};
                        wen_a25 = {1'b0, 1'b0};
                        wen_a24 = {1'b0, 1'b0};
                        wen_a23 = {1'b0, 1'b0};
                        wen_a22 = {1'b0, 1'b0};
                        wen_a21 = {1'b0, 1'b0};
                        wen_a20 = {1'b0, 1'b0};
                        wen_a19 = {1'b0, 1'b0};
                        wen_a18 = {1'b0, 1'b0};
                        wen_a17 = {1'b0, 1'b0};
                        wen_a16 = {1'b0, 1'b0};
                        wen_a15 = {1'b0, 1'b0};
                        wen_a14 = {1'b0, 1'b0};
                        wen_a13 = {1'b0, 1'b0};
                        wen_a12 = {1'b0, 1'b0};
                        wen_a11 = {1'b0, 1'b0};
                        wen_a10 = {1'b0, 1'b0};
                        wen_a9 = {1'b0, 1'b0};
                        wen_a8 = {1'b0, 1'b0};
                        wen_a7 = {1'b0, 1'b0};
                        wen_a6 = {1'b0, 1'b0};
                        wen_a5 = {1'b0, 1'b0};
                        wen_a4 = {1'b0, 1'b0};
                        wen_a3 = {1'b0, 1'b0};
                        wen_a2 = {1'b0, 1'b0};
                        wen_a1 = {1'b0, 1'b0};
                        wen_a0 = {wen, wen};
                        wen_b0 = {wen, wen};
                    end
                    default : begin
                        wen_a56 = {1'b0, 1'b0};
                        wen_a55 = {1'b0, 1'b0};
                        wen_a54 = {1'b0, 1'b0};
                        wen_a53 = {1'b0, 1'b0};
                        wen_a52 = {1'b0, 1'b0};
                        wen_a51 = {1'b0, 1'b0};
                        wen_a50 = {1'b0, 1'b0};
                        wen_a49 = {1'b0, 1'b0};
                        wen_a48 = {1'b0, 1'b0};
                        wen_a47 = {1'b0, 1'b0};
                        wen_a46 = {1'b0, 1'b0};
                        wen_a45 = {1'b0, 1'b0};
                        wen_a44 = {1'b0, 1'b0};
                        wen_a43 = {1'b0, 1'b0};
                        wen_a42 = {1'b0, 1'b0};
                        wen_a41 = {1'b0, 1'b0};
                        wen_a40 = {1'b0, 1'b0};
                        wen_a39 = {1'b0, 1'b0};
                        wen_a38 = {1'b0, 1'b0};
                        wen_a37 = {1'b0, 1'b0};
                        wen_a36 = {1'b0, 1'b0};
                        wen_a35 = {1'b0, 1'b0};
                        wen_a34 = {1'b0, 1'b0};
                        wen_a33 = {1'b0, 1'b0};
                        wen_a32 = {1'b0, 1'b0};
                        wen_a31 = {1'b0, 1'b0};
                        wen_a30 = {1'b0, 1'b0};
                        wen_a29 = {1'b0, 1'b0};
                        wen_a28 = {1'b0, 1'b0};
                        wen_a27 = {1'b0, 1'b0};
                        wen_a26 = {1'b0, 1'b0};
                        wen_a25 = {1'b0, 1'b0};
                        wen_a24 = {1'b0, 1'b0};
                        wen_a23 = {1'b0, 1'b0};
                        wen_a22 = {1'b0, 1'b0};
                        wen_a21 = {1'b0, 1'b0};
                        wen_a20 = {1'b0, 1'b0};
                        wen_a19 = {1'b0, 1'b0};
                        wen_a18 = {1'b0, 1'b0};
                        wen_a17 = {1'b0, 1'b0};
                        wen_a16 = {1'b0, 1'b0};
                        wen_a15 = {1'b0, 1'b0};
                        wen_a14 = {1'b0, 1'b0};
                        wen_a13 = {1'b0, 1'b0};
                        wen_a12 = {1'b0, 1'b0};
                        wen_a11 = {1'b0, 1'b0};
                        wen_a10 = {1'b0, 1'b0};
                        wen_a9 = {1'b0, 1'b0};
                        wen_a8 = {1'b0, 1'b0};
                        wen_a7 = {1'b0, 1'b0};
                        wen_a6 = {1'b0, 1'b0};
                        wen_a5 = {1'b0, 1'b0};
                        wen_a4 = {1'b0, 1'b0};
                        wen_a3 = {1'b0, 1'b0};
                        wen_a2 = {1'b0, 1'b0};
                        wen_a1 = {1'b0, 1'b0};
                        wen_a0 = {1'b0, 1'b0};
                        wen_b0 = {1'b0, 1'b0};
                    end
                endcase

                case (ckRdAddr[14:9])
                    6'b000000, 6'b000001, 6'b000010, 6'b000011,
                    6'b000100, 6'b000101, 6'b000110, 6'b000111,
                    6'b001000, 6'b001001, 6'b001010, 6'b001011,
                    6'b001100, 6'b001101, 6'b001110, 6'b001111,
                    6'b010000, 6'b010001, 6'b010010, 6'b010011,
                    6'b010100, 6'b010101, 6'b010110, 6'b010111,
                    6'b011000, 6'b011001, 6'b011010, 6'b011011,
                    6'b011100, 6'b011101, 6'b011110, 6'b011111 : begin
                        readData = {
                                        readData56[0],
                                        readData55[0],
                                        readData54[0],
                                        readData53[0],
                                        readData52[0],
                                        readData51[0],
                                        readData50[0],
                                        readData49[0],
                                        readData48[0],
                                        readData47[0],
                                        readData46[0],
                                        readData45[0],
                                        readData44[0],
                                        readData43[0],
                                        readData42[0],
                                        readData41[0],
                                        readData40[0],
                                        readData39[0],
                                        readData38[0],
                                        readData37[0],
                                        readData36[0],
                                        readData35[0],
                                        readData34[0],
                                        readData33[0],
                                        readData32[0],
                                        readData31[0],
                                        readData30[0],
                                        readData29[0],
                                        readData28[0],
                                        readData27[0],
                                        readData26[0],
                                        readData25[0]
                        };
                    end
                    6'b100000, 6'b100001, 6'b100010, 6'b100011,
                    6'b100100, 6'b100101, 6'b100110, 6'b100111,
                    6'b101000, 6'b101001, 6'b101010, 6'b101011,
                    6'b101100, 6'b101101, 6'b101110, 6'b101111 : begin
                        readData = {
                                        readData24[1:0],
                                        readData23[1:0],
                                        readData22[1:0],
                                        readData21[1:0],
                                        readData20[1:0],
                                        readData19[1:0],
                                        readData18[1:0],
                                        readData17[1:0],
                                        readData16[1:0],
                                        readData15[1:0],
                                        readData14[1:0],
                                        readData13[1:0],
                                        readData12[1:0],
                                        readData11[1:0],
                                        readData10[1:0],
                                        readData9[1:0]
                        };
                    end
                    6'b110000, 6'b110001, 6'b110010, 6'b110011,
                    6'b110100, 6'b110101, 6'b110110, 6'b110111 : begin
                        readData = {
                                        readData8[3:0],
                                        readData7[3:0],
                                        readData6[3:0],
                                        readData5[3:0],
                                        readData4[3:0],
                                        readData3[3:0],
                                        readData2[3:0],
                                        readData1[3:0]
                        };
                    end
                    6'b111000 : begin
                        readData = {readData0[34:27],readData0[25:18],readData0[16:9],readData0[7:0]};
                    end
                    default : begin
                        readData = 32'b0;
                    end
                endcase
            end        
            29696: begin
                width58 = 3'b000;
                width57 = 3'b000;
                width56 = 3'b000;
                width55 = 3'b000;
                width54 = 3'b000;
                width53 = 3'b000;
                width52 = 3'b000;
                width51 = 3'b000;
                width50 = 3'b000;
                width49 = 3'b000;
                width48 = 3'b000;
                width47 = 3'b000;
                width46 = 3'b000;
                width45 = 3'b000;
                width44 = 3'b000;
                width43 = 3'b000;
                width42 = 3'b000;
                width41 = 3'b000;
                width40 = 3'b000;
                width39 = 3'b000;
                width38 = 3'b000;
                width37 = 3'b000;
                width36 = 3'b000;
                width35 = 3'b000;
                width34 = 3'b000;
                width33 = 3'b000;
                width32 = 3'b000;
                width31 = 3'b000;
                width30 = 3'b000;
                width29 = 3'b000;
                width28 = 3'b000;
                width27 = 3'b000;
                width26 = 3'b001;
                width25 = 3'b001;
                width24 = 3'b001;
                width23 = 3'b001;
                width22 = 3'b001;
                width21 = 3'b001;
                width20 = 3'b001;
                width19 = 3'b001;
                width18 = 3'b001;
                width17 = 3'b001;
                width16 = 3'b001;
                width15 = 3'b001;
                width14 = 3'b001;
                width13 = 3'b001;
                width12 = 3'b001;
                width11 = 3'b001;
                width10 = 3'b010;
                width9 = 3'b010;
                width8 = 3'b010;
                width7 = 3'b010;
                width6 = 3'b010;
                width5 = 3'b010;
                width4 = 3'b010;
                width3 = 3'b010;
                width2 = 3'b100;
                width1 = 3'b100;

                writeAddr58 = {writeAddr[13:0]};
                writeAddr57 = {writeAddr[13:0]};
                writeAddr56 = {writeAddr[13:0]};
                writeAddr55 = {writeAddr[13:0]};
                writeAddr54 = {writeAddr[13:0]};
                writeAddr53 = {writeAddr[13:0]};
                writeAddr52 = {writeAddr[13:0]};
                writeAddr51 = {writeAddr[13:0]};
                writeAddr50 = {writeAddr[13:0]};
                writeAddr49 = {writeAddr[13:0]};
                writeAddr48 = {writeAddr[13:0]};
                writeAddr47 = {writeAddr[13:0]};
                writeAddr46 = {writeAddr[13:0]};
                writeAddr45 = {writeAddr[13:0]};
                writeAddr44 = {writeAddr[13:0]};
                writeAddr43 = {writeAddr[13:0]};
                writeAddr42 = {writeAddr[13:0]};
                writeAddr41 = {writeAddr[13:0]};
                writeAddr40 = {writeAddr[13:0]};
                writeAddr39 = {writeAddr[13:0]};
                writeAddr38 = {writeAddr[13:0]};
                writeAddr37 = {writeAddr[13:0]};
                writeAddr36 = {writeAddr[13:0]};
                writeAddr35 = {writeAddr[13:0]};
                writeAddr34 = {writeAddr[13:0]};
                writeAddr33 = {writeAddr[13:0]};
                writeAddr32 = {writeAddr[13:0]};
                writeAddr31 = {writeAddr[13:0]};
                writeAddr30 = {writeAddr[13:0]};
                writeAddr29 = {writeAddr[13:0]};
                writeAddr28 = {writeAddr[13:0]};
                writeAddr27 = {writeAddr[13:0]};
                writeAddr26 = {writeAddr[12:0], 1'b0};
                writeAddr25 = {writeAddr[12:0], 1'b0};
                writeAddr24 = {writeAddr[12:0], 1'b0};
                writeAddr23 = {writeAddr[12:0], 1'b0};
                writeAddr22 = {writeAddr[12:0], 1'b0};
                writeAddr21 = {writeAddr[12:0], 1'b0};
                writeAddr20 = {writeAddr[12:0], 1'b0};
                writeAddr19 = {writeAddr[12:0], 1'b0};
                writeAddr18 = {writeAddr[12:0], 1'b0};
                writeAddr17 = {writeAddr[12:0], 1'b0};
                writeAddr16 = {writeAddr[12:0], 1'b0};
                writeAddr15 = {writeAddr[12:0], 1'b0};
                writeAddr14 = {writeAddr[12:0], 1'b0};
                writeAddr13 = {writeAddr[12:0], 1'b0};
                writeAddr12 = {writeAddr[12:0], 1'b0};
                writeAddr11 = {writeAddr[12:0], 1'b0};
                writeAddr10 = {writeAddr[11:0], 2'b0};
                writeAddr9 = {writeAddr[11:0], 2'b0};
                writeAddr8 = {writeAddr[11:0], 2'b0};
                writeAddr7 = {writeAddr[11:0], 2'b0};
                writeAddr6 = {writeAddr[11:0], 2'b0};
                writeAddr5 = {writeAddr[11:0], 2'b0};
                writeAddr4 = {writeAddr[11:0], 2'b0};
                writeAddr3 = {writeAddr[11:0], 2'b0};
                writeAddr2 = {writeAddr[9:0], 4'b0};
                writeAddr1 = {writeAddr[9:0], 4'b0};

                readAddr58 = {writeAddr[13:0]};
                readAddr57 = {writeAddr[13:0]};
                readAddr56 = {writeAddr[13:0]};
                readAddr55 = {writeAddr[13:0]};
                readAddr54 = {writeAddr[13:0]};
                readAddr53 = {writeAddr[13:0]};
                readAddr52 = {writeAddr[13:0]};
                readAddr51 = {writeAddr[13:0]};
                readAddr50 = {writeAddr[13:0]};
                readAddr49 = {writeAddr[13:0]};
                readAddr48 = {writeAddr[13:0]};
                readAddr47 = {writeAddr[13:0]};
                readAddr46 = {writeAddr[13:0]};
                readAddr45 = {writeAddr[13:0]};
                readAddr44 = {writeAddr[13:0]};
                readAddr43 = {writeAddr[13:0]};
                readAddr42 = {writeAddr[13:0]};
                readAddr41 = {writeAddr[13:0]};
                readAddr40 = {writeAddr[13:0]};
                readAddr39 = {writeAddr[13:0]};
                readAddr38 = {writeAddr[13:0]};
                readAddr37 = {writeAddr[13:0]};
                readAddr36 = {writeAddr[13:0]};
                readAddr35 = {writeAddr[13:0]};
                readAddr34 = {writeAddr[13:0]};
                readAddr33 = {writeAddr[13:0]};
                readAddr32 = {writeAddr[13:0]};
                readAddr31 = {writeAddr[13:0]};
                readAddr30 = {writeAddr[13:0]};
                readAddr29 = {writeAddr[13:0]};
                readAddr28 = {writeAddr[13:0]};
                readAddr27 = {writeAddr[13:0]};
                readAddr26  = {readAddr[12:0],  1'b0};
                readAddr25  = {readAddr[12:0],  1'b0};
                readAddr24  = {readAddr[12:0],  1'b0};
                readAddr23  = {readAddr[12:0],  1'b0};
                readAddr22  = {readAddr[12:0],  1'b0};
                readAddr21  = {readAddr[12:0],  1'b0};
                readAddr20  = {readAddr[12:0],  1'b0};
                readAddr19  = {readAddr[12:0],  1'b0};
                readAddr18  = {readAddr[12:0],  1'b0};
                readAddr17  = {readAddr[12:0],  1'b0};
                readAddr16  = {readAddr[12:0],  1'b0};
                readAddr15  = {readAddr[12:0],  1'b0};
                readAddr14  = {readAddr[12:0],  1'b0};
                readAddr13  = {readAddr[12:0],  1'b0};
                readAddr12  = {readAddr[12:0],  1'b0};
                readAddr11  = {readAddr[12:0],  1'b0};
                readAddr10  = {readAddr[11:0],  2'b0};
                readAddr9  = {readAddr[11:0],  2'b0};
                readAddr8  = {readAddr[11:0],  2'b0};
                readAddr7  = {readAddr[11:0],  2'b0};
                readAddr6  = {readAddr[11:0],  2'b0};
                readAddr5  = {readAddr[11:0],  2'b0};
                readAddr4  = {readAddr[11:0],  2'b0};
                readAddr3  = {readAddr[11:0],  2'b0};
                readAddr2  = {readAddr[9:0],  4'b0};
                readAddr1  = {readAddr[9:0],  4'b0};

                writeData58 = {17'b0, writeData[31]};
                writeData57 = {17'b0, writeData[30]};
                writeData56 = {17'b0, writeData[29]};
                writeData55 = {17'b0, writeData[28]};
                writeData54 = {17'b0, writeData[27]};
                writeData53 = {17'b0, writeData[26]};
                writeData52 = {17'b0, writeData[25]};
                writeData51 = {17'b0, writeData[24]};
                writeData50 = {17'b0, writeData[23]};
                writeData49 = {17'b0, writeData[22]};
                writeData48 = {17'b0, writeData[21]};
                writeData47 = {17'b0, writeData[20]};
                writeData46 = {17'b0, writeData[19]};
                writeData45 = {17'b0, writeData[18]};
                writeData44 = {17'b0, writeData[17]};
                writeData43 = {17'b0, writeData[16]};
                writeData42 = {17'b0, writeData[15]};
                writeData41 = {17'b0, writeData[14]};
                writeData40 = {17'b0, writeData[13]};
                writeData39 = {17'b0, writeData[12]};
                writeData38 = {17'b0, writeData[11]};
                writeData37 = {17'b0, writeData[10]};
                writeData36 = {17'b0, writeData[9]};
                writeData35 = {17'b0, writeData[8]};
                writeData34 = {17'b0, writeData[7]};
                writeData33 = {17'b0, writeData[6]};
                writeData32 = {17'b0, writeData[5]};
                writeData31 = {17'b0, writeData[4]};
                writeData30 = {17'b0, writeData[3]};
                writeData29 = {17'b0, writeData[2]};
                writeData28 = {17'b0, writeData[1]};
                writeData27 = {17'b0, writeData[0]};
                writeData26 = {16'b0, writeData[31:30]};
                writeData25 = {16'b0, writeData[29:28]};
                writeData24 = {16'b0, writeData[27:26]};
                writeData23 = {16'b0, writeData[25:24]};
                writeData22 = {16'b0, writeData[23:22]};
                writeData21 = {16'b0, writeData[21:20]};
                writeData20 = {16'b0, writeData[19:18]};
                writeData19 = {16'b0, writeData[17:16]};
                writeData18 = {16'b0, writeData[15:14]};
                writeData17 = {16'b0, writeData[13:12]};
                writeData16 = {16'b0, writeData[11:10]};
                writeData15 = {16'b0, writeData[9:8]};
                writeData14 = {16'b0, writeData[7:6]};
                writeData13 = {16'b0, writeData[5:4]};
                writeData12 = {16'b0, writeData[3:2]};
                writeData11 = {16'b0, writeData[1:0]};
                writeData10 = {14'b0, writeData[31:28]};
                writeData9 = {14'b0, writeData[27:24]};
                writeData8 = {14'b0, writeData[23:20]};
                writeData7 = {14'b0, writeData[19:16]};
                writeData6 = {14'b0, writeData[15:12]};
                writeData5 = {14'b0, writeData[11:8]};
                writeData4 = {14'b0, writeData[7:4]};
                writeData3 = {14'b0, writeData[3:0]};
                writeData2 = {1'b0, writeData[31:24], 1'b0, writeData[23:16]};
                writeData1 = {1'b0, writeData[15:8], 1'b0, writeData[7:0]};

                case (writeAddr[14:9])
                    6'b000000, 6'b000001, 6'b000010, 6'b000011,
                    6'b000100, 6'b000101, 6'b000110, 6'b000111,
                    6'b001000, 6'b001001, 6'b001010, 6'b001011,
                    6'b001100, 6'b001101, 6'b001110, 6'b001111,
                    6'b010000, 6'b010001, 6'b010010, 6'b010011,
                    6'b010100, 6'b010101, 6'b010110, 6'b010111,
                    6'b011000, 6'b011001, 6'b011010, 6'b011011,
                    6'b011100, 6'b011101, 6'b011110, 6'b011111 : begin
                        wen_a58 = {1'b0, wen};
                        wen_a57 = {1'b0, wen};
                        wen_a56 = {1'b0, wen};
                        wen_a55 = {1'b0, wen};
                        wen_a54 = {1'b0, wen};
                        wen_a53 = {1'b0, wen};
                        wen_a52 = {1'b0, wen};
                        wen_a51 = {1'b0, wen};
                        wen_a50 = {1'b0, wen};
                        wen_a49 = {1'b0, wen};
                        wen_a48 = {1'b0, wen};
                        wen_a47 = {1'b0, wen};
                        wen_a46 = {1'b0, wen};
                        wen_a45 = {1'b0, wen};
                        wen_a44 = {1'b0, wen};
                        wen_a43 = {1'b0, wen};
                        wen_a42 = {1'b0, wen};
                        wen_a41 = {1'b0, wen};
                        wen_a40 = {1'b0, wen};
                        wen_a39 = {1'b0, wen};
                        wen_a38 = {1'b0, wen};
                        wen_a37 = {1'b0, wen};
                        wen_a36 = {1'b0, wen};
                        wen_a35 = {1'b0, wen};
                        wen_a34 = {1'b0, wen};
                        wen_a33 = {1'b0, wen};
                        wen_a32 = {1'b0, wen};
                        wen_a31 = {1'b0, wen};
                        wen_a30 = {1'b0, wen};
                        wen_a29 = {1'b0, wen};
                        wen_a28 = {1'b0, wen};
                        wen_a27 = {1'b0, wen};
                        wen_a26 = {1'b0, 1'b0};
                        wen_a25 = {1'b0, 1'b0};
                        wen_a24 = {1'b0, 1'b0};
                        wen_a23 = {1'b0, 1'b0};
                        wen_a22 = {1'b0, 1'b0};
                        wen_a21 = {1'b0, 1'b0};
                        wen_a20 = {1'b0, 1'b0};
                        wen_a19 = {1'b0, 1'b0};
                        wen_a18 = {1'b0, 1'b0};
                        wen_a17 = {1'b0, 1'b0};
                        wen_a16 = {1'b0, 1'b0};
                        wen_a15 = {1'b0, 1'b0};
                        wen_a14 = {1'b0, 1'b0};
                        wen_a13 = {1'b0, 1'b0};
                        wen_a12 = {1'b0, 1'b0};
                        wen_a11 = {1'b0, 1'b0};
                        wen_a10 = {1'b0, 1'b0};
                        wen_a9 = {1'b0, 1'b0};
                        wen_a8 = {1'b0, 1'b0};
                        wen_a7 = {1'b0, 1'b0};
                        wen_a6 = {1'b0, 1'b0};
                        wen_a5 = {1'b0, 1'b0};
                        wen_a4 = {1'b0, 1'b0};
                        wen_a3 = {1'b0, 1'b0};
                        wen_a2 = {1'b0, 1'b0};
                        wen_a1 = {1'b0, 1'b0};
                    end
                    6'b100000, 6'b100001, 6'b100010, 6'b100011,
                    6'b100100, 6'b100101, 6'b100110, 6'b100111,
                    6'b101000, 6'b101001, 6'b101010, 6'b101011,
                    6'b101100, 6'b101101, 6'b101110, 6'b101111 : begin
                        wen_a58 = {1'b0, 1'b0};
                        wen_a57 = {1'b0, 1'b0};
                        wen_a56 = {1'b0, 1'b0};
                        wen_a55 = {1'b0, 1'b0};
                        wen_a54 = {1'b0, 1'b0};
                        wen_a53 = {1'b0, 1'b0};
                        wen_a52 = {1'b0, 1'b0};
                        wen_a51 = {1'b0, 1'b0};
                        wen_a50 = {1'b0, 1'b0};
                        wen_a49 = {1'b0, 1'b0};
                        wen_a48 = {1'b0, 1'b0};
                        wen_a47 = {1'b0, 1'b0};
                        wen_a46 = {1'b0, 1'b0};
                        wen_a45 = {1'b0, 1'b0};
                        wen_a44 = {1'b0, 1'b0};
                        wen_a43 = {1'b0, 1'b0};
                        wen_a42 = {1'b0, 1'b0};
                        wen_a41 = {1'b0, 1'b0};
                        wen_a40 = {1'b0, 1'b0};
                        wen_a39 = {1'b0, 1'b0};
                        wen_a38 = {1'b0, 1'b0};
                        wen_a37 = {1'b0, 1'b0};
                        wen_a36 = {1'b0, 1'b0};
                        wen_a35 = {1'b0, 1'b0};
                        wen_a34 = {1'b0, 1'b0};
                        wen_a33 = {1'b0, 1'b0};
                        wen_a32 = {1'b0, 1'b0};
                        wen_a31 = {1'b0, 1'b0};
                        wen_a30 = {1'b0, 1'b0};
                        wen_a29 = {1'b0, 1'b0};
                        wen_a28 = {1'b0, 1'b0};
                        wen_a27 = {1'b0, 1'b0};
                        wen_a26 = {1'b0, wen};
                        wen_a25 = {1'b0, wen};
                        wen_a24 = {1'b0, wen};
                        wen_a23 = {1'b0, wen};
                        wen_a22 = {1'b0, wen};
                        wen_a21 = {1'b0, wen};
                        wen_a20 = {1'b0, wen};
                        wen_a19 = {1'b0, wen};
                        wen_a18 = {1'b0, wen};
                        wen_a17 = {1'b0, wen};
                        wen_a16 = {1'b0, wen};
                        wen_a15 = {1'b0, wen};
                        wen_a14 = {1'b0, wen};
                        wen_a13 = {1'b0, wen};
                        wen_a12 = {1'b0, wen};
                        wen_a11 = {1'b0, wen};
                        wen_a10 = {1'b0, 1'b0};
                        wen_a9 = {1'b0, 1'b0};
                        wen_a8 = {1'b0, 1'b0};
                        wen_a7 = {1'b0, 1'b0};
                        wen_a6 = {1'b0, 1'b0};
                        wen_a5 = {1'b0, 1'b0};
                        wen_a4 = {1'b0, 1'b0};
                        wen_a3 = {1'b0, 1'b0};
                        wen_a2 = {1'b0, 1'b0};
                        wen_a1 = {1'b0, 1'b0};
                    end
                    6'b110000, 6'b110001, 6'b110010, 6'b110011,
                    6'b110100, 6'b110101, 6'b110110, 6'b110111 : begin
                        wen_a58 = {1'b0, 1'b0};
                        wen_a57 = {1'b0, 1'b0};
                        wen_a56 = {1'b0, 1'b0};
                        wen_a55 = {1'b0, 1'b0};
                        wen_a54 = {1'b0, 1'b0};
                        wen_a53 = {1'b0, 1'b0};
                        wen_a52 = {1'b0, 1'b0};
                        wen_a51 = {1'b0, 1'b0};
                        wen_a50 = {1'b0, 1'b0};
                        wen_a49 = {1'b0, 1'b0};
                        wen_a48 = {1'b0, 1'b0};
                        wen_a47 = {1'b0, 1'b0};
                        wen_a46 = {1'b0, 1'b0};
                        wen_a45 = {1'b0, 1'b0};
                        wen_a44 = {1'b0, 1'b0};
                        wen_a43 = {1'b0, 1'b0};
                        wen_a42 = {1'b0, 1'b0};
                        wen_a41 = {1'b0, 1'b0};
                        wen_a40 = {1'b0, 1'b0};
                        wen_a39 = {1'b0, 1'b0};
                        wen_a38 = {1'b0, 1'b0};
                        wen_a37 = {1'b0, 1'b0};
                        wen_a36 = {1'b0, 1'b0};
                        wen_a35 = {1'b0, 1'b0};
                        wen_a34 = {1'b0, 1'b0};
                        wen_a33 = {1'b0, 1'b0};
                        wen_a32 = {1'b0, 1'b0};
                        wen_a31 = {1'b0, 1'b0};
                        wen_a30 = {1'b0, 1'b0};
                        wen_a29 = {1'b0, 1'b0};
                        wen_a28 = {1'b0, 1'b0};
                        wen_a27 = {1'b0, 1'b0};
                        wen_a26 = {1'b0, 1'b0};
                        wen_a25 = {1'b0, 1'b0};
                        wen_a24 = {1'b0, 1'b0};
                        wen_a23 = {1'b0, 1'b0};
                        wen_a22 = {1'b0, 1'b0};
                        wen_a21 = {1'b0, 1'b0};
                        wen_a20 = {1'b0, 1'b0};
                        wen_a19 = {1'b0, 1'b0};
                        wen_a18 = {1'b0, 1'b0};
                        wen_a17 = {1'b0, 1'b0};
                        wen_a16 = {1'b0, 1'b0};
                        wen_a15 = {1'b0, 1'b0};
                        wen_a14 = {1'b0, 1'b0};
                        wen_a13 = {1'b0, 1'b0};
                        wen_a12 = {1'b0, 1'b0};
                        wen_a11 = {1'b0, 1'b0};
                        wen_a10 = {1'b0, wen};
                        wen_a9 = {1'b0, wen};
                        wen_a8 = {1'b0, wen};
                        wen_a7 = {1'b0, wen};
                        wen_a6 = {1'b0, wen};
                        wen_a5 = {1'b0, wen};
                        wen_a4 = {1'b0, wen};
                        wen_a3 = {1'b0, wen};
                        wen_a2 = {1'b0, 1'b0};
                        wen_a1 = {1'b0, 1'b0};
                    end
                    6'b111000, 6'b111001 : begin
                        wen_a58 = {1'b0, 1'b0};
                        wen_a57 = {1'b0, 1'b0};
                        wen_a56 = {1'b0, 1'b0};
                        wen_a55 = {1'b0, 1'b0};
                        wen_a54 = {1'b0, 1'b0};
                        wen_a53 = {1'b0, 1'b0};
                        wen_a52 = {1'b0, 1'b0};
                        wen_a51 = {1'b0, 1'b0};
                        wen_a50 = {1'b0, 1'b0};
                        wen_a49 = {1'b0, 1'b0};
                        wen_a48 = {1'b0, 1'b0};
                        wen_a47 = {1'b0, 1'b0};
                        wen_a46 = {1'b0, 1'b0};
                        wen_a45 = {1'b0, 1'b0};
                        wen_a44 = {1'b0, 1'b0};
                        wen_a43 = {1'b0, 1'b0};
                        wen_a42 = {1'b0, 1'b0};
                        wen_a41 = {1'b0, 1'b0};
                        wen_a40 = {1'b0, 1'b0};
                        wen_a39 = {1'b0, 1'b0};
                        wen_a38 = {1'b0, 1'b0};
                        wen_a37 = {1'b0, 1'b0};
                        wen_a36 = {1'b0, 1'b0};
                        wen_a35 = {1'b0, 1'b0};
                        wen_a34 = {1'b0, 1'b0};
                        wen_a33 = {1'b0, 1'b0};
                        wen_a32 = {1'b0, 1'b0};
                        wen_a31 = {1'b0, 1'b0};
                        wen_a30 = {1'b0, 1'b0};
                        wen_a29 = {1'b0, 1'b0};
                        wen_a28 = {1'b0, 1'b0};
                        wen_a27 = {1'b0, 1'b0};
                        wen_a26 = {1'b0, 1'b0};
                        wen_a25 = {1'b0, 1'b0};
                        wen_a24 = {1'b0, 1'b0};
                        wen_a23 = {1'b0, 1'b0};
                        wen_a22 = {1'b0, 1'b0};
                        wen_a21 = {1'b0, 1'b0};
                        wen_a20 = {1'b0, 1'b0};
                        wen_a19 = {1'b0, 1'b0};
                        wen_a18 = {1'b0, 1'b0};
                        wen_a17 = {1'b0, 1'b0};
                        wen_a16 = {1'b0, 1'b0};
                        wen_a15 = {1'b0, 1'b0};
                        wen_a14 = {1'b0, 1'b0};
                        wen_a13 = {1'b0, 1'b0};
                        wen_a12 = {1'b0, 1'b0};
                        wen_a11 = {1'b0, 1'b0};
                        wen_a10 = {1'b0, 1'b0};
                        wen_a9 = {1'b0, 1'b0};
                        wen_a8 = {1'b0, 1'b0};
                        wen_a7 = {1'b0, 1'b0};
                        wen_a6 = {1'b0, 1'b0};
                        wen_a5 = {1'b0, 1'b0};
                        wen_a4 = {1'b0, 1'b0};
                        wen_a3 = {1'b0, 1'b0};
                        wen_a2 = {wen, wen};
                        wen_a1 = {wen, wen};
                    end
                    default : begin
                        wen_a58 = {1'b0, 1'b0};
                        wen_a57 = {1'b0, 1'b0};
                        wen_a56 = {1'b0, 1'b0};
                        wen_a55 = {1'b0, 1'b0};
                        wen_a54 = {1'b0, 1'b0};
                        wen_a53 = {1'b0, 1'b0};
                        wen_a52 = {1'b0, 1'b0};
                        wen_a51 = {1'b0, 1'b0};
                        wen_a50 = {1'b0, 1'b0};
                        wen_a49 = {1'b0, 1'b0};
                        wen_a48 = {1'b0, 1'b0};
                        wen_a47 = {1'b0, 1'b0};
                        wen_a46 = {1'b0, 1'b0};
                        wen_a45 = {1'b0, 1'b0};
                        wen_a44 = {1'b0, 1'b0};
                        wen_a43 = {1'b0, 1'b0};
                        wen_a42 = {1'b0, 1'b0};
                        wen_a41 = {1'b0, 1'b0};
                        wen_a40 = {1'b0, 1'b0};
                        wen_a39 = {1'b0, 1'b0};
                        wen_a38 = {1'b0, 1'b0};
                        wen_a37 = {1'b0, 1'b0};
                        wen_a36 = {1'b0, 1'b0};
                        wen_a35 = {1'b0, 1'b0};
                        wen_a34 = {1'b0, 1'b0};
                        wen_a33 = {1'b0, 1'b0};
                        wen_a32 = {1'b0, 1'b0};
                        wen_a31 = {1'b0, 1'b0};
                        wen_a30 = {1'b0, 1'b0};
                        wen_a29 = {1'b0, 1'b0};
                        wen_a28 = {1'b0, 1'b0};
                        wen_a27 = {1'b0, 1'b0};
                        wen_a26 = {1'b0, 1'b0};
                        wen_a25 = {1'b0, 1'b0};
                        wen_a24 = {1'b0, 1'b0};
                        wen_a23 = {1'b0, 1'b0};
                        wen_a22 = {1'b0, 1'b0};
                        wen_a21 = {1'b0, 1'b0};
                        wen_a20 = {1'b0, 1'b0};
                        wen_a19 = {1'b0, 1'b0};
                        wen_a18 = {1'b0, 1'b0};
                        wen_a17 = {1'b0, 1'b0};
                        wen_a16 = {1'b0, 1'b0};
                        wen_a15 = {1'b0, 1'b0};
                        wen_a14 = {1'b0, 1'b0};
                        wen_a13 = {1'b0, 1'b0};
                        wen_a12 = {1'b0, 1'b0};
                        wen_a11 = {1'b0, 1'b0};
                        wen_a10 = {1'b0, 1'b0};
                        wen_a9 = {1'b0, 1'b0};
                        wen_a8 = {1'b0, 1'b0};
                        wen_a7 = {1'b0, 1'b0};
                        wen_a6 = {1'b0, 1'b0};
                        wen_a5 = {1'b0, 1'b0};
                        wen_a4 = {1'b0, 1'b0};
                        wen_a3 = {1'b0, 1'b0};
                        wen_a2 = {1'b0, 1'b0};
                        wen_a1 = {1'b0, 1'b0};
                    end
                endcase

                case (ckRdAddr[14:9])
                    6'b000000, 6'b000001, 6'b000010, 6'b000011,
                    6'b000100, 6'b000101, 6'b000110, 6'b000111,
                    6'b001000, 6'b001001, 6'b001010, 6'b001011,
                    6'b001100, 6'b001101, 6'b001110, 6'b001111,
                    6'b010000, 6'b010001, 6'b010010, 6'b010011,
                    6'b010100, 6'b010101, 6'b010110, 6'b010111,
                    6'b011000, 6'b011001, 6'b011010, 6'b011011,
                    6'b011100, 6'b011101, 6'b011110, 6'b011111 : begin
                        readData = {
                                        readData58[0],
                                        readData57[0],
                                        readData56[0],
                                        readData55[0],
                                        readData54[0],
                                        readData53[0],
                                        readData52[0],
                                        readData51[0],
                                        readData50[0],
                                        readData49[0],
                                        readData48[0],
                                        readData47[0],
                                        readData46[0],
                                        readData45[0],
                                        readData44[0],
                                        readData43[0],
                                        readData42[0],
                                        readData41[0],
                                        readData40[0],
                                        readData39[0],
                                        readData38[0],
                                        readData37[0],
                                        readData36[0],
                                        readData35[0],
                                        readData34[0],
                                        readData33[0],
                                        readData32[0],
                                        readData31[0],
                                        readData30[0],
                                        readData29[0],
                                        readData28[0],
                                        readData27[0]
                        };
                    end
                    6'b100000, 6'b100001, 6'b100010, 6'b100011,
                    6'b100100, 6'b100101, 6'b100110, 6'b100111,
                    6'b101000, 6'b101001, 6'b101010, 6'b101011,
                    6'b101100, 6'b101101, 6'b101110, 6'b101111 : begin
                        readData = {
                                        readData26[1:0],
                                        readData25[1:0],
                                        readData24[1:0],
                                        readData23[1:0],
                                        readData22[1:0],
                                        readData21[1:0],
                                        readData20[1:0],
                                        readData19[1:0],
                                        readData18[1:0],
                                        readData17[1:0],
                                        readData16[1:0],
                                        readData15[1:0],
                                        readData14[1:0],
                                        readData13[1:0],
                                        readData12[1:0],
                                        readData11[1:0]
                        };
                    end
                    6'b110000, 6'b110001, 6'b110010, 6'b110011,
                    6'b110100, 6'b110101, 6'b110110, 6'b110111 : begin
                        readData = {
                                        readData10[3:0],
                                        readData9[3:0],
                                        readData8[3:0],
                                        readData7[3:0],
                                        readData6[3:0],
                                        readData5[3:0],
                                        readData4[3:0],
                                        readData3[3:0]
                        };
                    end
                    6'b111000, 6'b111001 : begin
                        readData = {readData2[16:9],readData2[7:0],readData1[16:9],readData1[7:0]};
                    end
                    default : begin
                        readData = 32'b0;
                    end
                endcase
            end        
            30208: begin
                width58 = 3'b000;
                width57 = 3'b000;
                width56 = 3'b000;
                width55 = 3'b000;
                width54 = 3'b000;
                width53 = 3'b000;
                width52 = 3'b000;
                width51 = 3'b000;
                width50 = 3'b000;
                width49 = 3'b000;
                width48 = 3'b000;
                width47 = 3'b000;
                width46 = 3'b000;
                width45 = 3'b000;
                width44 = 3'b000;
                width43 = 3'b000;
                width42 = 3'b000;
                width41 = 3'b000;
                width40 = 3'b000;
                width39 = 3'b000;
                width38 = 3'b000;
                width37 = 3'b000;
                width36 = 3'b000;
                width35 = 3'b000;
                width34 = 3'b000;
                width33 = 3'b000;
                width32 = 3'b000;
                width31 = 3'b000;
                width30 = 3'b000;
                width29 = 3'b000;
                width28 = 3'b000;
                width27 = 3'b000;
                width26 = 3'b001;
                width25 = 3'b001;
                width24 = 3'b001;
                width23 = 3'b001;
                width22 = 3'b001;
                width21 = 3'b001;
                width20 = 3'b001;
                width19 = 3'b001;
                width18 = 3'b001;
                width17 = 3'b001;
                width16 = 3'b001;
                width15 = 3'b001;
                width14 = 3'b001;
                width13 = 3'b001;
                width12 = 3'b001;
                width11 = 3'b001;
                width10 = 3'b010;
                width9 = 3'b010;
                width8 = 3'b010;
                width7 = 3'b010;
                width6 = 3'b010;
                width5 = 3'b010;
                width4 = 3'b010;
                width3 = 3'b010;
                width2 = 3'b100;
                width1 = 3'b100;
                width0 = 3'b101;

                writeAddr58 = {writeAddr[13:0]};
                writeAddr57 = {writeAddr[13:0]};
                writeAddr56 = {writeAddr[13:0]};
                writeAddr55 = {writeAddr[13:0]};
                writeAddr54 = {writeAddr[13:0]};
                writeAddr53 = {writeAddr[13:0]};
                writeAddr52 = {writeAddr[13:0]};
                writeAddr51 = {writeAddr[13:0]};
                writeAddr50 = {writeAddr[13:0]};
                writeAddr49 = {writeAddr[13:0]};
                writeAddr48 = {writeAddr[13:0]};
                writeAddr47 = {writeAddr[13:0]};
                writeAddr46 = {writeAddr[13:0]};
                writeAddr45 = {writeAddr[13:0]};
                writeAddr44 = {writeAddr[13:0]};
                writeAddr43 = {writeAddr[13:0]};
                writeAddr42 = {writeAddr[13:0]};
                writeAddr41 = {writeAddr[13:0]};
                writeAddr40 = {writeAddr[13:0]};
                writeAddr39 = {writeAddr[13:0]};
                writeAddr38 = {writeAddr[13:0]};
                writeAddr37 = {writeAddr[13:0]};
                writeAddr36 = {writeAddr[13:0]};
                writeAddr35 = {writeAddr[13:0]};
                writeAddr34 = {writeAddr[13:0]};
                writeAddr33 = {writeAddr[13:0]};
                writeAddr32 = {writeAddr[13:0]};
                writeAddr31 = {writeAddr[13:0]};
                writeAddr30 = {writeAddr[13:0]};
                writeAddr29 = {writeAddr[13:0]};
                writeAddr28 = {writeAddr[13:0]};
                writeAddr27 = {writeAddr[13:0]};
                writeAddr26 = {writeAddr[12:0], 1'b0};
                writeAddr25 = {writeAddr[12:0], 1'b0};
                writeAddr24 = {writeAddr[12:0], 1'b0};
                writeAddr23 = {writeAddr[12:0], 1'b0};
                writeAddr22 = {writeAddr[12:0], 1'b0};
                writeAddr21 = {writeAddr[12:0], 1'b0};
                writeAddr20 = {writeAddr[12:0], 1'b0};
                writeAddr19 = {writeAddr[12:0], 1'b0};
                writeAddr18 = {writeAddr[12:0], 1'b0};
                writeAddr17 = {writeAddr[12:0], 1'b0};
                writeAddr16 = {writeAddr[12:0], 1'b0};
                writeAddr15 = {writeAddr[12:0], 1'b0};
                writeAddr14 = {writeAddr[12:0], 1'b0};
                writeAddr13 = {writeAddr[12:0], 1'b0};
                writeAddr12 = {writeAddr[12:0], 1'b0};
                writeAddr11 = {writeAddr[12:0], 1'b0};
                writeAddr10 = {writeAddr[11:0], 2'b0};
                writeAddr9 = {writeAddr[11:0], 2'b0};
                writeAddr8 = {writeAddr[11:0], 2'b0};
                writeAddr7 = {writeAddr[11:0], 2'b0};
                writeAddr6 = {writeAddr[11:0], 2'b0};
                writeAddr5 = {writeAddr[11:0], 2'b0};
                writeAddr4 = {writeAddr[11:0], 2'b0};
                writeAddr3 = {writeAddr[11:0], 2'b0};
                writeAddr2 = {writeAddr[9:0], 4'b0};
                writeAddr1 = {writeAddr[9:0], 4'b0};
                writeAddr0 = {writeAddr[8:0], 5'b0};

                readAddr58 = {writeAddr[13:0]};
                readAddr57 = {writeAddr[13:0]};
                readAddr56 = {writeAddr[13:0]};
                readAddr55 = {writeAddr[13:0]};
                readAddr54 = {writeAddr[13:0]};
                readAddr53 = {writeAddr[13:0]};
                readAddr52 = {writeAddr[13:0]};
                readAddr51 = {writeAddr[13:0]};
                readAddr50 = {writeAddr[13:0]};
                readAddr49 = {writeAddr[13:0]};
                readAddr48 = {writeAddr[13:0]};
                readAddr47 = {writeAddr[13:0]};
                readAddr46 = {writeAddr[13:0]};
                readAddr45 = {writeAddr[13:0]};
                readAddr44 = {writeAddr[13:0]};
                readAddr43 = {writeAddr[13:0]};
                readAddr42 = {writeAddr[13:0]};
                readAddr41 = {writeAddr[13:0]};
                readAddr40 = {writeAddr[13:0]};
                readAddr39 = {writeAddr[13:0]};
                readAddr38 = {writeAddr[13:0]};
                readAddr37 = {writeAddr[13:0]};
                readAddr36 = {writeAddr[13:0]};
                readAddr35 = {writeAddr[13:0]};
                readAddr34 = {writeAddr[13:0]};
                readAddr33 = {writeAddr[13:0]};
                readAddr32 = {writeAddr[13:0]};
                readAddr31 = {writeAddr[13:0]};
                readAddr30 = {writeAddr[13:0]};
                readAddr29 = {writeAddr[13:0]};
                readAddr28 = {writeAddr[13:0]};
                readAddr27 = {writeAddr[13:0]};
                readAddr26  = {readAddr[12:0],  1'b0};
                readAddr25  = {readAddr[12:0],  1'b0};
                readAddr24  = {readAddr[12:0],  1'b0};
                readAddr23  = {readAddr[12:0],  1'b0};
                readAddr22  = {readAddr[12:0],  1'b0};
                readAddr21  = {readAddr[12:0],  1'b0};
                readAddr20  = {readAddr[12:0],  1'b0};
                readAddr19  = {readAddr[12:0],  1'b0};
                readAddr18  = {readAddr[12:0],  1'b0};
                readAddr17  = {readAddr[12:0],  1'b0};
                readAddr16  = {readAddr[12:0],  1'b0};
                readAddr15  = {readAddr[12:0],  1'b0};
                readAddr14  = {readAddr[12:0],  1'b0};
                readAddr13  = {readAddr[12:0],  1'b0};
                readAddr12  = {readAddr[12:0],  1'b0};
                readAddr11  = {readAddr[12:0],  1'b0};
                readAddr10  = {readAddr[11:0],  2'b0};
                readAddr9  = {readAddr[11:0],  2'b0};
                readAddr8  = {readAddr[11:0],  2'b0};
                readAddr7  = {readAddr[11:0],  2'b0};
                readAddr6  = {readAddr[11:0],  2'b0};
                readAddr5  = {readAddr[11:0],  2'b0};
                readAddr4  = {readAddr[11:0],  2'b0};
                readAddr3  = {readAddr[11:0],  2'b0};
                readAddr2  = {readAddr[9:0],  4'b0};
                readAddr1  = {readAddr[9:0],  4'b0};
                readAddr0  = {readAddr[8:0],  5'b0};

                writeData58 = {17'b0, writeData[31]};
                writeData57 = {17'b0, writeData[30]};
                writeData56 = {17'b0, writeData[29]};
                writeData55 = {17'b0, writeData[28]};
                writeData54 = {17'b0, writeData[27]};
                writeData53 = {17'b0, writeData[26]};
                writeData52 = {17'b0, writeData[25]};
                writeData51 = {17'b0, writeData[24]};
                writeData50 = {17'b0, writeData[23]};
                writeData49 = {17'b0, writeData[22]};
                writeData48 = {17'b0, writeData[21]};
                writeData47 = {17'b0, writeData[20]};
                writeData46 = {17'b0, writeData[19]};
                writeData45 = {17'b0, writeData[18]};
                writeData44 = {17'b0, writeData[17]};
                writeData43 = {17'b0, writeData[16]};
                writeData42 = {17'b0, writeData[15]};
                writeData41 = {17'b0, writeData[14]};
                writeData40 = {17'b0, writeData[13]};
                writeData39 = {17'b0, writeData[12]};
                writeData38 = {17'b0, writeData[11]};
                writeData37 = {17'b0, writeData[10]};
                writeData36 = {17'b0, writeData[9]};
                writeData35 = {17'b0, writeData[8]};
                writeData34 = {17'b0, writeData[7]};
                writeData33 = {17'b0, writeData[6]};
                writeData32 = {17'b0, writeData[5]};
                writeData31 = {17'b0, writeData[4]};
                writeData30 = {17'b0, writeData[3]};
                writeData29 = {17'b0, writeData[2]};
                writeData28 = {17'b0, writeData[1]};
                writeData27 = {17'b0, writeData[0]};
                writeData26 = {16'b0, writeData[31:30]};
                writeData25 = {16'b0, writeData[29:28]};
                writeData24 = {16'b0, writeData[27:26]};
                writeData23 = {16'b0, writeData[25:24]};
                writeData22 = {16'b0, writeData[23:22]};
                writeData21 = {16'b0, writeData[21:20]};
                writeData20 = {16'b0, writeData[19:18]};
                writeData19 = {16'b0, writeData[17:16]};
                writeData18 = {16'b0, writeData[15:14]};
                writeData17 = {16'b0, writeData[13:12]};
                writeData16 = {16'b0, writeData[11:10]};
                writeData15 = {16'b0, writeData[9:8]};
                writeData14 = {16'b0, writeData[7:6]};
                writeData13 = {16'b0, writeData[5:4]};
                writeData12 = {16'b0, writeData[3:2]};
                writeData11 = {16'b0, writeData[1:0]};
                writeData10 = {14'b0, writeData[31:28]};
                writeData9 = {14'b0, writeData[27:24]};
                writeData8 = {14'b0, writeData[23:20]};
                writeData7 = {14'b0, writeData[19:16]};
                writeData6 = {14'b0, writeData[15:12]};
                writeData5 = {14'b0, writeData[11:8]};
                writeData4 = {14'b0, writeData[7:4]};
                writeData3 = {14'b0, writeData[3:0]};
                writeData2 = {1'b0, writeData[31:24], 1'b0, writeData[23:16]};
                writeData1 = {1'b0, writeData[15:8], 1'b0, writeData[7:0]};
                writeData0 = {1'b0, writeData[31:24], 1'b0, writeData[23:16], 1'b0, writeData[15:8], 1'b0, writeData[7:0]};

                case (writeAddr[14:9])
                    6'b000000, 6'b000001, 6'b000010, 6'b000011,
                    6'b000100, 6'b000101, 6'b000110, 6'b000111,
                    6'b001000, 6'b001001, 6'b001010, 6'b001011,
                    6'b001100, 6'b001101, 6'b001110, 6'b001111,
                    6'b010000, 6'b010001, 6'b010010, 6'b010011,
                    6'b010100, 6'b010101, 6'b010110, 6'b010111,
                    6'b011000, 6'b011001, 6'b011010, 6'b011011,
                    6'b011100, 6'b011101, 6'b011110, 6'b011111 : begin
                        wen_a58 = {1'b0, wen};
                        wen_a57 = {1'b0, wen};
                        wen_a56 = {1'b0, wen};
                        wen_a55 = {1'b0, wen};
                        wen_a54 = {1'b0, wen};
                        wen_a53 = {1'b0, wen};
                        wen_a52 = {1'b0, wen};
                        wen_a51 = {1'b0, wen};
                        wen_a50 = {1'b0, wen};
                        wen_a49 = {1'b0, wen};
                        wen_a48 = {1'b0, wen};
                        wen_a47 = {1'b0, wen};
                        wen_a46 = {1'b0, wen};
                        wen_a45 = {1'b0, wen};
                        wen_a44 = {1'b0, wen};
                        wen_a43 = {1'b0, wen};
                        wen_a42 = {1'b0, wen};
                        wen_a41 = {1'b0, wen};
                        wen_a40 = {1'b0, wen};
                        wen_a39 = {1'b0, wen};
                        wen_a38 = {1'b0, wen};
                        wen_a37 = {1'b0, wen};
                        wen_a36 = {1'b0, wen};
                        wen_a35 = {1'b0, wen};
                        wen_a34 = {1'b0, wen};
                        wen_a33 = {1'b0, wen};
                        wen_a32 = {1'b0, wen};
                        wen_a31 = {1'b0, wen};
                        wen_a30 = {1'b0, wen};
                        wen_a29 = {1'b0, wen};
                        wen_a28 = {1'b0, wen};
                        wen_a27 = {1'b0, wen};
                        wen_a26 = {1'b0, 1'b0};
                        wen_a25 = {1'b0, 1'b0};
                        wen_a24 = {1'b0, 1'b0};
                        wen_a23 = {1'b0, 1'b0};
                        wen_a22 = {1'b0, 1'b0};
                        wen_a21 = {1'b0, 1'b0};
                        wen_a20 = {1'b0, 1'b0};
                        wen_a19 = {1'b0, 1'b0};
                        wen_a18 = {1'b0, 1'b0};
                        wen_a17 = {1'b0, 1'b0};
                        wen_a16 = {1'b0, 1'b0};
                        wen_a15 = {1'b0, 1'b0};
                        wen_a14 = {1'b0, 1'b0};
                        wen_a13 = {1'b0, 1'b0};
                        wen_a12 = {1'b0, 1'b0};
                        wen_a11 = {1'b0, 1'b0};
                        wen_a10 = {1'b0, 1'b0};
                        wen_a9 = {1'b0, 1'b0};
                        wen_a8 = {1'b0, 1'b0};
                        wen_a7 = {1'b0, 1'b0};
                        wen_a6 = {1'b0, 1'b0};
                        wen_a5 = {1'b0, 1'b0};
                        wen_a4 = {1'b0, 1'b0};
                        wen_a3 = {1'b0, 1'b0};
                        wen_a2 = {1'b0, 1'b0};
                        wen_a1 = {1'b0, 1'b0};
                        wen_a0 = {1'b0, 1'b0};
                        wen_b0 = {1'b0, 1'b0};
                    end
                    6'b100000, 6'b100001, 6'b100010, 6'b100011,
                    6'b100100, 6'b100101, 6'b100110, 6'b100111,
                    6'b101000, 6'b101001, 6'b101010, 6'b101011,
                    6'b101100, 6'b101101, 6'b101110, 6'b101111 : begin
                        wen_a58 = {1'b0, 1'b0};
                        wen_a57 = {1'b0, 1'b0};
                        wen_a56 = {1'b0, 1'b0};
                        wen_a55 = {1'b0, 1'b0};
                        wen_a54 = {1'b0, 1'b0};
                        wen_a53 = {1'b0, 1'b0};
                        wen_a52 = {1'b0, 1'b0};
                        wen_a51 = {1'b0, 1'b0};
                        wen_a50 = {1'b0, 1'b0};
                        wen_a49 = {1'b0, 1'b0};
                        wen_a48 = {1'b0, 1'b0};
                        wen_a47 = {1'b0, 1'b0};
                        wen_a46 = {1'b0, 1'b0};
                        wen_a45 = {1'b0, 1'b0};
                        wen_a44 = {1'b0, 1'b0};
                        wen_a43 = {1'b0, 1'b0};
                        wen_a42 = {1'b0, 1'b0};
                        wen_a41 = {1'b0, 1'b0};
                        wen_a40 = {1'b0, 1'b0};
                        wen_a39 = {1'b0, 1'b0};
                        wen_a38 = {1'b0, 1'b0};
                        wen_a37 = {1'b0, 1'b0};
                        wen_a36 = {1'b0, 1'b0};
                        wen_a35 = {1'b0, 1'b0};
                        wen_a34 = {1'b0, 1'b0};
                        wen_a33 = {1'b0, 1'b0};
                        wen_a32 = {1'b0, 1'b0};
                        wen_a31 = {1'b0, 1'b0};
                        wen_a30 = {1'b0, 1'b0};
                        wen_a29 = {1'b0, 1'b0};
                        wen_a28 = {1'b0, 1'b0};
                        wen_a27 = {1'b0, 1'b0};
                        wen_a26 = {1'b0, wen};
                        wen_a25 = {1'b0, wen};
                        wen_a24 = {1'b0, wen};
                        wen_a23 = {1'b0, wen};
                        wen_a22 = {1'b0, wen};
                        wen_a21 = {1'b0, wen};
                        wen_a20 = {1'b0, wen};
                        wen_a19 = {1'b0, wen};
                        wen_a18 = {1'b0, wen};
                        wen_a17 = {1'b0, wen};
                        wen_a16 = {1'b0, wen};
                        wen_a15 = {1'b0, wen};
                        wen_a14 = {1'b0, wen};
                        wen_a13 = {1'b0, wen};
                        wen_a12 = {1'b0, wen};
                        wen_a11 = {1'b0, wen};
                        wen_a10 = {1'b0, 1'b0};
                        wen_a9 = {1'b0, 1'b0};
                        wen_a8 = {1'b0, 1'b0};
                        wen_a7 = {1'b0, 1'b0};
                        wen_a6 = {1'b0, 1'b0};
                        wen_a5 = {1'b0, 1'b0};
                        wen_a4 = {1'b0, 1'b0};
                        wen_a3 = {1'b0, 1'b0};
                        wen_a2 = {1'b0, 1'b0};
                        wen_a1 = {1'b0, 1'b0};
                        wen_a0 = {1'b0, 1'b0};
                        wen_b0 = {1'b0, 1'b0};
                    end
                    6'b110000, 6'b110001, 6'b110010, 6'b110011,
                    6'b110100, 6'b110101, 6'b110110, 6'b110111 : begin
                        wen_a58 = {1'b0, 1'b0};
                        wen_a57 = {1'b0, 1'b0};
                        wen_a56 = {1'b0, 1'b0};
                        wen_a55 = {1'b0, 1'b0};
                        wen_a54 = {1'b0, 1'b0};
                        wen_a53 = {1'b0, 1'b0};
                        wen_a52 = {1'b0, 1'b0};
                        wen_a51 = {1'b0, 1'b0};
                        wen_a50 = {1'b0, 1'b0};
                        wen_a49 = {1'b0, 1'b0};
                        wen_a48 = {1'b0, 1'b0};
                        wen_a47 = {1'b0, 1'b0};
                        wen_a46 = {1'b0, 1'b0};
                        wen_a45 = {1'b0, 1'b0};
                        wen_a44 = {1'b0, 1'b0};
                        wen_a43 = {1'b0, 1'b0};
                        wen_a42 = {1'b0, 1'b0};
                        wen_a41 = {1'b0, 1'b0};
                        wen_a40 = {1'b0, 1'b0};
                        wen_a39 = {1'b0, 1'b0};
                        wen_a38 = {1'b0, 1'b0};
                        wen_a37 = {1'b0, 1'b0};
                        wen_a36 = {1'b0, 1'b0};
                        wen_a35 = {1'b0, 1'b0};
                        wen_a34 = {1'b0, 1'b0};
                        wen_a33 = {1'b0, 1'b0};
                        wen_a32 = {1'b0, 1'b0};
                        wen_a31 = {1'b0, 1'b0};
                        wen_a30 = {1'b0, 1'b0};
                        wen_a29 = {1'b0, 1'b0};
                        wen_a28 = {1'b0, 1'b0};
                        wen_a27 = {1'b0, 1'b0};
                        wen_a26 = {1'b0, 1'b0};
                        wen_a25 = {1'b0, 1'b0};
                        wen_a24 = {1'b0, 1'b0};
                        wen_a23 = {1'b0, 1'b0};
                        wen_a22 = {1'b0, 1'b0};
                        wen_a21 = {1'b0, 1'b0};
                        wen_a20 = {1'b0, 1'b0};
                        wen_a19 = {1'b0, 1'b0};
                        wen_a18 = {1'b0, 1'b0};
                        wen_a17 = {1'b0, 1'b0};
                        wen_a16 = {1'b0, 1'b0};
                        wen_a15 = {1'b0, 1'b0};
                        wen_a14 = {1'b0, 1'b0};
                        wen_a13 = {1'b0, 1'b0};
                        wen_a12 = {1'b0, 1'b0};
                        wen_a11 = {1'b0, 1'b0};
                        wen_a10 = {1'b0, wen};
                        wen_a9 = {1'b0, wen};
                        wen_a8 = {1'b0, wen};
                        wen_a7 = {1'b0, wen};
                        wen_a6 = {1'b0, wen};
                        wen_a5 = {1'b0, wen};
                        wen_a4 = {1'b0, wen};
                        wen_a3 = {1'b0, wen};
                        wen_a2 = {1'b0, 1'b0};
                        wen_a1 = {1'b0, 1'b0};
                        wen_a0 = {1'b0, 1'b0};
                        wen_b0 = {1'b0, 1'b0};
                    end
                    6'b111000, 6'b111001 : begin
                        wen_a58 = {1'b0, 1'b0};
                        wen_a57 = {1'b0, 1'b0};
                        wen_a56 = {1'b0, 1'b0};
                        wen_a55 = {1'b0, 1'b0};
                        wen_a54 = {1'b0, 1'b0};
                        wen_a53 = {1'b0, 1'b0};
                        wen_a52 = {1'b0, 1'b0};
                        wen_a51 = {1'b0, 1'b0};
                        wen_a50 = {1'b0, 1'b0};
                        wen_a49 = {1'b0, 1'b0};
                        wen_a48 = {1'b0, 1'b0};
                        wen_a47 = {1'b0, 1'b0};
                        wen_a46 = {1'b0, 1'b0};
                        wen_a45 = {1'b0, 1'b0};
                        wen_a44 = {1'b0, 1'b0};
                        wen_a43 = {1'b0, 1'b0};
                        wen_a42 = {1'b0, 1'b0};
                        wen_a41 = {1'b0, 1'b0};
                        wen_a40 = {1'b0, 1'b0};
                        wen_a39 = {1'b0, 1'b0};
                        wen_a38 = {1'b0, 1'b0};
                        wen_a37 = {1'b0, 1'b0};
                        wen_a36 = {1'b0, 1'b0};
                        wen_a35 = {1'b0, 1'b0};
                        wen_a34 = {1'b0, 1'b0};
                        wen_a33 = {1'b0, 1'b0};
                        wen_a32 = {1'b0, 1'b0};
                        wen_a31 = {1'b0, 1'b0};
                        wen_a30 = {1'b0, 1'b0};
                        wen_a29 = {1'b0, 1'b0};
                        wen_a28 = {1'b0, 1'b0};
                        wen_a27 = {1'b0, 1'b0};
                        wen_a26 = {1'b0, 1'b0};
                        wen_a25 = {1'b0, 1'b0};
                        wen_a24 = {1'b0, 1'b0};
                        wen_a23 = {1'b0, 1'b0};
                        wen_a22 = {1'b0, 1'b0};
                        wen_a21 = {1'b0, 1'b0};
                        wen_a20 = {1'b0, 1'b0};
                        wen_a19 = {1'b0, 1'b0};
                        wen_a18 = {1'b0, 1'b0};
                        wen_a17 = {1'b0, 1'b0};
                        wen_a16 = {1'b0, 1'b0};
                        wen_a15 = {1'b0, 1'b0};
                        wen_a14 = {1'b0, 1'b0};
                        wen_a13 = {1'b0, 1'b0};
                        wen_a12 = {1'b0, 1'b0};
                        wen_a11 = {1'b0, 1'b0};
                        wen_a10 = {1'b0, 1'b0};
                        wen_a9 = {1'b0, 1'b0};
                        wen_a8 = {1'b0, 1'b0};
                        wen_a7 = {1'b0, 1'b0};
                        wen_a6 = {1'b0, 1'b0};
                        wen_a5 = {1'b0, 1'b0};
                        wen_a4 = {1'b0, 1'b0};
                        wen_a3 = {1'b0, 1'b0};
                        wen_a2 = {wen, wen};
                        wen_a1 = {wen, wen};
                        wen_a0 = {1'b0, 1'b0};
                        wen_b0 = {1'b0, 1'b0};
                    end
                    6'b111010 : begin
                        wen_a58 = {1'b0, 1'b0};
                        wen_a57 = {1'b0, 1'b0};
                        wen_a56 = {1'b0, 1'b0};
                        wen_a55 = {1'b0, 1'b0};
                        wen_a54 = {1'b0, 1'b0};
                        wen_a53 = {1'b0, 1'b0};
                        wen_a52 = {1'b0, 1'b0};
                        wen_a51 = {1'b0, 1'b0};
                        wen_a50 = {1'b0, 1'b0};
                        wen_a49 = {1'b0, 1'b0};
                        wen_a48 = {1'b0, 1'b0};
                        wen_a47 = {1'b0, 1'b0};
                        wen_a46 = {1'b0, 1'b0};
                        wen_a45 = {1'b0, 1'b0};
                        wen_a44 = {1'b0, 1'b0};
                        wen_a43 = {1'b0, 1'b0};
                        wen_a42 = {1'b0, 1'b0};
                        wen_a41 = {1'b0, 1'b0};
                        wen_a40 = {1'b0, 1'b0};
                        wen_a39 = {1'b0, 1'b0};
                        wen_a38 = {1'b0, 1'b0};
                        wen_a37 = {1'b0, 1'b0};
                        wen_a36 = {1'b0, 1'b0};
                        wen_a35 = {1'b0, 1'b0};
                        wen_a34 = {1'b0, 1'b0};
                        wen_a33 = {1'b0, 1'b0};
                        wen_a32 = {1'b0, 1'b0};
                        wen_a31 = {1'b0, 1'b0};
                        wen_a30 = {1'b0, 1'b0};
                        wen_a29 = {1'b0, 1'b0};
                        wen_a28 = {1'b0, 1'b0};
                        wen_a27 = {1'b0, 1'b0};
                        wen_a26 = {1'b0, 1'b0};
                        wen_a25 = {1'b0, 1'b0};
                        wen_a24 = {1'b0, 1'b0};
                        wen_a23 = {1'b0, 1'b0};
                        wen_a22 = {1'b0, 1'b0};
                        wen_a21 = {1'b0, 1'b0};
                        wen_a20 = {1'b0, 1'b0};
                        wen_a19 = {1'b0, 1'b0};
                        wen_a18 = {1'b0, 1'b0};
                        wen_a17 = {1'b0, 1'b0};
                        wen_a16 = {1'b0, 1'b0};
                        wen_a15 = {1'b0, 1'b0};
                        wen_a14 = {1'b0, 1'b0};
                        wen_a13 = {1'b0, 1'b0};
                        wen_a12 = {1'b0, 1'b0};
                        wen_a11 = {1'b0, 1'b0};
                        wen_a10 = {1'b0, 1'b0};
                        wen_a9 = {1'b0, 1'b0};
                        wen_a8 = {1'b0, 1'b0};
                        wen_a7 = {1'b0, 1'b0};
                        wen_a6 = {1'b0, 1'b0};
                        wen_a5 = {1'b0, 1'b0};
                        wen_a4 = {1'b0, 1'b0};
                        wen_a3 = {1'b0, 1'b0};
                        wen_a2 = {1'b0, 1'b0};
                        wen_a1 = {1'b0, 1'b0};
                        wen_a0 = {wen, wen};
                        wen_b0 = {wen, wen};
                    end
                    default : begin
                        wen_a58 = {1'b0, 1'b0};
                        wen_a57 = {1'b0, 1'b0};
                        wen_a56 = {1'b0, 1'b0};
                        wen_a55 = {1'b0, 1'b0};
                        wen_a54 = {1'b0, 1'b0};
                        wen_a53 = {1'b0, 1'b0};
                        wen_a52 = {1'b0, 1'b0};
                        wen_a51 = {1'b0, 1'b0};
                        wen_a50 = {1'b0, 1'b0};
                        wen_a49 = {1'b0, 1'b0};
                        wen_a48 = {1'b0, 1'b0};
                        wen_a47 = {1'b0, 1'b0};
                        wen_a46 = {1'b0, 1'b0};
                        wen_a45 = {1'b0, 1'b0};
                        wen_a44 = {1'b0, 1'b0};
                        wen_a43 = {1'b0, 1'b0};
                        wen_a42 = {1'b0, 1'b0};
                        wen_a41 = {1'b0, 1'b0};
                        wen_a40 = {1'b0, 1'b0};
                        wen_a39 = {1'b0, 1'b0};
                        wen_a38 = {1'b0, 1'b0};
                        wen_a37 = {1'b0, 1'b0};
                        wen_a36 = {1'b0, 1'b0};
                        wen_a35 = {1'b0, 1'b0};
                        wen_a34 = {1'b0, 1'b0};
                        wen_a33 = {1'b0, 1'b0};
                        wen_a32 = {1'b0, 1'b0};
                        wen_a31 = {1'b0, 1'b0};
                        wen_a30 = {1'b0, 1'b0};
                        wen_a29 = {1'b0, 1'b0};
                        wen_a28 = {1'b0, 1'b0};
                        wen_a27 = {1'b0, 1'b0};
                        wen_a26 = {1'b0, 1'b0};
                        wen_a25 = {1'b0, 1'b0};
                        wen_a24 = {1'b0, 1'b0};
                        wen_a23 = {1'b0, 1'b0};
                        wen_a22 = {1'b0, 1'b0};
                        wen_a21 = {1'b0, 1'b0};
                        wen_a20 = {1'b0, 1'b0};
                        wen_a19 = {1'b0, 1'b0};
                        wen_a18 = {1'b0, 1'b0};
                        wen_a17 = {1'b0, 1'b0};
                        wen_a16 = {1'b0, 1'b0};
                        wen_a15 = {1'b0, 1'b0};
                        wen_a14 = {1'b0, 1'b0};
                        wen_a13 = {1'b0, 1'b0};
                        wen_a12 = {1'b0, 1'b0};
                        wen_a11 = {1'b0, 1'b0};
                        wen_a10 = {1'b0, 1'b0};
                        wen_a9 = {1'b0, 1'b0};
                        wen_a8 = {1'b0, 1'b0};
                        wen_a7 = {1'b0, 1'b0};
                        wen_a6 = {1'b0, 1'b0};
                        wen_a5 = {1'b0, 1'b0};
                        wen_a4 = {1'b0, 1'b0};
                        wen_a3 = {1'b0, 1'b0};
                        wen_a2 = {1'b0, 1'b0};
                        wen_a1 = {1'b0, 1'b0};
                        wen_a0 = {1'b0, 1'b0};
                        wen_b0 = {1'b0, 1'b0};
                    end
                endcase

                case (ckRdAddr[14:9])
                    6'b000000, 6'b000001, 6'b000010, 6'b000011,
                    6'b000100, 6'b000101, 6'b000110, 6'b000111,
                    6'b001000, 6'b001001, 6'b001010, 6'b001011,
                    6'b001100, 6'b001101, 6'b001110, 6'b001111,
                    6'b010000, 6'b010001, 6'b010010, 6'b010011,
                    6'b010100, 6'b010101, 6'b010110, 6'b010111,
                    6'b011000, 6'b011001, 6'b011010, 6'b011011,
                    6'b011100, 6'b011101, 6'b011110, 6'b011111 : begin
                        readData = {
                                        readData58[0],
                                        readData57[0],
                                        readData56[0],
                                        readData55[0],
                                        readData54[0],
                                        readData53[0],
                                        readData52[0],
                                        readData51[0],
                                        readData50[0],
                                        readData49[0],
                                        readData48[0],
                                        readData47[0],
                                        readData46[0],
                                        readData45[0],
                                        readData44[0],
                                        readData43[0],
                                        readData42[0],
                                        readData41[0],
                                        readData40[0],
                                        readData39[0],
                                        readData38[0],
                                        readData37[0],
                                        readData36[0],
                                        readData35[0],
                                        readData34[0],
                                        readData33[0],
                                        readData32[0],
                                        readData31[0],
                                        readData30[0],
                                        readData29[0],
                                        readData28[0],
                                        readData27[0]
                        };
                    end
                    6'b100000, 6'b100001, 6'b100010, 6'b100011,
                    6'b100100, 6'b100101, 6'b100110, 6'b100111,
                    6'b101000, 6'b101001, 6'b101010, 6'b101011,
                    6'b101100, 6'b101101, 6'b101110, 6'b101111 : begin
                        readData = {
                                        readData26[1:0],
                                        readData25[1:0],
                                        readData24[1:0],
                                        readData23[1:0],
                                        readData22[1:0],
                                        readData21[1:0],
                                        readData20[1:0],
                                        readData19[1:0],
                                        readData18[1:0],
                                        readData17[1:0],
                                        readData16[1:0],
                                        readData15[1:0],
                                        readData14[1:0],
                                        readData13[1:0],
                                        readData12[1:0],
                                        readData11[1:0]
                        };
                    end
                    6'b110000, 6'b110001, 6'b110010, 6'b110011,
                    6'b110100, 6'b110101, 6'b110110, 6'b110111 : begin
                        readData = {
                                        readData10[3:0],
                                        readData9[3:0],
                                        readData8[3:0],
                                        readData7[3:0],
                                        readData6[3:0],
                                        readData5[3:0],
                                        readData4[3:0],
                                        readData3[3:0]
                        };
                    end
                    6'b111000, 6'b111001 : begin
                        readData = {readData2[16:9],readData2[7:0],readData1[16:9],readData1[7:0]};
                    end
                    6'b111010 : begin
                        readData = {readData0[34:27],readData0[25:18],readData0[16:9],readData0[7:0]};
                    end
                    default : begin
                        readData = 32'b0;
                    end
                endcase
            end        
            30720: begin
                width60 = 3'b000;
                width59 = 3'b000;
                width58 = 3'b000;
                width57 = 3'b000;
                width56 = 3'b000;
                width55 = 3'b000;
                width54 = 3'b000;
                width53 = 3'b000;
                width52 = 3'b000;
                width51 = 3'b000;
                width50 = 3'b000;
                width49 = 3'b000;
                width48 = 3'b000;
                width47 = 3'b000;
                width46 = 3'b000;
                width45 = 3'b000;
                width44 = 3'b000;
                width43 = 3'b000;
                width42 = 3'b000;
                width41 = 3'b000;
                width40 = 3'b000;
                width39 = 3'b000;
                width38 = 3'b000;
                width37 = 3'b000;
                width36 = 3'b000;
                width35 = 3'b000;
                width34 = 3'b000;
                width33 = 3'b000;
                width32 = 3'b000;
                width31 = 3'b000;
                width30 = 3'b000;
                width29 = 3'b000;
                width28 = 3'b001;
                width27 = 3'b001;
                width26 = 3'b001;
                width25 = 3'b001;
                width24 = 3'b001;
                width23 = 3'b001;
                width22 = 3'b001;
                width21 = 3'b001;
                width20 = 3'b001;
                width19 = 3'b001;
                width18 = 3'b001;
                width17 = 3'b001;
                width16 = 3'b001;
                width15 = 3'b001;
                width14 = 3'b001;
                width13 = 3'b001;
                width12 = 3'b010;
                width11 = 3'b010;
                width10 = 3'b010;
                width9 = 3'b010;
                width8 = 3'b010;
                width7 = 3'b010;
                width6 = 3'b010;
                width5 = 3'b010;
                width4 = 3'b011;
                width3 = 3'b011;
                width2 = 3'b011;
                width1 = 3'b011;

                writeAddr60 = {writeAddr[13:0]};
                writeAddr59 = {writeAddr[13:0]};
                writeAddr58 = {writeAddr[13:0]};
                writeAddr57 = {writeAddr[13:0]};
                writeAddr56 = {writeAddr[13:0]};
                writeAddr55 = {writeAddr[13:0]};
                writeAddr54 = {writeAddr[13:0]};
                writeAddr53 = {writeAddr[13:0]};
                writeAddr52 = {writeAddr[13:0]};
                writeAddr51 = {writeAddr[13:0]};
                writeAddr50 = {writeAddr[13:0]};
                writeAddr49 = {writeAddr[13:0]};
                writeAddr48 = {writeAddr[13:0]};
                writeAddr47 = {writeAddr[13:0]};
                writeAddr46 = {writeAddr[13:0]};
                writeAddr45 = {writeAddr[13:0]};
                writeAddr44 = {writeAddr[13:0]};
                writeAddr43 = {writeAddr[13:0]};
                writeAddr42 = {writeAddr[13:0]};
                writeAddr41 = {writeAddr[13:0]};
                writeAddr40 = {writeAddr[13:0]};
                writeAddr39 = {writeAddr[13:0]};
                writeAddr38 = {writeAddr[13:0]};
                writeAddr37 = {writeAddr[13:0]};
                writeAddr36 = {writeAddr[13:0]};
                writeAddr35 = {writeAddr[13:0]};
                writeAddr34 = {writeAddr[13:0]};
                writeAddr33 = {writeAddr[13:0]};
                writeAddr32 = {writeAddr[13:0]};
                writeAddr31 = {writeAddr[13:0]};
                writeAddr30 = {writeAddr[13:0]};
                writeAddr29 = {writeAddr[13:0]};
                writeAddr28 = {writeAddr[12:0], 1'b0};
                writeAddr27 = {writeAddr[12:0], 1'b0};
                writeAddr26 = {writeAddr[12:0], 1'b0};
                writeAddr25 = {writeAddr[12:0], 1'b0};
                writeAddr24 = {writeAddr[12:0], 1'b0};
                writeAddr23 = {writeAddr[12:0], 1'b0};
                writeAddr22 = {writeAddr[12:0], 1'b0};
                writeAddr21 = {writeAddr[12:0], 1'b0};
                writeAddr20 = {writeAddr[12:0], 1'b0};
                writeAddr19 = {writeAddr[12:0], 1'b0};
                writeAddr18 = {writeAddr[12:0], 1'b0};
                writeAddr17 = {writeAddr[12:0], 1'b0};
                writeAddr16 = {writeAddr[12:0], 1'b0};
                writeAddr15 = {writeAddr[12:0], 1'b0};
                writeAddr14 = {writeAddr[12:0], 1'b0};
                writeAddr13 = {writeAddr[12:0], 1'b0};
                writeAddr12 = {writeAddr[11:0], 2'b0};
                writeAddr11 = {writeAddr[11:0], 2'b0};
                writeAddr10 = {writeAddr[11:0], 2'b0};
                writeAddr9 = {writeAddr[11:0], 2'b0};
                writeAddr8 = {writeAddr[11:0], 2'b0};
                writeAddr7 = {writeAddr[11:0], 2'b0};
                writeAddr6 = {writeAddr[11:0], 2'b0};
                writeAddr5 = {writeAddr[11:0], 2'b0};
                writeAddr4 = {writeAddr[10:0], 3'b0};
                writeAddr3 = {writeAddr[10:0], 3'b0};
                writeAddr2 = {writeAddr[10:0], 3'b0};
                writeAddr1 = {writeAddr[10:0], 3'b0};

                readAddr60 = {writeAddr[13:0]};
                readAddr59 = {writeAddr[13:0]};
                readAddr58 = {writeAddr[13:0]};
                readAddr57 = {writeAddr[13:0]};
                readAddr56 = {writeAddr[13:0]};
                readAddr55 = {writeAddr[13:0]};
                readAddr54 = {writeAddr[13:0]};
                readAddr53 = {writeAddr[13:0]};
                readAddr52 = {writeAddr[13:0]};
                readAddr51 = {writeAddr[13:0]};
                readAddr50 = {writeAddr[13:0]};
                readAddr49 = {writeAddr[13:0]};
                readAddr48 = {writeAddr[13:0]};
                readAddr47 = {writeAddr[13:0]};
                readAddr46 = {writeAddr[13:0]};
                readAddr45 = {writeAddr[13:0]};
                readAddr44 = {writeAddr[13:0]};
                readAddr43 = {writeAddr[13:0]};
                readAddr42 = {writeAddr[13:0]};
                readAddr41 = {writeAddr[13:0]};
                readAddr40 = {writeAddr[13:0]};
                readAddr39 = {writeAddr[13:0]};
                readAddr38 = {writeAddr[13:0]};
                readAddr37 = {writeAddr[13:0]};
                readAddr36 = {writeAddr[13:0]};
                readAddr35 = {writeAddr[13:0]};
                readAddr34 = {writeAddr[13:0]};
                readAddr33 = {writeAddr[13:0]};
                readAddr32 = {writeAddr[13:0]};
                readAddr31 = {writeAddr[13:0]};
                readAddr30 = {writeAddr[13:0]};
                readAddr29 = {writeAddr[13:0]};
                readAddr28  = {readAddr[12:0],  1'b0};
                readAddr27  = {readAddr[12:0],  1'b0};
                readAddr26  = {readAddr[12:0],  1'b0};
                readAddr25  = {readAddr[12:0],  1'b0};
                readAddr24  = {readAddr[12:0],  1'b0};
                readAddr23  = {readAddr[12:0],  1'b0};
                readAddr22  = {readAddr[12:0],  1'b0};
                readAddr21  = {readAddr[12:0],  1'b0};
                readAddr20  = {readAddr[12:0],  1'b0};
                readAddr19  = {readAddr[12:0],  1'b0};
                readAddr18  = {readAddr[12:0],  1'b0};
                readAddr17  = {readAddr[12:0],  1'b0};
                readAddr16  = {readAddr[12:0],  1'b0};
                readAddr15  = {readAddr[12:0],  1'b0};
                readAddr14  = {readAddr[12:0],  1'b0};
                readAddr13  = {readAddr[12:0],  1'b0};
                readAddr12  = {readAddr[11:0],  2'b0};
                readAddr11  = {readAddr[11:0],  2'b0};
                readAddr10  = {readAddr[11:0],  2'b0};
                readAddr9  = {readAddr[11:0],  2'b0};
                readAddr8  = {readAddr[11:0],  2'b0};
                readAddr7  = {readAddr[11:0],  2'b0};
                readAddr6  = {readAddr[11:0],  2'b0};
                readAddr5  = {readAddr[11:0],  2'b0};
                readAddr4  = {readAddr[10:0],  3'b0};
                readAddr3  = {readAddr[10:0],  3'b0};
                readAddr2  = {readAddr[10:0],  3'b0};
                readAddr1  = {readAddr[10:0],  3'b0};

                writeData60 = {17'b0, writeData[31]};
                writeData59 = {17'b0, writeData[30]};
                writeData58 = {17'b0, writeData[29]};
                writeData57 = {17'b0, writeData[28]};
                writeData56 = {17'b0, writeData[27]};
                writeData55 = {17'b0, writeData[26]};
                writeData54 = {17'b0, writeData[25]};
                writeData53 = {17'b0, writeData[24]};
                writeData52 = {17'b0, writeData[23]};
                writeData51 = {17'b0, writeData[22]};
                writeData50 = {17'b0, writeData[21]};
                writeData49 = {17'b0, writeData[20]};
                writeData48 = {17'b0, writeData[19]};
                writeData47 = {17'b0, writeData[18]};
                writeData46 = {17'b0, writeData[17]};
                writeData45 = {17'b0, writeData[16]};
                writeData44 = {17'b0, writeData[15]};
                writeData43 = {17'b0, writeData[14]};
                writeData42 = {17'b0, writeData[13]};
                writeData41 = {17'b0, writeData[12]};
                writeData40 = {17'b0, writeData[11]};
                writeData39 = {17'b0, writeData[10]};
                writeData38 = {17'b0, writeData[9]};
                writeData37 = {17'b0, writeData[8]};
                writeData36 = {17'b0, writeData[7]};
                writeData35 = {17'b0, writeData[6]};
                writeData34 = {17'b0, writeData[5]};
                writeData33 = {17'b0, writeData[4]};
                writeData32 = {17'b0, writeData[3]};
                writeData31 = {17'b0, writeData[2]};
                writeData30 = {17'b0, writeData[1]};
                writeData29 = {17'b0, writeData[0]};
                writeData28 = {16'b0, writeData[31:30]};
                writeData27 = {16'b0, writeData[29:28]};
                writeData26 = {16'b0, writeData[27:26]};
                writeData25 = {16'b0, writeData[25:24]};
                writeData24 = {16'b0, writeData[23:22]};
                writeData23 = {16'b0, writeData[21:20]};
                writeData22 = {16'b0, writeData[19:18]};
                writeData21 = {16'b0, writeData[17:16]};
                writeData20 = {16'b0, writeData[15:14]};
                writeData19 = {16'b0, writeData[13:12]};
                writeData18 = {16'b0, writeData[11:10]};
                writeData17 = {16'b0, writeData[9:8]};
                writeData16 = {16'b0, writeData[7:6]};
                writeData15 = {16'b0, writeData[5:4]};
                writeData14 = {16'b0, writeData[3:2]};
                writeData13 = {16'b0, writeData[1:0]};
                writeData12 = {14'b0, writeData[31:28]};
                writeData11 = {14'b0, writeData[27:24]};
                writeData10 = {14'b0, writeData[23:20]};
                writeData9 = {14'b0, writeData[19:16]};
                writeData8 = {14'b0, writeData[15:12]};
                writeData7 = {14'b0, writeData[11:8]};
                writeData6 = {14'b0, writeData[7:4]};
                writeData5 = {14'b0, writeData[3:0]};
                writeData4 = {10'b0, writeData[31:24]};
                writeData3 = {10'b0, writeData[23:16]};
                writeData2 = {10'b0, writeData[15:8]};
                writeData1 = {10'b0, writeData[7:0]};

                case (writeAddr[14:9])
                    6'b000000, 6'b000001, 6'b000010, 6'b000011,
                    6'b000100, 6'b000101, 6'b000110, 6'b000111,
                    6'b001000, 6'b001001, 6'b001010, 6'b001011,
                    6'b001100, 6'b001101, 6'b001110, 6'b001111,
                    6'b010000, 6'b010001, 6'b010010, 6'b010011,
                    6'b010100, 6'b010101, 6'b010110, 6'b010111,
                    6'b011000, 6'b011001, 6'b011010, 6'b011011,
                    6'b011100, 6'b011101, 6'b011110, 6'b011111 : begin
                        wen_a60 = {1'b0, wen};
                        wen_a59 = {1'b0, wen};
                        wen_a58 = {1'b0, wen};
                        wen_a57 = {1'b0, wen};
                        wen_a56 = {1'b0, wen};
                        wen_a55 = {1'b0, wen};
                        wen_a54 = {1'b0, wen};
                        wen_a53 = {1'b0, wen};
                        wen_a52 = {1'b0, wen};
                        wen_a51 = {1'b0, wen};
                        wen_a50 = {1'b0, wen};
                        wen_a49 = {1'b0, wen};
                        wen_a48 = {1'b0, wen};
                        wen_a47 = {1'b0, wen};
                        wen_a46 = {1'b0, wen};
                        wen_a45 = {1'b0, wen};
                        wen_a44 = {1'b0, wen};
                        wen_a43 = {1'b0, wen};
                        wen_a42 = {1'b0, wen};
                        wen_a41 = {1'b0, wen};
                        wen_a40 = {1'b0, wen};
                        wen_a39 = {1'b0, wen};
                        wen_a38 = {1'b0, wen};
                        wen_a37 = {1'b0, wen};
                        wen_a36 = {1'b0, wen};
                        wen_a35 = {1'b0, wen};
                        wen_a34 = {1'b0, wen};
                        wen_a33 = {1'b0, wen};
                        wen_a32 = {1'b0, wen};
                        wen_a31 = {1'b0, wen};
                        wen_a30 = {1'b0, wen};
                        wen_a29 = {1'b0, wen};
                        wen_a28 = {1'b0, 1'b0};
                        wen_a27 = {1'b0, 1'b0};
                        wen_a26 = {1'b0, 1'b0};
                        wen_a25 = {1'b0, 1'b0};
                        wen_a24 = {1'b0, 1'b0};
                        wen_a23 = {1'b0, 1'b0};
                        wen_a22 = {1'b0, 1'b0};
                        wen_a21 = {1'b0, 1'b0};
                        wen_a20 = {1'b0, 1'b0};
                        wen_a19 = {1'b0, 1'b0};
                        wen_a18 = {1'b0, 1'b0};
                        wen_a17 = {1'b0, 1'b0};
                        wen_a16 = {1'b0, 1'b0};
                        wen_a15 = {1'b0, 1'b0};
                        wen_a14 = {1'b0, 1'b0};
                        wen_a13 = {1'b0, 1'b0};
                        wen_a12 = {1'b0, 1'b0};
                        wen_a11 = {1'b0, 1'b0};
                        wen_a10 = {1'b0, 1'b0};
                        wen_a9 = {1'b0, 1'b0};
                        wen_a8 = {1'b0, 1'b0};
                        wen_a7 = {1'b0, 1'b0};
                        wen_a6 = {1'b0, 1'b0};
                        wen_a5 = {1'b0, 1'b0};
                        wen_a4 = {1'b0, 1'b0};
                        wen_a3 = {1'b0, 1'b0};
                        wen_a2 = {1'b0, 1'b0};
                        wen_a1 = {1'b0, 1'b0};
                    end
                    6'b100000, 6'b100001, 6'b100010, 6'b100011,
                    6'b100100, 6'b100101, 6'b100110, 6'b100111,
                    6'b101000, 6'b101001, 6'b101010, 6'b101011,
                    6'b101100, 6'b101101, 6'b101110, 6'b101111 : begin
                        wen_a60 = {1'b0, 1'b0};
                        wen_a59 = {1'b0, 1'b0};
                        wen_a58 = {1'b0, 1'b0};
                        wen_a57 = {1'b0, 1'b0};
                        wen_a56 = {1'b0, 1'b0};
                        wen_a55 = {1'b0, 1'b0};
                        wen_a54 = {1'b0, 1'b0};
                        wen_a53 = {1'b0, 1'b0};
                        wen_a52 = {1'b0, 1'b0};
                        wen_a51 = {1'b0, 1'b0};
                        wen_a50 = {1'b0, 1'b0};
                        wen_a49 = {1'b0, 1'b0};
                        wen_a48 = {1'b0, 1'b0};
                        wen_a47 = {1'b0, 1'b0};
                        wen_a46 = {1'b0, 1'b0};
                        wen_a45 = {1'b0, 1'b0};
                        wen_a44 = {1'b0, 1'b0};
                        wen_a43 = {1'b0, 1'b0};
                        wen_a42 = {1'b0, 1'b0};
                        wen_a41 = {1'b0, 1'b0};
                        wen_a40 = {1'b0, 1'b0};
                        wen_a39 = {1'b0, 1'b0};
                        wen_a38 = {1'b0, 1'b0};
                        wen_a37 = {1'b0, 1'b0};
                        wen_a36 = {1'b0, 1'b0};
                        wen_a35 = {1'b0, 1'b0};
                        wen_a34 = {1'b0, 1'b0};
                        wen_a33 = {1'b0, 1'b0};
                        wen_a32 = {1'b0, 1'b0};
                        wen_a31 = {1'b0, 1'b0};
                        wen_a30 = {1'b0, 1'b0};
                        wen_a29 = {1'b0, 1'b0};
                        wen_a28 = {1'b0, wen};
                        wen_a27 = {1'b0, wen};
                        wen_a26 = {1'b0, wen};
                        wen_a25 = {1'b0, wen};
                        wen_a24 = {1'b0, wen};
                        wen_a23 = {1'b0, wen};
                        wen_a22 = {1'b0, wen};
                        wen_a21 = {1'b0, wen};
                        wen_a20 = {1'b0, wen};
                        wen_a19 = {1'b0, wen};
                        wen_a18 = {1'b0, wen};
                        wen_a17 = {1'b0, wen};
                        wen_a16 = {1'b0, wen};
                        wen_a15 = {1'b0, wen};
                        wen_a14 = {1'b0, wen};
                        wen_a13 = {1'b0, wen};
                        wen_a12 = {1'b0, 1'b0};
                        wen_a11 = {1'b0, 1'b0};
                        wen_a10 = {1'b0, 1'b0};
                        wen_a9 = {1'b0, 1'b0};
                        wen_a8 = {1'b0, 1'b0};
                        wen_a7 = {1'b0, 1'b0};
                        wen_a6 = {1'b0, 1'b0};
                        wen_a5 = {1'b0, 1'b0};
                        wen_a4 = {1'b0, 1'b0};
                        wen_a3 = {1'b0, 1'b0};
                        wen_a2 = {1'b0, 1'b0};
                        wen_a1 = {1'b0, 1'b0};
                    end
                    6'b110000, 6'b110001, 6'b110010, 6'b110011,
                    6'b110100, 6'b110101, 6'b110110, 6'b110111 : begin
                        wen_a60 = {1'b0, 1'b0};
                        wen_a59 = {1'b0, 1'b0};
                        wen_a58 = {1'b0, 1'b0};
                        wen_a57 = {1'b0, 1'b0};
                        wen_a56 = {1'b0, 1'b0};
                        wen_a55 = {1'b0, 1'b0};
                        wen_a54 = {1'b0, 1'b0};
                        wen_a53 = {1'b0, 1'b0};
                        wen_a52 = {1'b0, 1'b0};
                        wen_a51 = {1'b0, 1'b0};
                        wen_a50 = {1'b0, 1'b0};
                        wen_a49 = {1'b0, 1'b0};
                        wen_a48 = {1'b0, 1'b0};
                        wen_a47 = {1'b0, 1'b0};
                        wen_a46 = {1'b0, 1'b0};
                        wen_a45 = {1'b0, 1'b0};
                        wen_a44 = {1'b0, 1'b0};
                        wen_a43 = {1'b0, 1'b0};
                        wen_a42 = {1'b0, 1'b0};
                        wen_a41 = {1'b0, 1'b0};
                        wen_a40 = {1'b0, 1'b0};
                        wen_a39 = {1'b0, 1'b0};
                        wen_a38 = {1'b0, 1'b0};
                        wen_a37 = {1'b0, 1'b0};
                        wen_a36 = {1'b0, 1'b0};
                        wen_a35 = {1'b0, 1'b0};
                        wen_a34 = {1'b0, 1'b0};
                        wen_a33 = {1'b0, 1'b0};
                        wen_a32 = {1'b0, 1'b0};
                        wen_a31 = {1'b0, 1'b0};
                        wen_a30 = {1'b0, 1'b0};
                        wen_a29 = {1'b0, 1'b0};
                        wen_a28 = {1'b0, 1'b0};
                        wen_a27 = {1'b0, 1'b0};
                        wen_a26 = {1'b0, 1'b0};
                        wen_a25 = {1'b0, 1'b0};
                        wen_a24 = {1'b0, 1'b0};
                        wen_a23 = {1'b0, 1'b0};
                        wen_a22 = {1'b0, 1'b0};
                        wen_a21 = {1'b0, 1'b0};
                        wen_a20 = {1'b0, 1'b0};
                        wen_a19 = {1'b0, 1'b0};
                        wen_a18 = {1'b0, 1'b0};
                        wen_a17 = {1'b0, 1'b0};
                        wen_a16 = {1'b0, 1'b0};
                        wen_a15 = {1'b0, 1'b0};
                        wen_a14 = {1'b0, 1'b0};
                        wen_a13 = {1'b0, 1'b0};
                        wen_a12 = {1'b0, wen};
                        wen_a11 = {1'b0, wen};
                        wen_a10 = {1'b0, wen};
                        wen_a9 = {1'b0, wen};
                        wen_a8 = {1'b0, wen};
                        wen_a7 = {1'b0, wen};
                        wen_a6 = {1'b0, wen};
                        wen_a5 = {1'b0, wen};
                        wen_a4 = {1'b0, 1'b0};
                        wen_a3 = {1'b0, 1'b0};
                        wen_a2 = {1'b0, 1'b0};
                        wen_a1 = {1'b0, 1'b0};
                    end
                    6'b111000, 6'b111001, 6'b111010, 6'b111011 : begin
                        wen_a60 = {1'b0, 1'b0};
                        wen_a59 = {1'b0, 1'b0};
                        wen_a58 = {1'b0, 1'b0};
                        wen_a57 = {1'b0, 1'b0};
                        wen_a56 = {1'b0, 1'b0};
                        wen_a55 = {1'b0, 1'b0};
                        wen_a54 = {1'b0, 1'b0};
                        wen_a53 = {1'b0, 1'b0};
                        wen_a52 = {1'b0, 1'b0};
                        wen_a51 = {1'b0, 1'b0};
                        wen_a50 = {1'b0, 1'b0};
                        wen_a49 = {1'b0, 1'b0};
                        wen_a48 = {1'b0, 1'b0};
                        wen_a47 = {1'b0, 1'b0};
                        wen_a46 = {1'b0, 1'b0};
                        wen_a45 = {1'b0, 1'b0};
                        wen_a44 = {1'b0, 1'b0};
                        wen_a43 = {1'b0, 1'b0};
                        wen_a42 = {1'b0, 1'b0};
                        wen_a41 = {1'b0, 1'b0};
                        wen_a40 = {1'b0, 1'b0};
                        wen_a39 = {1'b0, 1'b0};
                        wen_a38 = {1'b0, 1'b0};
                        wen_a37 = {1'b0, 1'b0};
                        wen_a36 = {1'b0, 1'b0};
                        wen_a35 = {1'b0, 1'b0};
                        wen_a34 = {1'b0, 1'b0};
                        wen_a33 = {1'b0, 1'b0};
                        wen_a32 = {1'b0, 1'b0};
                        wen_a31 = {1'b0, 1'b0};
                        wen_a30 = {1'b0, 1'b0};
                        wen_a29 = {1'b0, 1'b0};
                        wen_a28 = {1'b0, 1'b0};
                        wen_a27 = {1'b0, 1'b0};
                        wen_a26 = {1'b0, 1'b0};
                        wen_a25 = {1'b0, 1'b0};
                        wen_a24 = {1'b0, 1'b0};
                        wen_a23 = {1'b0, 1'b0};
                        wen_a22 = {1'b0, 1'b0};
                        wen_a21 = {1'b0, 1'b0};
                        wen_a20 = {1'b0, 1'b0};
                        wen_a19 = {1'b0, 1'b0};
                        wen_a18 = {1'b0, 1'b0};
                        wen_a17 = {1'b0, 1'b0};
                        wen_a16 = {1'b0, 1'b0};
                        wen_a15 = {1'b0, 1'b0};
                        wen_a14 = {1'b0, 1'b0};
                        wen_a13 = {1'b0, 1'b0};
                        wen_a12 = {1'b0, 1'b0};
                        wen_a11 = {1'b0, 1'b0};
                        wen_a10 = {1'b0, 1'b0};
                        wen_a9 = {1'b0, 1'b0};
                        wen_a8 = {1'b0, 1'b0};
                        wen_a7 = {1'b0, 1'b0};
                        wen_a6 = {1'b0, 1'b0};
                        wen_a5 = {1'b0, 1'b0};
                        wen_a4 = {1'b0, wen};
                        wen_a3 = {1'b0, wen};
                        wen_a2 = {1'b0, wen};
                        wen_a1 = {1'b0, wen};
                    end
                    default : begin
                        wen_a60 = {1'b0, 1'b0};
                        wen_a59 = {1'b0, 1'b0};
                        wen_a58 = {1'b0, 1'b0};
                        wen_a57 = {1'b0, 1'b0};
                        wen_a56 = {1'b0, 1'b0};
                        wen_a55 = {1'b0, 1'b0};
                        wen_a54 = {1'b0, 1'b0};
                        wen_a53 = {1'b0, 1'b0};
                        wen_a52 = {1'b0, 1'b0};
                        wen_a51 = {1'b0, 1'b0};
                        wen_a50 = {1'b0, 1'b0};
                        wen_a49 = {1'b0, 1'b0};
                        wen_a48 = {1'b0, 1'b0};
                        wen_a47 = {1'b0, 1'b0};
                        wen_a46 = {1'b0, 1'b0};
                        wen_a45 = {1'b0, 1'b0};
                        wen_a44 = {1'b0, 1'b0};
                        wen_a43 = {1'b0, 1'b0};
                        wen_a42 = {1'b0, 1'b0};
                        wen_a41 = {1'b0, 1'b0};
                        wen_a40 = {1'b0, 1'b0};
                        wen_a39 = {1'b0, 1'b0};
                        wen_a38 = {1'b0, 1'b0};
                        wen_a37 = {1'b0, 1'b0};
                        wen_a36 = {1'b0, 1'b0};
                        wen_a35 = {1'b0, 1'b0};
                        wen_a34 = {1'b0, 1'b0};
                        wen_a33 = {1'b0, 1'b0};
                        wen_a32 = {1'b0, 1'b0};
                        wen_a31 = {1'b0, 1'b0};
                        wen_a30 = {1'b0, 1'b0};
                        wen_a29 = {1'b0, 1'b0};
                        wen_a28 = {1'b0, 1'b0};
                        wen_a27 = {1'b0, 1'b0};
                        wen_a26 = {1'b0, 1'b0};
                        wen_a25 = {1'b0, 1'b0};
                        wen_a24 = {1'b0, 1'b0};
                        wen_a23 = {1'b0, 1'b0};
                        wen_a22 = {1'b0, 1'b0};
                        wen_a21 = {1'b0, 1'b0};
                        wen_a20 = {1'b0, 1'b0};
                        wen_a19 = {1'b0, 1'b0};
                        wen_a18 = {1'b0, 1'b0};
                        wen_a17 = {1'b0, 1'b0};
                        wen_a16 = {1'b0, 1'b0};
                        wen_a15 = {1'b0, 1'b0};
                        wen_a14 = {1'b0, 1'b0};
                        wen_a13 = {1'b0, 1'b0};
                        wen_a12 = {1'b0, 1'b0};
                        wen_a11 = {1'b0, 1'b0};
                        wen_a10 = {1'b0, 1'b0};
                        wen_a9 = {1'b0, 1'b0};
                        wen_a8 = {1'b0, 1'b0};
                        wen_a7 = {1'b0, 1'b0};
                        wen_a6 = {1'b0, 1'b0};
                        wen_a5 = {1'b0, 1'b0};
                        wen_a4 = {1'b0, 1'b0};
                        wen_a3 = {1'b0, 1'b0};
                        wen_a2 = {1'b0, 1'b0};
                        wen_a1 = {1'b0, 1'b0};
                    end
                endcase

                case (ckRdAddr[14:9])
                    6'b000000, 6'b000001, 6'b000010, 6'b000011,
                    6'b000100, 6'b000101, 6'b000110, 6'b000111,
                    6'b001000, 6'b001001, 6'b001010, 6'b001011,
                    6'b001100, 6'b001101, 6'b001110, 6'b001111,
                    6'b010000, 6'b010001, 6'b010010, 6'b010011,
                    6'b010100, 6'b010101, 6'b010110, 6'b010111,
                    6'b011000, 6'b011001, 6'b011010, 6'b011011,
                    6'b011100, 6'b011101, 6'b011110, 6'b011111 : begin
                        readData = {
                                        readData60[0],
                                        readData59[0],
                                        readData58[0],
                                        readData57[0],
                                        readData56[0],
                                        readData55[0],
                                        readData54[0],
                                        readData53[0],
                                        readData52[0],
                                        readData51[0],
                                        readData50[0],
                                        readData49[0],
                                        readData48[0],
                                        readData47[0],
                                        readData46[0],
                                        readData45[0],
                                        readData44[0],
                                        readData43[0],
                                        readData42[0],
                                        readData41[0],
                                        readData40[0],
                                        readData39[0],
                                        readData38[0],
                                        readData37[0],
                                        readData36[0],
                                        readData35[0],
                                        readData34[0],
                                        readData33[0],
                                        readData32[0],
                                        readData31[0],
                                        readData30[0],
                                        readData29[0]
                        };
                    end
                    6'b100000, 6'b100001, 6'b100010, 6'b100011,
                    6'b100100, 6'b100101, 6'b100110, 6'b100111,
                    6'b101000, 6'b101001, 6'b101010, 6'b101011,
                    6'b101100, 6'b101101, 6'b101110, 6'b101111 : begin
                        readData = {
                                        readData28[1:0],
                                        readData27[1:0],
                                        readData26[1:0],
                                        readData25[1:0],
                                        readData24[1:0],
                                        readData23[1:0],
                                        readData22[1:0],
                                        readData21[1:0],
                                        readData20[1:0],
                                        readData19[1:0],
                                        readData18[1:0],
                                        readData17[1:0],
                                        readData16[1:0],
                                        readData15[1:0],
                                        readData14[1:0],
                                        readData13[1:0]
                        };
                    end
                    6'b110000, 6'b110001, 6'b110010, 6'b110011,
                    6'b110100, 6'b110101, 6'b110110, 6'b110111 : begin
                        readData = {
                                        readData12[3:0],
                                        readData11[3:0],
                                        readData10[3:0],
                                        readData9[3:0],
                                        readData8[3:0],
                                        readData7[3:0],
                                        readData6[3:0],
                                        readData5[3:0]
                        };
                    end
                    6'b111000, 6'b111001, 6'b111010, 6'b111011 : begin
                        readData = {readData4[7:0],readData3[7:0],readData2[7:0],readData1[7:0]};
                    end
                    default : begin
                        readData = 32'b0;
                    end
                endcase
            end        
            31232: begin
                width60 = 3'b000;
                width59 = 3'b000;
                width58 = 3'b000;
                width57 = 3'b000;
                width56 = 3'b000;
                width55 = 3'b000;
                width54 = 3'b000;
                width53 = 3'b000;
                width52 = 3'b000;
                width51 = 3'b000;
                width50 = 3'b000;
                width49 = 3'b000;
                width48 = 3'b000;
                width47 = 3'b000;
                width46 = 3'b000;
                width45 = 3'b000;
                width44 = 3'b000;
                width43 = 3'b000;
                width42 = 3'b000;
                width41 = 3'b000;
                width40 = 3'b000;
                width39 = 3'b000;
                width38 = 3'b000;
                width37 = 3'b000;
                width36 = 3'b000;
                width35 = 3'b000;
                width34 = 3'b000;
                width33 = 3'b000;
                width32 = 3'b000;
                width31 = 3'b000;
                width30 = 3'b000;
                width29 = 3'b000;
                width28 = 3'b001;
                width27 = 3'b001;
                width26 = 3'b001;
                width25 = 3'b001;
                width24 = 3'b001;
                width23 = 3'b001;
                width22 = 3'b001;
                width21 = 3'b001;
                width20 = 3'b001;
                width19 = 3'b001;
                width18 = 3'b001;
                width17 = 3'b001;
                width16 = 3'b001;
                width15 = 3'b001;
                width14 = 3'b001;
                width13 = 3'b001;
                width12 = 3'b010;
                width11 = 3'b010;
                width10 = 3'b010;
                width9 = 3'b010;
                width8 = 3'b010;
                width7 = 3'b010;
                width6 = 3'b010;
                width5 = 3'b010;
                width4 = 3'b011;
                width3 = 3'b011;
                width2 = 3'b011;
                width1 = 3'b011;
                width0 = 3'b101;

                writeAddr60 = {writeAddr[13:0]};
                writeAddr59 = {writeAddr[13:0]};
                writeAddr58 = {writeAddr[13:0]};
                writeAddr57 = {writeAddr[13:0]};
                writeAddr56 = {writeAddr[13:0]};
                writeAddr55 = {writeAddr[13:0]};
                writeAddr54 = {writeAddr[13:0]};
                writeAddr53 = {writeAddr[13:0]};
                writeAddr52 = {writeAddr[13:0]};
                writeAddr51 = {writeAddr[13:0]};
                writeAddr50 = {writeAddr[13:0]};
                writeAddr49 = {writeAddr[13:0]};
                writeAddr48 = {writeAddr[13:0]};
                writeAddr47 = {writeAddr[13:0]};
                writeAddr46 = {writeAddr[13:0]};
                writeAddr45 = {writeAddr[13:0]};
                writeAddr44 = {writeAddr[13:0]};
                writeAddr43 = {writeAddr[13:0]};
                writeAddr42 = {writeAddr[13:0]};
                writeAddr41 = {writeAddr[13:0]};
                writeAddr40 = {writeAddr[13:0]};
                writeAddr39 = {writeAddr[13:0]};
                writeAddr38 = {writeAddr[13:0]};
                writeAddr37 = {writeAddr[13:0]};
                writeAddr36 = {writeAddr[13:0]};
                writeAddr35 = {writeAddr[13:0]};
                writeAddr34 = {writeAddr[13:0]};
                writeAddr33 = {writeAddr[13:0]};
                writeAddr32 = {writeAddr[13:0]};
                writeAddr31 = {writeAddr[13:0]};
                writeAddr30 = {writeAddr[13:0]};
                writeAddr29 = {writeAddr[13:0]};
                writeAddr28 = {writeAddr[12:0], 1'b0};
                writeAddr27 = {writeAddr[12:0], 1'b0};
                writeAddr26 = {writeAddr[12:0], 1'b0};
                writeAddr25 = {writeAddr[12:0], 1'b0};
                writeAddr24 = {writeAddr[12:0], 1'b0};
                writeAddr23 = {writeAddr[12:0], 1'b0};
                writeAddr22 = {writeAddr[12:0], 1'b0};
                writeAddr21 = {writeAddr[12:0], 1'b0};
                writeAddr20 = {writeAddr[12:0], 1'b0};
                writeAddr19 = {writeAddr[12:0], 1'b0};
                writeAddr18 = {writeAddr[12:0], 1'b0};
                writeAddr17 = {writeAddr[12:0], 1'b0};
                writeAddr16 = {writeAddr[12:0], 1'b0};
                writeAddr15 = {writeAddr[12:0], 1'b0};
                writeAddr14 = {writeAddr[12:0], 1'b0};
                writeAddr13 = {writeAddr[12:0], 1'b0};
                writeAddr12 = {writeAddr[11:0], 2'b0};
                writeAddr11 = {writeAddr[11:0], 2'b0};
                writeAddr10 = {writeAddr[11:0], 2'b0};
                writeAddr9 = {writeAddr[11:0], 2'b0};
                writeAddr8 = {writeAddr[11:0], 2'b0};
                writeAddr7 = {writeAddr[11:0], 2'b0};
                writeAddr6 = {writeAddr[11:0], 2'b0};
                writeAddr5 = {writeAddr[11:0], 2'b0};
                writeAddr4 = {writeAddr[10:0], 3'b0};
                writeAddr3 = {writeAddr[10:0], 3'b0};
                writeAddr2 = {writeAddr[10:0], 3'b0};
                writeAddr1 = {writeAddr[10:0], 3'b0};
                writeAddr0 = {writeAddr[8:0], 5'b0};

                readAddr60 = {writeAddr[13:0]};
                readAddr59 = {writeAddr[13:0]};
                readAddr58 = {writeAddr[13:0]};
                readAddr57 = {writeAddr[13:0]};
                readAddr56 = {writeAddr[13:0]};
                readAddr55 = {writeAddr[13:0]};
                readAddr54 = {writeAddr[13:0]};
                readAddr53 = {writeAddr[13:0]};
                readAddr52 = {writeAddr[13:0]};
                readAddr51 = {writeAddr[13:0]};
                readAddr50 = {writeAddr[13:0]};
                readAddr49 = {writeAddr[13:0]};
                readAddr48 = {writeAddr[13:0]};
                readAddr47 = {writeAddr[13:0]};
                readAddr46 = {writeAddr[13:0]};
                readAddr45 = {writeAddr[13:0]};
                readAddr44 = {writeAddr[13:0]};
                readAddr43 = {writeAddr[13:0]};
                readAddr42 = {writeAddr[13:0]};
                readAddr41 = {writeAddr[13:0]};
                readAddr40 = {writeAddr[13:0]};
                readAddr39 = {writeAddr[13:0]};
                readAddr38 = {writeAddr[13:0]};
                readAddr37 = {writeAddr[13:0]};
                readAddr36 = {writeAddr[13:0]};
                readAddr35 = {writeAddr[13:0]};
                readAddr34 = {writeAddr[13:0]};
                readAddr33 = {writeAddr[13:0]};
                readAddr32 = {writeAddr[13:0]};
                readAddr31 = {writeAddr[13:0]};
                readAddr30 = {writeAddr[13:0]};
                readAddr29 = {writeAddr[13:0]};
                readAddr28  = {readAddr[12:0],  1'b0};
                readAddr27  = {readAddr[12:0],  1'b0};
                readAddr26  = {readAddr[12:0],  1'b0};
                readAddr25  = {readAddr[12:0],  1'b0};
                readAddr24  = {readAddr[12:0],  1'b0};
                readAddr23  = {readAddr[12:0],  1'b0};
                readAddr22  = {readAddr[12:0],  1'b0};
                readAddr21  = {readAddr[12:0],  1'b0};
                readAddr20  = {readAddr[12:0],  1'b0};
                readAddr19  = {readAddr[12:0],  1'b0};
                readAddr18  = {readAddr[12:0],  1'b0};
                readAddr17  = {readAddr[12:0],  1'b0};
                readAddr16  = {readAddr[12:0],  1'b0};
                readAddr15  = {readAddr[12:0],  1'b0};
                readAddr14  = {readAddr[12:0],  1'b0};
                readAddr13  = {readAddr[12:0],  1'b0};
                readAddr12  = {readAddr[11:0],  2'b0};
                readAddr11  = {readAddr[11:0],  2'b0};
                readAddr10  = {readAddr[11:0],  2'b0};
                readAddr9  = {readAddr[11:0],  2'b0};
                readAddr8  = {readAddr[11:0],  2'b0};
                readAddr7  = {readAddr[11:0],  2'b0};
                readAddr6  = {readAddr[11:0],  2'b0};
                readAddr5  = {readAddr[11:0],  2'b0};
                readAddr4  = {readAddr[10:0],  3'b0};
                readAddr3  = {readAddr[10:0],  3'b0};
                readAddr2  = {readAddr[10:0],  3'b0};
                readAddr1  = {readAddr[10:0],  3'b0};
                readAddr0  = {readAddr[8:0],  5'b0};

                writeData60 = {17'b0, writeData[31]};
                writeData59 = {17'b0, writeData[30]};
                writeData58 = {17'b0, writeData[29]};
                writeData57 = {17'b0, writeData[28]};
                writeData56 = {17'b0, writeData[27]};
                writeData55 = {17'b0, writeData[26]};
                writeData54 = {17'b0, writeData[25]};
                writeData53 = {17'b0, writeData[24]};
                writeData52 = {17'b0, writeData[23]};
                writeData51 = {17'b0, writeData[22]};
                writeData50 = {17'b0, writeData[21]};
                writeData49 = {17'b0, writeData[20]};
                writeData48 = {17'b0, writeData[19]};
                writeData47 = {17'b0, writeData[18]};
                writeData46 = {17'b0, writeData[17]};
                writeData45 = {17'b0, writeData[16]};
                writeData44 = {17'b0, writeData[15]};
                writeData43 = {17'b0, writeData[14]};
                writeData42 = {17'b0, writeData[13]};
                writeData41 = {17'b0, writeData[12]};
                writeData40 = {17'b0, writeData[11]};
                writeData39 = {17'b0, writeData[10]};
                writeData38 = {17'b0, writeData[9]};
                writeData37 = {17'b0, writeData[8]};
                writeData36 = {17'b0, writeData[7]};
                writeData35 = {17'b0, writeData[6]};
                writeData34 = {17'b0, writeData[5]};
                writeData33 = {17'b0, writeData[4]};
                writeData32 = {17'b0, writeData[3]};
                writeData31 = {17'b0, writeData[2]};
                writeData30 = {17'b0, writeData[1]};
                writeData29 = {17'b0, writeData[0]};
                writeData28 = {16'b0, writeData[31:30]};
                writeData27 = {16'b0, writeData[29:28]};
                writeData26 = {16'b0, writeData[27:26]};
                writeData25 = {16'b0, writeData[25:24]};
                writeData24 = {16'b0, writeData[23:22]};
                writeData23 = {16'b0, writeData[21:20]};
                writeData22 = {16'b0, writeData[19:18]};
                writeData21 = {16'b0, writeData[17:16]};
                writeData20 = {16'b0, writeData[15:14]};
                writeData19 = {16'b0, writeData[13:12]};
                writeData18 = {16'b0, writeData[11:10]};
                writeData17 = {16'b0, writeData[9:8]};
                writeData16 = {16'b0, writeData[7:6]};
                writeData15 = {16'b0, writeData[5:4]};
                writeData14 = {16'b0, writeData[3:2]};
                writeData13 = {16'b0, writeData[1:0]};
                writeData12 = {14'b0, writeData[31:28]};
                writeData11 = {14'b0, writeData[27:24]};
                writeData10 = {14'b0, writeData[23:20]};
                writeData9 = {14'b0, writeData[19:16]};
                writeData8 = {14'b0, writeData[15:12]};
                writeData7 = {14'b0, writeData[11:8]};
                writeData6 = {14'b0, writeData[7:4]};
                writeData5 = {14'b0, writeData[3:0]};
                writeData4 = {10'b0, writeData[31:24]};
                writeData3 = {10'b0, writeData[23:16]};
                writeData2 = {10'b0, writeData[15:8]};
                writeData1 = {10'b0, writeData[7:0]};
                writeData0 = {1'b0, writeData[31:24], 1'b0, writeData[23:16], 1'b0, writeData[15:8], 1'b0, writeData[7:0]};

                case (writeAddr[14:9])
                    6'b000000, 6'b000001, 6'b000010, 6'b000011,
                    6'b000100, 6'b000101, 6'b000110, 6'b000111,
                    6'b001000, 6'b001001, 6'b001010, 6'b001011,
                    6'b001100, 6'b001101, 6'b001110, 6'b001111,
                    6'b010000, 6'b010001, 6'b010010, 6'b010011,
                    6'b010100, 6'b010101, 6'b010110, 6'b010111,
                    6'b011000, 6'b011001, 6'b011010, 6'b011011,
                    6'b011100, 6'b011101, 6'b011110, 6'b011111 : begin
                        wen_a60 = {1'b0, wen};
                        wen_a59 = {1'b0, wen};
                        wen_a58 = {1'b0, wen};
                        wen_a57 = {1'b0, wen};
                        wen_a56 = {1'b0, wen};
                        wen_a55 = {1'b0, wen};
                        wen_a54 = {1'b0, wen};
                        wen_a53 = {1'b0, wen};
                        wen_a52 = {1'b0, wen};
                        wen_a51 = {1'b0, wen};
                        wen_a50 = {1'b0, wen};
                        wen_a49 = {1'b0, wen};
                        wen_a48 = {1'b0, wen};
                        wen_a47 = {1'b0, wen};
                        wen_a46 = {1'b0, wen};
                        wen_a45 = {1'b0, wen};
                        wen_a44 = {1'b0, wen};
                        wen_a43 = {1'b0, wen};
                        wen_a42 = {1'b0, wen};
                        wen_a41 = {1'b0, wen};
                        wen_a40 = {1'b0, wen};
                        wen_a39 = {1'b0, wen};
                        wen_a38 = {1'b0, wen};
                        wen_a37 = {1'b0, wen};
                        wen_a36 = {1'b0, wen};
                        wen_a35 = {1'b0, wen};
                        wen_a34 = {1'b0, wen};
                        wen_a33 = {1'b0, wen};
                        wen_a32 = {1'b0, wen};
                        wen_a31 = {1'b0, wen};
                        wen_a30 = {1'b0, wen};
                        wen_a29 = {1'b0, wen};
                        wen_a28 = {1'b0, 1'b0};
                        wen_a27 = {1'b0, 1'b0};
                        wen_a26 = {1'b0, 1'b0};
                        wen_a25 = {1'b0, 1'b0};
                        wen_a24 = {1'b0, 1'b0};
                        wen_a23 = {1'b0, 1'b0};
                        wen_a22 = {1'b0, 1'b0};
                        wen_a21 = {1'b0, 1'b0};
                        wen_a20 = {1'b0, 1'b0};
                        wen_a19 = {1'b0, 1'b0};
                        wen_a18 = {1'b0, 1'b0};
                        wen_a17 = {1'b0, 1'b0};
                        wen_a16 = {1'b0, 1'b0};
                        wen_a15 = {1'b0, 1'b0};
                        wen_a14 = {1'b0, 1'b0};
                        wen_a13 = {1'b0, 1'b0};
                        wen_a12 = {1'b0, 1'b0};
                        wen_a11 = {1'b0, 1'b0};
                        wen_a10 = {1'b0, 1'b0};
                        wen_a9 = {1'b0, 1'b0};
                        wen_a8 = {1'b0, 1'b0};
                        wen_a7 = {1'b0, 1'b0};
                        wen_a6 = {1'b0, 1'b0};
                        wen_a5 = {1'b0, 1'b0};
                        wen_a4 = {1'b0, 1'b0};
                        wen_a3 = {1'b0, 1'b0};
                        wen_a2 = {1'b0, 1'b0};
                        wen_a1 = {1'b0, 1'b0};
                        wen_a0 = {1'b0, 1'b0};
                        wen_b0 = {1'b0, 1'b0};
                    end
                    6'b100000, 6'b100001, 6'b100010, 6'b100011,
                    6'b100100, 6'b100101, 6'b100110, 6'b100111,
                    6'b101000, 6'b101001, 6'b101010, 6'b101011,
                    6'b101100, 6'b101101, 6'b101110, 6'b101111 : begin
                        wen_a60 = {1'b0, 1'b0};
                        wen_a59 = {1'b0, 1'b0};
                        wen_a58 = {1'b0, 1'b0};
                        wen_a57 = {1'b0, 1'b0};
                        wen_a56 = {1'b0, 1'b0};
                        wen_a55 = {1'b0, 1'b0};
                        wen_a54 = {1'b0, 1'b0};
                        wen_a53 = {1'b0, 1'b0};
                        wen_a52 = {1'b0, 1'b0};
                        wen_a51 = {1'b0, 1'b0};
                        wen_a50 = {1'b0, 1'b0};
                        wen_a49 = {1'b0, 1'b0};
                        wen_a48 = {1'b0, 1'b0};
                        wen_a47 = {1'b0, 1'b0};
                        wen_a46 = {1'b0, 1'b0};
                        wen_a45 = {1'b0, 1'b0};
                        wen_a44 = {1'b0, 1'b0};
                        wen_a43 = {1'b0, 1'b0};
                        wen_a42 = {1'b0, 1'b0};
                        wen_a41 = {1'b0, 1'b0};
                        wen_a40 = {1'b0, 1'b0};
                        wen_a39 = {1'b0, 1'b0};
                        wen_a38 = {1'b0, 1'b0};
                        wen_a37 = {1'b0, 1'b0};
                        wen_a36 = {1'b0, 1'b0};
                        wen_a35 = {1'b0, 1'b0};
                        wen_a34 = {1'b0, 1'b0};
                        wen_a33 = {1'b0, 1'b0};
                        wen_a32 = {1'b0, 1'b0};
                        wen_a31 = {1'b0, 1'b0};
                        wen_a30 = {1'b0, 1'b0};
                        wen_a29 = {1'b0, 1'b0};
                        wen_a28 = {1'b0, wen};
                        wen_a27 = {1'b0, wen};
                        wen_a26 = {1'b0, wen};
                        wen_a25 = {1'b0, wen};
                        wen_a24 = {1'b0, wen};
                        wen_a23 = {1'b0, wen};
                        wen_a22 = {1'b0, wen};
                        wen_a21 = {1'b0, wen};
                        wen_a20 = {1'b0, wen};
                        wen_a19 = {1'b0, wen};
                        wen_a18 = {1'b0, wen};
                        wen_a17 = {1'b0, wen};
                        wen_a16 = {1'b0, wen};
                        wen_a15 = {1'b0, wen};
                        wen_a14 = {1'b0, wen};
                        wen_a13 = {1'b0, wen};
                        wen_a12 = {1'b0, 1'b0};
                        wen_a11 = {1'b0, 1'b0};
                        wen_a10 = {1'b0, 1'b0};
                        wen_a9 = {1'b0, 1'b0};
                        wen_a8 = {1'b0, 1'b0};
                        wen_a7 = {1'b0, 1'b0};
                        wen_a6 = {1'b0, 1'b0};
                        wen_a5 = {1'b0, 1'b0};
                        wen_a4 = {1'b0, 1'b0};
                        wen_a3 = {1'b0, 1'b0};
                        wen_a2 = {1'b0, 1'b0};
                        wen_a1 = {1'b0, 1'b0};
                        wen_a0 = {1'b0, 1'b0};
                        wen_b0 = {1'b0, 1'b0};
                    end
                    6'b110000, 6'b110001, 6'b110010, 6'b110011,
                    6'b110100, 6'b110101, 6'b110110, 6'b110111 : begin
                        wen_a60 = {1'b0, 1'b0};
                        wen_a59 = {1'b0, 1'b0};
                        wen_a58 = {1'b0, 1'b0};
                        wen_a57 = {1'b0, 1'b0};
                        wen_a56 = {1'b0, 1'b0};
                        wen_a55 = {1'b0, 1'b0};
                        wen_a54 = {1'b0, 1'b0};
                        wen_a53 = {1'b0, 1'b0};
                        wen_a52 = {1'b0, 1'b0};
                        wen_a51 = {1'b0, 1'b0};
                        wen_a50 = {1'b0, 1'b0};
                        wen_a49 = {1'b0, 1'b0};
                        wen_a48 = {1'b0, 1'b0};
                        wen_a47 = {1'b0, 1'b0};
                        wen_a46 = {1'b0, 1'b0};
                        wen_a45 = {1'b0, 1'b0};
                        wen_a44 = {1'b0, 1'b0};
                        wen_a43 = {1'b0, 1'b0};
                        wen_a42 = {1'b0, 1'b0};
                        wen_a41 = {1'b0, 1'b0};
                        wen_a40 = {1'b0, 1'b0};
                        wen_a39 = {1'b0, 1'b0};
                        wen_a38 = {1'b0, 1'b0};
                        wen_a37 = {1'b0, 1'b0};
                        wen_a36 = {1'b0, 1'b0};
                        wen_a35 = {1'b0, 1'b0};
                        wen_a34 = {1'b0, 1'b0};
                        wen_a33 = {1'b0, 1'b0};
                        wen_a32 = {1'b0, 1'b0};
                        wen_a31 = {1'b0, 1'b0};
                        wen_a30 = {1'b0, 1'b0};
                        wen_a29 = {1'b0, 1'b0};
                        wen_a28 = {1'b0, 1'b0};
                        wen_a27 = {1'b0, 1'b0};
                        wen_a26 = {1'b0, 1'b0};
                        wen_a25 = {1'b0, 1'b0};
                        wen_a24 = {1'b0, 1'b0};
                        wen_a23 = {1'b0, 1'b0};
                        wen_a22 = {1'b0, 1'b0};
                        wen_a21 = {1'b0, 1'b0};
                        wen_a20 = {1'b0, 1'b0};
                        wen_a19 = {1'b0, 1'b0};
                        wen_a18 = {1'b0, 1'b0};
                        wen_a17 = {1'b0, 1'b0};
                        wen_a16 = {1'b0, 1'b0};
                        wen_a15 = {1'b0, 1'b0};
                        wen_a14 = {1'b0, 1'b0};
                        wen_a13 = {1'b0, 1'b0};
                        wen_a12 = {1'b0, wen};
                        wen_a11 = {1'b0, wen};
                        wen_a10 = {1'b0, wen};
                        wen_a9 = {1'b0, wen};
                        wen_a8 = {1'b0, wen};
                        wen_a7 = {1'b0, wen};
                        wen_a6 = {1'b0, wen};
                        wen_a5 = {1'b0, wen};
                        wen_a4 = {1'b0, 1'b0};
                        wen_a3 = {1'b0, 1'b0};
                        wen_a2 = {1'b0, 1'b0};
                        wen_a1 = {1'b0, 1'b0};
                        wen_a0 = {1'b0, 1'b0};
                        wen_b0 = {1'b0, 1'b0};
                    end
                    6'b111000, 6'b111001, 6'b111010, 6'b111011 : begin
                        wen_a60 = {1'b0, 1'b0};
                        wen_a59 = {1'b0, 1'b0};
                        wen_a58 = {1'b0, 1'b0};
                        wen_a57 = {1'b0, 1'b0};
                        wen_a56 = {1'b0, 1'b0};
                        wen_a55 = {1'b0, 1'b0};
                        wen_a54 = {1'b0, 1'b0};
                        wen_a53 = {1'b0, 1'b0};
                        wen_a52 = {1'b0, 1'b0};
                        wen_a51 = {1'b0, 1'b0};
                        wen_a50 = {1'b0, 1'b0};
                        wen_a49 = {1'b0, 1'b0};
                        wen_a48 = {1'b0, 1'b0};
                        wen_a47 = {1'b0, 1'b0};
                        wen_a46 = {1'b0, 1'b0};
                        wen_a45 = {1'b0, 1'b0};
                        wen_a44 = {1'b0, 1'b0};
                        wen_a43 = {1'b0, 1'b0};
                        wen_a42 = {1'b0, 1'b0};
                        wen_a41 = {1'b0, 1'b0};
                        wen_a40 = {1'b0, 1'b0};
                        wen_a39 = {1'b0, 1'b0};
                        wen_a38 = {1'b0, 1'b0};
                        wen_a37 = {1'b0, 1'b0};
                        wen_a36 = {1'b0, 1'b0};
                        wen_a35 = {1'b0, 1'b0};
                        wen_a34 = {1'b0, 1'b0};
                        wen_a33 = {1'b0, 1'b0};
                        wen_a32 = {1'b0, 1'b0};
                        wen_a31 = {1'b0, 1'b0};
                        wen_a30 = {1'b0, 1'b0};
                        wen_a29 = {1'b0, 1'b0};
                        wen_a28 = {1'b0, 1'b0};
                        wen_a27 = {1'b0, 1'b0};
                        wen_a26 = {1'b0, 1'b0};
                        wen_a25 = {1'b0, 1'b0};
                        wen_a24 = {1'b0, 1'b0};
                        wen_a23 = {1'b0, 1'b0};
                        wen_a22 = {1'b0, 1'b0};
                        wen_a21 = {1'b0, 1'b0};
                        wen_a20 = {1'b0, 1'b0};
                        wen_a19 = {1'b0, 1'b0};
                        wen_a18 = {1'b0, 1'b0};
                        wen_a17 = {1'b0, 1'b0};
                        wen_a16 = {1'b0, 1'b0};
                        wen_a15 = {1'b0, 1'b0};
                        wen_a14 = {1'b0, 1'b0};
                        wen_a13 = {1'b0, 1'b0};
                        wen_a12 = {1'b0, 1'b0};
                        wen_a11 = {1'b0, 1'b0};
                        wen_a10 = {1'b0, 1'b0};
                        wen_a9 = {1'b0, 1'b0};
                        wen_a8 = {1'b0, 1'b0};
                        wen_a7 = {1'b0, 1'b0};
                        wen_a6 = {1'b0, 1'b0};
                        wen_a5 = {1'b0, 1'b0};
                        wen_a4 = {1'b0, wen};
                        wen_a3 = {1'b0, wen};
                        wen_a2 = {1'b0, wen};
                        wen_a1 = {1'b0, wen};
                        wen_a0 = {1'b0, 1'b0};
                        wen_b0 = {1'b0, 1'b0};
                    end
                    6'b111100 : begin
                        wen_a60 = {1'b0, 1'b0};
                        wen_a59 = {1'b0, 1'b0};
                        wen_a58 = {1'b0, 1'b0};
                        wen_a57 = {1'b0, 1'b0};
                        wen_a56 = {1'b0, 1'b0};
                        wen_a55 = {1'b0, 1'b0};
                        wen_a54 = {1'b0, 1'b0};
                        wen_a53 = {1'b0, 1'b0};
                        wen_a52 = {1'b0, 1'b0};
                        wen_a51 = {1'b0, 1'b0};
                        wen_a50 = {1'b0, 1'b0};
                        wen_a49 = {1'b0, 1'b0};
                        wen_a48 = {1'b0, 1'b0};
                        wen_a47 = {1'b0, 1'b0};
                        wen_a46 = {1'b0, 1'b0};
                        wen_a45 = {1'b0, 1'b0};
                        wen_a44 = {1'b0, 1'b0};
                        wen_a43 = {1'b0, 1'b0};
                        wen_a42 = {1'b0, 1'b0};
                        wen_a41 = {1'b0, 1'b0};
                        wen_a40 = {1'b0, 1'b0};
                        wen_a39 = {1'b0, 1'b0};
                        wen_a38 = {1'b0, 1'b0};
                        wen_a37 = {1'b0, 1'b0};
                        wen_a36 = {1'b0, 1'b0};
                        wen_a35 = {1'b0, 1'b0};
                        wen_a34 = {1'b0, 1'b0};
                        wen_a33 = {1'b0, 1'b0};
                        wen_a32 = {1'b0, 1'b0};
                        wen_a31 = {1'b0, 1'b0};
                        wen_a30 = {1'b0, 1'b0};
                        wen_a29 = {1'b0, 1'b0};
                        wen_a28 = {1'b0, 1'b0};
                        wen_a27 = {1'b0, 1'b0};
                        wen_a26 = {1'b0, 1'b0};
                        wen_a25 = {1'b0, 1'b0};
                        wen_a24 = {1'b0, 1'b0};
                        wen_a23 = {1'b0, 1'b0};
                        wen_a22 = {1'b0, 1'b0};
                        wen_a21 = {1'b0, 1'b0};
                        wen_a20 = {1'b0, 1'b0};
                        wen_a19 = {1'b0, 1'b0};
                        wen_a18 = {1'b0, 1'b0};
                        wen_a17 = {1'b0, 1'b0};
                        wen_a16 = {1'b0, 1'b0};
                        wen_a15 = {1'b0, 1'b0};
                        wen_a14 = {1'b0, 1'b0};
                        wen_a13 = {1'b0, 1'b0};
                        wen_a12 = {1'b0, 1'b0};
                        wen_a11 = {1'b0, 1'b0};
                        wen_a10 = {1'b0, 1'b0};
                        wen_a9 = {1'b0, 1'b0};
                        wen_a8 = {1'b0, 1'b0};
                        wen_a7 = {1'b0, 1'b0};
                        wen_a6 = {1'b0, 1'b0};
                        wen_a5 = {1'b0, 1'b0};
                        wen_a4 = {1'b0, 1'b0};
                        wen_a3 = {1'b0, 1'b0};
                        wen_a2 = {1'b0, 1'b0};
                        wen_a1 = {1'b0, 1'b0};
                        wen_a0 = {wen, wen};
                        wen_b0 = {wen, wen};
                    end
                    default : begin
                        wen_a60 = {1'b0, 1'b0};
                        wen_a59 = {1'b0, 1'b0};
                        wen_a58 = {1'b0, 1'b0};
                        wen_a57 = {1'b0, 1'b0};
                        wen_a56 = {1'b0, 1'b0};
                        wen_a55 = {1'b0, 1'b0};
                        wen_a54 = {1'b0, 1'b0};
                        wen_a53 = {1'b0, 1'b0};
                        wen_a52 = {1'b0, 1'b0};
                        wen_a51 = {1'b0, 1'b0};
                        wen_a50 = {1'b0, 1'b0};
                        wen_a49 = {1'b0, 1'b0};
                        wen_a48 = {1'b0, 1'b0};
                        wen_a47 = {1'b0, 1'b0};
                        wen_a46 = {1'b0, 1'b0};
                        wen_a45 = {1'b0, 1'b0};
                        wen_a44 = {1'b0, 1'b0};
                        wen_a43 = {1'b0, 1'b0};
                        wen_a42 = {1'b0, 1'b0};
                        wen_a41 = {1'b0, 1'b0};
                        wen_a40 = {1'b0, 1'b0};
                        wen_a39 = {1'b0, 1'b0};
                        wen_a38 = {1'b0, 1'b0};
                        wen_a37 = {1'b0, 1'b0};
                        wen_a36 = {1'b0, 1'b0};
                        wen_a35 = {1'b0, 1'b0};
                        wen_a34 = {1'b0, 1'b0};
                        wen_a33 = {1'b0, 1'b0};
                        wen_a32 = {1'b0, 1'b0};
                        wen_a31 = {1'b0, 1'b0};
                        wen_a30 = {1'b0, 1'b0};
                        wen_a29 = {1'b0, 1'b0};
                        wen_a28 = {1'b0, 1'b0};
                        wen_a27 = {1'b0, 1'b0};
                        wen_a26 = {1'b0, 1'b0};
                        wen_a25 = {1'b0, 1'b0};
                        wen_a24 = {1'b0, 1'b0};
                        wen_a23 = {1'b0, 1'b0};
                        wen_a22 = {1'b0, 1'b0};
                        wen_a21 = {1'b0, 1'b0};
                        wen_a20 = {1'b0, 1'b0};
                        wen_a19 = {1'b0, 1'b0};
                        wen_a18 = {1'b0, 1'b0};
                        wen_a17 = {1'b0, 1'b0};
                        wen_a16 = {1'b0, 1'b0};
                        wen_a15 = {1'b0, 1'b0};
                        wen_a14 = {1'b0, 1'b0};
                        wen_a13 = {1'b0, 1'b0};
                        wen_a12 = {1'b0, 1'b0};
                        wen_a11 = {1'b0, 1'b0};
                        wen_a10 = {1'b0, 1'b0};
                        wen_a9 = {1'b0, 1'b0};
                        wen_a8 = {1'b0, 1'b0};
                        wen_a7 = {1'b0, 1'b0};
                        wen_a6 = {1'b0, 1'b0};
                        wen_a5 = {1'b0, 1'b0};
                        wen_a4 = {1'b0, 1'b0};
                        wen_a3 = {1'b0, 1'b0};
                        wen_a2 = {1'b0, 1'b0};
                        wen_a1 = {1'b0, 1'b0};
                        wen_a0 = {1'b0, 1'b0};
                        wen_b0 = {1'b0, 1'b0};
                    end
                endcase

                case (ckRdAddr[14:9])
                    6'b000000, 6'b000001, 6'b000010, 6'b000011,
                    6'b000100, 6'b000101, 6'b000110, 6'b000111,
                    6'b001000, 6'b001001, 6'b001010, 6'b001011,
                    6'b001100, 6'b001101, 6'b001110, 6'b001111,
                    6'b010000, 6'b010001, 6'b010010, 6'b010011,
                    6'b010100, 6'b010101, 6'b010110, 6'b010111,
                    6'b011000, 6'b011001, 6'b011010, 6'b011011,
                    6'b011100, 6'b011101, 6'b011110, 6'b011111 : begin
                        readData = {
                                        readData60[0],
                                        readData59[0],
                                        readData58[0],
                                        readData57[0],
                                        readData56[0],
                                        readData55[0],
                                        readData54[0],
                                        readData53[0],
                                        readData52[0],
                                        readData51[0],
                                        readData50[0],
                                        readData49[0],
                                        readData48[0],
                                        readData47[0],
                                        readData46[0],
                                        readData45[0],
                                        readData44[0],
                                        readData43[0],
                                        readData42[0],
                                        readData41[0],
                                        readData40[0],
                                        readData39[0],
                                        readData38[0],
                                        readData37[0],
                                        readData36[0],
                                        readData35[0],
                                        readData34[0],
                                        readData33[0],
                                        readData32[0],
                                        readData31[0],
                                        readData30[0],
                                        readData29[0]
                        };
                    end
                    6'b100000, 6'b100001, 6'b100010, 6'b100011,
                    6'b100100, 6'b100101, 6'b100110, 6'b100111,
                    6'b101000, 6'b101001, 6'b101010, 6'b101011,
                    6'b101100, 6'b101101, 6'b101110, 6'b101111 : begin
                        readData = {
                                        readData28[1:0],
                                        readData27[1:0],
                                        readData26[1:0],
                                        readData25[1:0],
                                        readData24[1:0],
                                        readData23[1:0],
                                        readData22[1:0],
                                        readData21[1:0],
                                        readData20[1:0],
                                        readData19[1:0],
                                        readData18[1:0],
                                        readData17[1:0],
                                        readData16[1:0],
                                        readData15[1:0],
                                        readData14[1:0],
                                        readData13[1:0]
                        };
                    end
                    6'b110000, 6'b110001, 6'b110010, 6'b110011,
                    6'b110100, 6'b110101, 6'b110110, 6'b110111 : begin
                        readData = {
                                        readData12[3:0],
                                        readData11[3:0],
                                        readData10[3:0],
                                        readData9[3:0],
                                        readData8[3:0],
                                        readData7[3:0],
                                        readData6[3:0],
                                        readData5[3:0]
                        };
                    end
                    6'b111000, 6'b111001, 6'b111010, 6'b111011 : begin
                        readData = {readData4[7:0],readData3[7:0],readData2[7:0],readData1[7:0]};
                    end
                    6'b111100 : begin
                        readData = {readData0[34:27],readData0[25:18],readData0[16:9],readData0[7:0]};
                    end
                    default : begin
                        readData = 32'b0;
                    end
                endcase
            end        
            31744: begin
                width62 = 3'b000;
                width61 = 3'b000;
                width60 = 3'b000;
                width59 = 3'b000;
                width58 = 3'b000;
                width57 = 3'b000;
                width56 = 3'b000;
                width55 = 3'b000;
                width54 = 3'b000;
                width53 = 3'b000;
                width52 = 3'b000;
                width51 = 3'b000;
                width50 = 3'b000;
                width49 = 3'b000;
                width48 = 3'b000;
                width47 = 3'b000;
                width46 = 3'b000;
                width45 = 3'b000;
                width44 = 3'b000;
                width43 = 3'b000;
                width42 = 3'b000;
                width41 = 3'b000;
                width40 = 3'b000;
                width39 = 3'b000;
                width38 = 3'b000;
                width37 = 3'b000;
                width36 = 3'b000;
                width35 = 3'b000;
                width34 = 3'b000;
                width33 = 3'b000;
                width32 = 3'b000;
                width31 = 3'b000;
                width30 = 3'b001;
                width29 = 3'b001;
                width28 = 3'b001;
                width27 = 3'b001;
                width26 = 3'b001;
                width25 = 3'b001;
                width24 = 3'b001;
                width23 = 3'b001;
                width22 = 3'b001;
                width21 = 3'b001;
                width20 = 3'b001;
                width19 = 3'b001;
                width18 = 3'b001;
                width17 = 3'b001;
                width16 = 3'b001;
                width15 = 3'b001;
                width14 = 3'b010;
                width13 = 3'b010;
                width12 = 3'b010;
                width11 = 3'b010;
                width10 = 3'b010;
                width9 = 3'b010;
                width8 = 3'b010;
                width7 = 3'b010;
                width6 = 3'b011;
                width5 = 3'b011;
                width4 = 3'b011;
                width3 = 3'b011;
                width2 = 3'b100;
                width1 = 3'b100;

                writeAddr62 = {writeAddr[13:0]};
                writeAddr61 = {writeAddr[13:0]};
                writeAddr60 = {writeAddr[13:0]};
                writeAddr59 = {writeAddr[13:0]};
                writeAddr58 = {writeAddr[13:0]};
                writeAddr57 = {writeAddr[13:0]};
                writeAddr56 = {writeAddr[13:0]};
                writeAddr55 = {writeAddr[13:0]};
                writeAddr54 = {writeAddr[13:0]};
                writeAddr53 = {writeAddr[13:0]};
                writeAddr52 = {writeAddr[13:0]};
                writeAddr51 = {writeAddr[13:0]};
                writeAddr50 = {writeAddr[13:0]};
                writeAddr49 = {writeAddr[13:0]};
                writeAddr48 = {writeAddr[13:0]};
                writeAddr47 = {writeAddr[13:0]};
                writeAddr46 = {writeAddr[13:0]};
                writeAddr45 = {writeAddr[13:0]};
                writeAddr44 = {writeAddr[13:0]};
                writeAddr43 = {writeAddr[13:0]};
                writeAddr42 = {writeAddr[13:0]};
                writeAddr41 = {writeAddr[13:0]};
                writeAddr40 = {writeAddr[13:0]};
                writeAddr39 = {writeAddr[13:0]};
                writeAddr38 = {writeAddr[13:0]};
                writeAddr37 = {writeAddr[13:0]};
                writeAddr36 = {writeAddr[13:0]};
                writeAddr35 = {writeAddr[13:0]};
                writeAddr34 = {writeAddr[13:0]};
                writeAddr33 = {writeAddr[13:0]};
                writeAddr32 = {writeAddr[13:0]};
                writeAddr31 = {writeAddr[13:0]};
                writeAddr30 = {writeAddr[12:0], 1'b0};
                writeAddr29 = {writeAddr[12:0], 1'b0};
                writeAddr28 = {writeAddr[12:0], 1'b0};
                writeAddr27 = {writeAddr[12:0], 1'b0};
                writeAddr26 = {writeAddr[12:0], 1'b0};
                writeAddr25 = {writeAddr[12:0], 1'b0};
                writeAddr24 = {writeAddr[12:0], 1'b0};
                writeAddr23 = {writeAddr[12:0], 1'b0};
                writeAddr22 = {writeAddr[12:0], 1'b0};
                writeAddr21 = {writeAddr[12:0], 1'b0};
                writeAddr20 = {writeAddr[12:0], 1'b0};
                writeAddr19 = {writeAddr[12:0], 1'b0};
                writeAddr18 = {writeAddr[12:0], 1'b0};
                writeAddr17 = {writeAddr[12:0], 1'b0};
                writeAddr16 = {writeAddr[12:0], 1'b0};
                writeAddr15 = {writeAddr[12:0], 1'b0};
                writeAddr14 = {writeAddr[11:0], 2'b0};
                writeAddr13 = {writeAddr[11:0], 2'b0};
                writeAddr12 = {writeAddr[11:0], 2'b0};
                writeAddr11 = {writeAddr[11:0], 2'b0};
                writeAddr10 = {writeAddr[11:0], 2'b0};
                writeAddr9 = {writeAddr[11:0], 2'b0};
                writeAddr8 = {writeAddr[11:0], 2'b0};
                writeAddr7 = {writeAddr[11:0], 2'b0};
                writeAddr6 = {writeAddr[10:0], 3'b0};
                writeAddr5 = {writeAddr[10:0], 3'b0};
                writeAddr4 = {writeAddr[10:0], 3'b0};
                writeAddr3 = {writeAddr[10:0], 3'b0};
                writeAddr2 = {writeAddr[9:0], 4'b0};
                writeAddr1 = {writeAddr[9:0], 4'b0};

                readAddr62 = {writeAddr[13:0]};
                readAddr61 = {writeAddr[13:0]};
                readAddr60 = {writeAddr[13:0]};
                readAddr59 = {writeAddr[13:0]};
                readAddr58 = {writeAddr[13:0]};
                readAddr57 = {writeAddr[13:0]};
                readAddr56 = {writeAddr[13:0]};
                readAddr55 = {writeAddr[13:0]};
                readAddr54 = {writeAddr[13:0]};
                readAddr53 = {writeAddr[13:0]};
                readAddr52 = {writeAddr[13:0]};
                readAddr51 = {writeAddr[13:0]};
                readAddr50 = {writeAddr[13:0]};
                readAddr49 = {writeAddr[13:0]};
                readAddr48 = {writeAddr[13:0]};
                readAddr47 = {writeAddr[13:0]};
                readAddr46 = {writeAddr[13:0]};
                readAddr45 = {writeAddr[13:0]};
                readAddr44 = {writeAddr[13:0]};
                readAddr43 = {writeAddr[13:0]};
                readAddr42 = {writeAddr[13:0]};
                readAddr41 = {writeAddr[13:0]};
                readAddr40 = {writeAddr[13:0]};
                readAddr39 = {writeAddr[13:0]};
                readAddr38 = {writeAddr[13:0]};
                readAddr37 = {writeAddr[13:0]};
                readAddr36 = {writeAddr[13:0]};
                readAddr35 = {writeAddr[13:0]};
                readAddr34 = {writeAddr[13:0]};
                readAddr33 = {writeAddr[13:0]};
                readAddr32 = {writeAddr[13:0]};
                readAddr31 = {writeAddr[13:0]};
                readAddr30  = {readAddr[12:0],  1'b0};
                readAddr29  = {readAddr[12:0],  1'b0};
                readAddr28  = {readAddr[12:0],  1'b0};
                readAddr27  = {readAddr[12:0],  1'b0};
                readAddr26  = {readAddr[12:0],  1'b0};
                readAddr25  = {readAddr[12:0],  1'b0};
                readAddr24  = {readAddr[12:0],  1'b0};
                readAddr23  = {readAddr[12:0],  1'b0};
                readAddr22  = {readAddr[12:0],  1'b0};
                readAddr21  = {readAddr[12:0],  1'b0};
                readAddr20  = {readAddr[12:0],  1'b0};
                readAddr19  = {readAddr[12:0],  1'b0};
                readAddr18  = {readAddr[12:0],  1'b0};
                readAddr17  = {readAddr[12:0],  1'b0};
                readAddr16  = {readAddr[12:0],  1'b0};
                readAddr15  = {readAddr[12:0],  1'b0};
                readAddr14  = {readAddr[11:0],  2'b0};
                readAddr13  = {readAddr[11:0],  2'b0};
                readAddr12  = {readAddr[11:0],  2'b0};
                readAddr11  = {readAddr[11:0],  2'b0};
                readAddr10  = {readAddr[11:0],  2'b0};
                readAddr9  = {readAddr[11:0],  2'b0};
                readAddr8  = {readAddr[11:0],  2'b0};
                readAddr7  = {readAddr[11:0],  2'b0};
                readAddr6  = {readAddr[10:0],  3'b0};
                readAddr5  = {readAddr[10:0],  3'b0};
                readAddr4  = {readAddr[10:0],  3'b0};
                readAddr3  = {readAddr[10:0],  3'b0};
                readAddr2  = {readAddr[9:0],  4'b0};
                readAddr1  = {readAddr[9:0],  4'b0};

                writeData62 = {17'b0, writeData[31]};
                writeData61 = {17'b0, writeData[30]};
                writeData60 = {17'b0, writeData[29]};
                writeData59 = {17'b0, writeData[28]};
                writeData58 = {17'b0, writeData[27]};
                writeData57 = {17'b0, writeData[26]};
                writeData56 = {17'b0, writeData[25]};
                writeData55 = {17'b0, writeData[24]};
                writeData54 = {17'b0, writeData[23]};
                writeData53 = {17'b0, writeData[22]};
                writeData52 = {17'b0, writeData[21]};
                writeData51 = {17'b0, writeData[20]};
                writeData50 = {17'b0, writeData[19]};
                writeData49 = {17'b0, writeData[18]};
                writeData48 = {17'b0, writeData[17]};
                writeData47 = {17'b0, writeData[16]};
                writeData46 = {17'b0, writeData[15]};
                writeData45 = {17'b0, writeData[14]};
                writeData44 = {17'b0, writeData[13]};
                writeData43 = {17'b0, writeData[12]};
                writeData42 = {17'b0, writeData[11]};
                writeData41 = {17'b0, writeData[10]};
                writeData40 = {17'b0, writeData[9]};
                writeData39 = {17'b0, writeData[8]};
                writeData38 = {17'b0, writeData[7]};
                writeData37 = {17'b0, writeData[6]};
                writeData36 = {17'b0, writeData[5]};
                writeData35 = {17'b0, writeData[4]};
                writeData34 = {17'b0, writeData[3]};
                writeData33 = {17'b0, writeData[2]};
                writeData32 = {17'b0, writeData[1]};
                writeData31 = {17'b0, writeData[0]};
                writeData30 = {16'b0, writeData[31:30]};
                writeData29 = {16'b0, writeData[29:28]};
                writeData28 = {16'b0, writeData[27:26]};
                writeData27 = {16'b0, writeData[25:24]};
                writeData26 = {16'b0, writeData[23:22]};
                writeData25 = {16'b0, writeData[21:20]};
                writeData24 = {16'b0, writeData[19:18]};
                writeData23 = {16'b0, writeData[17:16]};
                writeData22 = {16'b0, writeData[15:14]};
                writeData21 = {16'b0, writeData[13:12]};
                writeData20 = {16'b0, writeData[11:10]};
                writeData19 = {16'b0, writeData[9:8]};
                writeData18 = {16'b0, writeData[7:6]};
                writeData17 = {16'b0, writeData[5:4]};
                writeData16 = {16'b0, writeData[3:2]};
                writeData15 = {16'b0, writeData[1:0]};
                writeData14 = {14'b0, writeData[31:28]};
                writeData13 = {14'b0, writeData[27:24]};
                writeData12 = {14'b0, writeData[23:20]};
                writeData11 = {14'b0, writeData[19:16]};
                writeData10 = {14'b0, writeData[15:12]};
                writeData9 = {14'b0, writeData[11:8]};
                writeData8 = {14'b0, writeData[7:4]};
                writeData7 = {14'b0, writeData[3:0]};
                writeData6 = {10'b0, writeData[31:24]};
                writeData5 = {10'b0, writeData[23:16]};
                writeData4 = {10'b0, writeData[15:8]};
                writeData3 = {10'b0, writeData[7:0]};
                writeData2 = {1'b0, writeData[31:24], 1'b0, writeData[23:16]};
                writeData1 = {1'b0, writeData[15:8], 1'b0, writeData[7:0]};

                case (writeAddr[14:9])
                    6'b000000, 6'b000001, 6'b000010, 6'b000011,
                    6'b000100, 6'b000101, 6'b000110, 6'b000111,
                    6'b001000, 6'b001001, 6'b001010, 6'b001011,
                    6'b001100, 6'b001101, 6'b001110, 6'b001111,
                    6'b010000, 6'b010001, 6'b010010, 6'b010011,
                    6'b010100, 6'b010101, 6'b010110, 6'b010111,
                    6'b011000, 6'b011001, 6'b011010, 6'b011011,
                    6'b011100, 6'b011101, 6'b011110, 6'b011111 : begin
                        wen_a62 = {1'b0, wen};
                        wen_a61 = {1'b0, wen};
                        wen_a60 = {1'b0, wen};
                        wen_a59 = {1'b0, wen};
                        wen_a58 = {1'b0, wen};
                        wen_a57 = {1'b0, wen};
                        wen_a56 = {1'b0, wen};
                        wen_a55 = {1'b0, wen};
                        wen_a54 = {1'b0, wen};
                        wen_a53 = {1'b0, wen};
                        wen_a52 = {1'b0, wen};
                        wen_a51 = {1'b0, wen};
                        wen_a50 = {1'b0, wen};
                        wen_a49 = {1'b0, wen};
                        wen_a48 = {1'b0, wen};
                        wen_a47 = {1'b0, wen};
                        wen_a46 = {1'b0, wen};
                        wen_a45 = {1'b0, wen};
                        wen_a44 = {1'b0, wen};
                        wen_a43 = {1'b0, wen};
                        wen_a42 = {1'b0, wen};
                        wen_a41 = {1'b0, wen};
                        wen_a40 = {1'b0, wen};
                        wen_a39 = {1'b0, wen};
                        wen_a38 = {1'b0, wen};
                        wen_a37 = {1'b0, wen};
                        wen_a36 = {1'b0, wen};
                        wen_a35 = {1'b0, wen};
                        wen_a34 = {1'b0, wen};
                        wen_a33 = {1'b0, wen};
                        wen_a32 = {1'b0, wen};
                        wen_a31 = {1'b0, wen};
                        wen_a30 = {1'b0, 1'b0};
                        wen_a29 = {1'b0, 1'b0};
                        wen_a28 = {1'b0, 1'b0};
                        wen_a27 = {1'b0, 1'b0};
                        wen_a26 = {1'b0, 1'b0};
                        wen_a25 = {1'b0, 1'b0};
                        wen_a24 = {1'b0, 1'b0};
                        wen_a23 = {1'b0, 1'b0};
                        wen_a22 = {1'b0, 1'b0};
                        wen_a21 = {1'b0, 1'b0};
                        wen_a20 = {1'b0, 1'b0};
                        wen_a19 = {1'b0, 1'b0};
                        wen_a18 = {1'b0, 1'b0};
                        wen_a17 = {1'b0, 1'b0};
                        wen_a16 = {1'b0, 1'b0};
                        wen_a15 = {1'b0, 1'b0};
                        wen_a14 = {1'b0, 1'b0};
                        wen_a13 = {1'b0, 1'b0};
                        wen_a12 = {1'b0, 1'b0};
                        wen_a11 = {1'b0, 1'b0};
                        wen_a10 = {1'b0, 1'b0};
                        wen_a9 = {1'b0, 1'b0};
                        wen_a8 = {1'b0, 1'b0};
                        wen_a7 = {1'b0, 1'b0};
                        wen_a6 = {1'b0, 1'b0};
                        wen_a5 = {1'b0, 1'b0};
                        wen_a4 = {1'b0, 1'b0};
                        wen_a3 = {1'b0, 1'b0};
                        wen_a2 = {1'b0, 1'b0};
                        wen_a1 = {1'b0, 1'b0};
                    end
                    6'b100000, 6'b100001, 6'b100010, 6'b100011,
                    6'b100100, 6'b100101, 6'b100110, 6'b100111,
                    6'b101000, 6'b101001, 6'b101010, 6'b101011,
                    6'b101100, 6'b101101, 6'b101110, 6'b101111 : begin
                        wen_a62 = {1'b0, 1'b0};
                        wen_a61 = {1'b0, 1'b0};
                        wen_a60 = {1'b0, 1'b0};
                        wen_a59 = {1'b0, 1'b0};
                        wen_a58 = {1'b0, 1'b0};
                        wen_a57 = {1'b0, 1'b0};
                        wen_a56 = {1'b0, 1'b0};
                        wen_a55 = {1'b0, 1'b0};
                        wen_a54 = {1'b0, 1'b0};
                        wen_a53 = {1'b0, 1'b0};
                        wen_a52 = {1'b0, 1'b0};
                        wen_a51 = {1'b0, 1'b0};
                        wen_a50 = {1'b0, 1'b0};
                        wen_a49 = {1'b0, 1'b0};
                        wen_a48 = {1'b0, 1'b0};
                        wen_a47 = {1'b0, 1'b0};
                        wen_a46 = {1'b0, 1'b0};
                        wen_a45 = {1'b0, 1'b0};
                        wen_a44 = {1'b0, 1'b0};
                        wen_a43 = {1'b0, 1'b0};
                        wen_a42 = {1'b0, 1'b0};
                        wen_a41 = {1'b0, 1'b0};
                        wen_a40 = {1'b0, 1'b0};
                        wen_a39 = {1'b0, 1'b0};
                        wen_a38 = {1'b0, 1'b0};
                        wen_a37 = {1'b0, 1'b0};
                        wen_a36 = {1'b0, 1'b0};
                        wen_a35 = {1'b0, 1'b0};
                        wen_a34 = {1'b0, 1'b0};
                        wen_a33 = {1'b0, 1'b0};
                        wen_a32 = {1'b0, 1'b0};
                        wen_a31 = {1'b0, 1'b0};
                        wen_a30 = {1'b0, wen};
                        wen_a29 = {1'b0, wen};
                        wen_a28 = {1'b0, wen};
                        wen_a27 = {1'b0, wen};
                        wen_a26 = {1'b0, wen};
                        wen_a25 = {1'b0, wen};
                        wen_a24 = {1'b0, wen};
                        wen_a23 = {1'b0, wen};
                        wen_a22 = {1'b0, wen};
                        wen_a21 = {1'b0, wen};
                        wen_a20 = {1'b0, wen};
                        wen_a19 = {1'b0, wen};
                        wen_a18 = {1'b0, wen};
                        wen_a17 = {1'b0, wen};
                        wen_a16 = {1'b0, wen};
                        wen_a15 = {1'b0, wen};
                        wen_a14 = {1'b0, 1'b0};
                        wen_a13 = {1'b0, 1'b0};
                        wen_a12 = {1'b0, 1'b0};
                        wen_a11 = {1'b0, 1'b0};
                        wen_a10 = {1'b0, 1'b0};
                        wen_a9 = {1'b0, 1'b0};
                        wen_a8 = {1'b0, 1'b0};
                        wen_a7 = {1'b0, 1'b0};
                        wen_a6 = {1'b0, 1'b0};
                        wen_a5 = {1'b0, 1'b0};
                        wen_a4 = {1'b0, 1'b0};
                        wen_a3 = {1'b0, 1'b0};
                        wen_a2 = {1'b0, 1'b0};
                        wen_a1 = {1'b0, 1'b0};
                    end
                    6'b110000, 6'b110001, 6'b110010, 6'b110011,
                    6'b110100, 6'b110101, 6'b110110, 6'b110111 : begin
                        wen_a62 = {1'b0, 1'b0};
                        wen_a61 = {1'b0, 1'b0};
                        wen_a60 = {1'b0, 1'b0};
                        wen_a59 = {1'b0, 1'b0};
                        wen_a58 = {1'b0, 1'b0};
                        wen_a57 = {1'b0, 1'b0};
                        wen_a56 = {1'b0, 1'b0};
                        wen_a55 = {1'b0, 1'b0};
                        wen_a54 = {1'b0, 1'b0};
                        wen_a53 = {1'b0, 1'b0};
                        wen_a52 = {1'b0, 1'b0};
                        wen_a51 = {1'b0, 1'b0};
                        wen_a50 = {1'b0, 1'b0};
                        wen_a49 = {1'b0, 1'b0};
                        wen_a48 = {1'b0, 1'b0};
                        wen_a47 = {1'b0, 1'b0};
                        wen_a46 = {1'b0, 1'b0};
                        wen_a45 = {1'b0, 1'b0};
                        wen_a44 = {1'b0, 1'b0};
                        wen_a43 = {1'b0, 1'b0};
                        wen_a42 = {1'b0, 1'b0};
                        wen_a41 = {1'b0, 1'b0};
                        wen_a40 = {1'b0, 1'b0};
                        wen_a39 = {1'b0, 1'b0};
                        wen_a38 = {1'b0, 1'b0};
                        wen_a37 = {1'b0, 1'b0};
                        wen_a36 = {1'b0, 1'b0};
                        wen_a35 = {1'b0, 1'b0};
                        wen_a34 = {1'b0, 1'b0};
                        wen_a33 = {1'b0, 1'b0};
                        wen_a32 = {1'b0, 1'b0};
                        wen_a31 = {1'b0, 1'b0};
                        wen_a30 = {1'b0, 1'b0};
                        wen_a29 = {1'b0, 1'b0};
                        wen_a28 = {1'b0, 1'b0};
                        wen_a27 = {1'b0, 1'b0};
                        wen_a26 = {1'b0, 1'b0};
                        wen_a25 = {1'b0, 1'b0};
                        wen_a24 = {1'b0, 1'b0};
                        wen_a23 = {1'b0, 1'b0};
                        wen_a22 = {1'b0, 1'b0};
                        wen_a21 = {1'b0, 1'b0};
                        wen_a20 = {1'b0, 1'b0};
                        wen_a19 = {1'b0, 1'b0};
                        wen_a18 = {1'b0, 1'b0};
                        wen_a17 = {1'b0, 1'b0};
                        wen_a16 = {1'b0, 1'b0};
                        wen_a15 = {1'b0, 1'b0};
                        wen_a14 = {1'b0, wen};
                        wen_a13 = {1'b0, wen};
                        wen_a12 = {1'b0, wen};
                        wen_a11 = {1'b0, wen};
                        wen_a10 = {1'b0, wen};
                        wen_a9 = {1'b0, wen};
                        wen_a8 = {1'b0, wen};
                        wen_a7 = {1'b0, wen};
                        wen_a6 = {1'b0, 1'b0};
                        wen_a5 = {1'b0, 1'b0};
                        wen_a4 = {1'b0, 1'b0};
                        wen_a3 = {1'b0, 1'b0};
                        wen_a2 = {1'b0, 1'b0};
                        wen_a1 = {1'b0, 1'b0};
                    end
                    6'b111000, 6'b111001, 6'b111010, 6'b111011 : begin
                        wen_a62 = {1'b0, 1'b0};
                        wen_a61 = {1'b0, 1'b0};
                        wen_a60 = {1'b0, 1'b0};
                        wen_a59 = {1'b0, 1'b0};
                        wen_a58 = {1'b0, 1'b0};
                        wen_a57 = {1'b0, 1'b0};
                        wen_a56 = {1'b0, 1'b0};
                        wen_a55 = {1'b0, 1'b0};
                        wen_a54 = {1'b0, 1'b0};
                        wen_a53 = {1'b0, 1'b0};
                        wen_a52 = {1'b0, 1'b0};
                        wen_a51 = {1'b0, 1'b0};
                        wen_a50 = {1'b0, 1'b0};
                        wen_a49 = {1'b0, 1'b0};
                        wen_a48 = {1'b0, 1'b0};
                        wen_a47 = {1'b0, 1'b0};
                        wen_a46 = {1'b0, 1'b0};
                        wen_a45 = {1'b0, 1'b0};
                        wen_a44 = {1'b0, 1'b0};
                        wen_a43 = {1'b0, 1'b0};
                        wen_a42 = {1'b0, 1'b0};
                        wen_a41 = {1'b0, 1'b0};
                        wen_a40 = {1'b0, 1'b0};
                        wen_a39 = {1'b0, 1'b0};
                        wen_a38 = {1'b0, 1'b0};
                        wen_a37 = {1'b0, 1'b0};
                        wen_a36 = {1'b0, 1'b0};
                        wen_a35 = {1'b0, 1'b0};
                        wen_a34 = {1'b0, 1'b0};
                        wen_a33 = {1'b0, 1'b0};
                        wen_a32 = {1'b0, 1'b0};
                        wen_a31 = {1'b0, 1'b0};
                        wen_a30 = {1'b0, 1'b0};
                        wen_a29 = {1'b0, 1'b0};
                        wen_a28 = {1'b0, 1'b0};
                        wen_a27 = {1'b0, 1'b0};
                        wen_a26 = {1'b0, 1'b0};
                        wen_a25 = {1'b0, 1'b0};
                        wen_a24 = {1'b0, 1'b0};
                        wen_a23 = {1'b0, 1'b0};
                        wen_a22 = {1'b0, 1'b0};
                        wen_a21 = {1'b0, 1'b0};
                        wen_a20 = {1'b0, 1'b0};
                        wen_a19 = {1'b0, 1'b0};
                        wen_a18 = {1'b0, 1'b0};
                        wen_a17 = {1'b0, 1'b0};
                        wen_a16 = {1'b0, 1'b0};
                        wen_a15 = {1'b0, 1'b0};
                        wen_a14 = {1'b0, 1'b0};
                        wen_a13 = {1'b0, 1'b0};
                        wen_a12 = {1'b0, 1'b0};
                        wen_a11 = {1'b0, 1'b0};
                        wen_a10 = {1'b0, 1'b0};
                        wen_a9 = {1'b0, 1'b0};
                        wen_a8 = {1'b0, 1'b0};
                        wen_a7 = {1'b0, 1'b0};
                        wen_a6 = {1'b0, wen};
                        wen_a5 = {1'b0, wen};
                        wen_a4 = {1'b0, wen};
                        wen_a3 = {1'b0, wen};
                        wen_a2 = {1'b0, 1'b0};
                        wen_a1 = {1'b0, 1'b0};
                    end
                    6'b111100, 6'b111101 : begin
                        wen_a62 = {1'b0, 1'b0};
                        wen_a61 = {1'b0, 1'b0};
                        wen_a60 = {1'b0, 1'b0};
                        wen_a59 = {1'b0, 1'b0};
                        wen_a58 = {1'b0, 1'b0};
                        wen_a57 = {1'b0, 1'b0};
                        wen_a56 = {1'b0, 1'b0};
                        wen_a55 = {1'b0, 1'b0};
                        wen_a54 = {1'b0, 1'b0};
                        wen_a53 = {1'b0, 1'b0};
                        wen_a52 = {1'b0, 1'b0};
                        wen_a51 = {1'b0, 1'b0};
                        wen_a50 = {1'b0, 1'b0};
                        wen_a49 = {1'b0, 1'b0};
                        wen_a48 = {1'b0, 1'b0};
                        wen_a47 = {1'b0, 1'b0};
                        wen_a46 = {1'b0, 1'b0};
                        wen_a45 = {1'b0, 1'b0};
                        wen_a44 = {1'b0, 1'b0};
                        wen_a43 = {1'b0, 1'b0};
                        wen_a42 = {1'b0, 1'b0};
                        wen_a41 = {1'b0, 1'b0};
                        wen_a40 = {1'b0, 1'b0};
                        wen_a39 = {1'b0, 1'b0};
                        wen_a38 = {1'b0, 1'b0};
                        wen_a37 = {1'b0, 1'b0};
                        wen_a36 = {1'b0, 1'b0};
                        wen_a35 = {1'b0, 1'b0};
                        wen_a34 = {1'b0, 1'b0};
                        wen_a33 = {1'b0, 1'b0};
                        wen_a32 = {1'b0, 1'b0};
                        wen_a31 = {1'b0, 1'b0};
                        wen_a30 = {1'b0, 1'b0};
                        wen_a29 = {1'b0, 1'b0};
                        wen_a28 = {1'b0, 1'b0};
                        wen_a27 = {1'b0, 1'b0};
                        wen_a26 = {1'b0, 1'b0};
                        wen_a25 = {1'b0, 1'b0};
                        wen_a24 = {1'b0, 1'b0};
                        wen_a23 = {1'b0, 1'b0};
                        wen_a22 = {1'b0, 1'b0};
                        wen_a21 = {1'b0, 1'b0};
                        wen_a20 = {1'b0, 1'b0};
                        wen_a19 = {1'b0, 1'b0};
                        wen_a18 = {1'b0, 1'b0};
                        wen_a17 = {1'b0, 1'b0};
                        wen_a16 = {1'b0, 1'b0};
                        wen_a15 = {1'b0, 1'b0};
                        wen_a14 = {1'b0, 1'b0};
                        wen_a13 = {1'b0, 1'b0};
                        wen_a12 = {1'b0, 1'b0};
                        wen_a11 = {1'b0, 1'b0};
                        wen_a10 = {1'b0, 1'b0};
                        wen_a9 = {1'b0, 1'b0};
                        wen_a8 = {1'b0, 1'b0};
                        wen_a7 = {1'b0, 1'b0};
                        wen_a6 = {1'b0, 1'b0};
                        wen_a5 = {1'b0, 1'b0};
                        wen_a4 = {1'b0, 1'b0};
                        wen_a3 = {1'b0, 1'b0};
                        wen_a2 = {wen, wen};
                        wen_a1 = {wen, wen};
                    end
                    default : begin
                        wen_a62 = {1'b0, 1'b0};
                        wen_a61 = {1'b0, 1'b0};
                        wen_a60 = {1'b0, 1'b0};
                        wen_a59 = {1'b0, 1'b0};
                        wen_a58 = {1'b0, 1'b0};
                        wen_a57 = {1'b0, 1'b0};
                        wen_a56 = {1'b0, 1'b0};
                        wen_a55 = {1'b0, 1'b0};
                        wen_a54 = {1'b0, 1'b0};
                        wen_a53 = {1'b0, 1'b0};
                        wen_a52 = {1'b0, 1'b0};
                        wen_a51 = {1'b0, 1'b0};
                        wen_a50 = {1'b0, 1'b0};
                        wen_a49 = {1'b0, 1'b0};
                        wen_a48 = {1'b0, 1'b0};
                        wen_a47 = {1'b0, 1'b0};
                        wen_a46 = {1'b0, 1'b0};
                        wen_a45 = {1'b0, 1'b0};
                        wen_a44 = {1'b0, 1'b0};
                        wen_a43 = {1'b0, 1'b0};
                        wen_a42 = {1'b0, 1'b0};
                        wen_a41 = {1'b0, 1'b0};
                        wen_a40 = {1'b0, 1'b0};
                        wen_a39 = {1'b0, 1'b0};
                        wen_a38 = {1'b0, 1'b0};
                        wen_a37 = {1'b0, 1'b0};
                        wen_a36 = {1'b0, 1'b0};
                        wen_a35 = {1'b0, 1'b0};
                        wen_a34 = {1'b0, 1'b0};
                        wen_a33 = {1'b0, 1'b0};
                        wen_a32 = {1'b0, 1'b0};
                        wen_a31 = {1'b0, 1'b0};
                        wen_a30 = {1'b0, 1'b0};
                        wen_a29 = {1'b0, 1'b0};
                        wen_a28 = {1'b0, 1'b0};
                        wen_a27 = {1'b0, 1'b0};
                        wen_a26 = {1'b0, 1'b0};
                        wen_a25 = {1'b0, 1'b0};
                        wen_a24 = {1'b0, 1'b0};
                        wen_a23 = {1'b0, 1'b0};
                        wen_a22 = {1'b0, 1'b0};
                        wen_a21 = {1'b0, 1'b0};
                        wen_a20 = {1'b0, 1'b0};
                        wen_a19 = {1'b0, 1'b0};
                        wen_a18 = {1'b0, 1'b0};
                        wen_a17 = {1'b0, 1'b0};
                        wen_a16 = {1'b0, 1'b0};
                        wen_a15 = {1'b0, 1'b0};
                        wen_a14 = {1'b0, 1'b0};
                        wen_a13 = {1'b0, 1'b0};
                        wen_a12 = {1'b0, 1'b0};
                        wen_a11 = {1'b0, 1'b0};
                        wen_a10 = {1'b0, 1'b0};
                        wen_a9 = {1'b0, 1'b0};
                        wen_a8 = {1'b0, 1'b0};
                        wen_a7 = {1'b0, 1'b0};
                        wen_a6 = {1'b0, 1'b0};
                        wen_a5 = {1'b0, 1'b0};
                        wen_a4 = {1'b0, 1'b0};
                        wen_a3 = {1'b0, 1'b0};
                        wen_a2 = {1'b0, 1'b0};
                        wen_a1 = {1'b0, 1'b0};
                    end
                endcase

                case (ckRdAddr[14:9])
                    6'b000000, 6'b000001, 6'b000010, 6'b000011,
                    6'b000100, 6'b000101, 6'b000110, 6'b000111,
                    6'b001000, 6'b001001, 6'b001010, 6'b001011,
                    6'b001100, 6'b001101, 6'b001110, 6'b001111,
                    6'b010000, 6'b010001, 6'b010010, 6'b010011,
                    6'b010100, 6'b010101, 6'b010110, 6'b010111,
                    6'b011000, 6'b011001, 6'b011010, 6'b011011,
                    6'b011100, 6'b011101, 6'b011110, 6'b011111 : begin
                        readData = {
                                        readData62[0],
                                        readData61[0],
                                        readData60[0],
                                        readData59[0],
                                        readData58[0],
                                        readData57[0],
                                        readData56[0],
                                        readData55[0],
                                        readData54[0],
                                        readData53[0],
                                        readData52[0],
                                        readData51[0],
                                        readData50[0],
                                        readData49[0],
                                        readData48[0],
                                        readData47[0],
                                        readData46[0],
                                        readData45[0],
                                        readData44[0],
                                        readData43[0],
                                        readData42[0],
                                        readData41[0],
                                        readData40[0],
                                        readData39[0],
                                        readData38[0],
                                        readData37[0],
                                        readData36[0],
                                        readData35[0],
                                        readData34[0],
                                        readData33[0],
                                        readData32[0],
                                        readData31[0]
                        };
                    end
                    6'b100000, 6'b100001, 6'b100010, 6'b100011,
                    6'b100100, 6'b100101, 6'b100110, 6'b100111,
                    6'b101000, 6'b101001, 6'b101010, 6'b101011,
                    6'b101100, 6'b101101, 6'b101110, 6'b101111 : begin
                        readData = {
                                        readData30[1:0],
                                        readData29[1:0],
                                        readData28[1:0],
                                        readData27[1:0],
                                        readData26[1:0],
                                        readData25[1:0],
                                        readData24[1:0],
                                        readData23[1:0],
                                        readData22[1:0],
                                        readData21[1:0],
                                        readData20[1:0],
                                        readData19[1:0],
                                        readData18[1:0],
                                        readData17[1:0],
                                        readData16[1:0],
                                        readData15[1:0]
                        };
                    end
                    6'b110000, 6'b110001, 6'b110010, 6'b110011,
                    6'b110100, 6'b110101, 6'b110110, 6'b110111 : begin
                        readData = {
                                        readData14[3:0],
                                        readData13[3:0],
                                        readData12[3:0],
                                        readData11[3:0],
                                        readData10[3:0],
                                        readData9[3:0],
                                        readData8[3:0],
                                        readData7[3:0]
                        };
                    end
                    6'b111000, 6'b111001, 6'b111010, 6'b111011 : begin
                        readData = {readData6[7:0],readData5[7:0],readData4[7:0],readData3[7:0]};
                    end
                    6'b111100, 6'b111101 : begin
                        readData = {readData2[16:9],readData2[7:0],readData1[16:9],readData1[7:0]};
                    end
                    default : begin
                        readData = 32'b0;
                    end
                endcase
            end        
            32256: begin
                width62 = 3'b000;
                width61 = 3'b000;
                width60 = 3'b000;
                width59 = 3'b000;
                width58 = 3'b000;
                width57 = 3'b000;
                width56 = 3'b000;
                width55 = 3'b000;
                width54 = 3'b000;
                width53 = 3'b000;
                width52 = 3'b000;
                width51 = 3'b000;
                width50 = 3'b000;
                width49 = 3'b000;
                width48 = 3'b000;
                width47 = 3'b000;
                width46 = 3'b000;
                width45 = 3'b000;
                width44 = 3'b000;
                width43 = 3'b000;
                width42 = 3'b000;
                width41 = 3'b000;
                width40 = 3'b000;
                width39 = 3'b000;
                width38 = 3'b000;
                width37 = 3'b000;
                width36 = 3'b000;
                width35 = 3'b000;
                width34 = 3'b000;
                width33 = 3'b000;
                width32 = 3'b000;
                width31 = 3'b000;
                width30 = 3'b001;
                width29 = 3'b001;
                width28 = 3'b001;
                width27 = 3'b001;
                width26 = 3'b001;
                width25 = 3'b001;
                width24 = 3'b001;
                width23 = 3'b001;
                width22 = 3'b001;
                width21 = 3'b001;
                width20 = 3'b001;
                width19 = 3'b001;
                width18 = 3'b001;
                width17 = 3'b001;
                width16 = 3'b001;
                width15 = 3'b001;
                width14 = 3'b010;
                width13 = 3'b010;
                width12 = 3'b010;
                width11 = 3'b010;
                width10 = 3'b010;
                width9 = 3'b010;
                width8 = 3'b010;
                width7 = 3'b010;
                width6 = 3'b011;
                width5 = 3'b011;
                width4 = 3'b011;
                width3 = 3'b011;
                width2 = 3'b100;
                width1 = 3'b100;
                width0 = 3'b101;

                writeAddr62 = {writeAddr[13:0]};
                writeAddr61 = {writeAddr[13:0]};
                writeAddr60 = {writeAddr[13:0]};
                writeAddr59 = {writeAddr[13:0]};
                writeAddr58 = {writeAddr[13:0]};
                writeAddr57 = {writeAddr[13:0]};
                writeAddr56 = {writeAddr[13:0]};
                writeAddr55 = {writeAddr[13:0]};
                writeAddr54 = {writeAddr[13:0]};
                writeAddr53 = {writeAddr[13:0]};
                writeAddr52 = {writeAddr[13:0]};
                writeAddr51 = {writeAddr[13:0]};
                writeAddr50 = {writeAddr[13:0]};
                writeAddr49 = {writeAddr[13:0]};
                writeAddr48 = {writeAddr[13:0]};
                writeAddr47 = {writeAddr[13:0]};
                writeAddr46 = {writeAddr[13:0]};
                writeAddr45 = {writeAddr[13:0]};
                writeAddr44 = {writeAddr[13:0]};
                writeAddr43 = {writeAddr[13:0]};
                writeAddr42 = {writeAddr[13:0]};
                writeAddr41 = {writeAddr[13:0]};
                writeAddr40 = {writeAddr[13:0]};
                writeAddr39 = {writeAddr[13:0]};
                writeAddr38 = {writeAddr[13:0]};
                writeAddr37 = {writeAddr[13:0]};
                writeAddr36 = {writeAddr[13:0]};
                writeAddr35 = {writeAddr[13:0]};
                writeAddr34 = {writeAddr[13:0]};
                writeAddr33 = {writeAddr[13:0]};
                writeAddr32 = {writeAddr[13:0]};
                writeAddr31 = {writeAddr[13:0]};
                writeAddr30 = {writeAddr[12:0], 1'b0};
                writeAddr29 = {writeAddr[12:0], 1'b0};
                writeAddr28 = {writeAddr[12:0], 1'b0};
                writeAddr27 = {writeAddr[12:0], 1'b0};
                writeAddr26 = {writeAddr[12:0], 1'b0};
                writeAddr25 = {writeAddr[12:0], 1'b0};
                writeAddr24 = {writeAddr[12:0], 1'b0};
                writeAddr23 = {writeAddr[12:0], 1'b0};
                writeAddr22 = {writeAddr[12:0], 1'b0};
                writeAddr21 = {writeAddr[12:0], 1'b0};
                writeAddr20 = {writeAddr[12:0], 1'b0};
                writeAddr19 = {writeAddr[12:0], 1'b0};
                writeAddr18 = {writeAddr[12:0], 1'b0};
                writeAddr17 = {writeAddr[12:0], 1'b0};
                writeAddr16 = {writeAddr[12:0], 1'b0};
                writeAddr15 = {writeAddr[12:0], 1'b0};
                writeAddr14 = {writeAddr[11:0], 2'b0};
                writeAddr13 = {writeAddr[11:0], 2'b0};
                writeAddr12 = {writeAddr[11:0], 2'b0};
                writeAddr11 = {writeAddr[11:0], 2'b0};
                writeAddr10 = {writeAddr[11:0], 2'b0};
                writeAddr9 = {writeAddr[11:0], 2'b0};
                writeAddr8 = {writeAddr[11:0], 2'b0};
                writeAddr7 = {writeAddr[11:0], 2'b0};
                writeAddr6 = {writeAddr[10:0], 3'b0};
                writeAddr5 = {writeAddr[10:0], 3'b0};
                writeAddr4 = {writeAddr[10:0], 3'b0};
                writeAddr3 = {writeAddr[10:0], 3'b0};
                writeAddr2 = {writeAddr[9:0], 4'b0};
                writeAddr1 = {writeAddr[9:0], 4'b0};
                writeAddr0 = {writeAddr[8:0], 5'b0};

                readAddr62 = {writeAddr[13:0]};
                readAddr61 = {writeAddr[13:0]};
                readAddr60 = {writeAddr[13:0]};
                readAddr59 = {writeAddr[13:0]};
                readAddr58 = {writeAddr[13:0]};
                readAddr57 = {writeAddr[13:0]};
                readAddr56 = {writeAddr[13:0]};
                readAddr55 = {writeAddr[13:0]};
                readAddr54 = {writeAddr[13:0]};
                readAddr53 = {writeAddr[13:0]};
                readAddr52 = {writeAddr[13:0]};
                readAddr51 = {writeAddr[13:0]};
                readAddr50 = {writeAddr[13:0]};
                readAddr49 = {writeAddr[13:0]};
                readAddr48 = {writeAddr[13:0]};
                readAddr47 = {writeAddr[13:0]};
                readAddr46 = {writeAddr[13:0]};
                readAddr45 = {writeAddr[13:0]};
                readAddr44 = {writeAddr[13:0]};
                readAddr43 = {writeAddr[13:0]};
                readAddr42 = {writeAddr[13:0]};
                readAddr41 = {writeAddr[13:0]};
                readAddr40 = {writeAddr[13:0]};
                readAddr39 = {writeAddr[13:0]};
                readAddr38 = {writeAddr[13:0]};
                readAddr37 = {writeAddr[13:0]};
                readAddr36 = {writeAddr[13:0]};
                readAddr35 = {writeAddr[13:0]};
                readAddr34 = {writeAddr[13:0]};
                readAddr33 = {writeAddr[13:0]};
                readAddr32 = {writeAddr[13:0]};
                readAddr31 = {writeAddr[13:0]};
                readAddr30  = {readAddr[12:0],  1'b0};
                readAddr29  = {readAddr[12:0],  1'b0};
                readAddr28  = {readAddr[12:0],  1'b0};
                readAddr27  = {readAddr[12:0],  1'b0};
                readAddr26  = {readAddr[12:0],  1'b0};
                readAddr25  = {readAddr[12:0],  1'b0};
                readAddr24  = {readAddr[12:0],  1'b0};
                readAddr23  = {readAddr[12:0],  1'b0};
                readAddr22  = {readAddr[12:0],  1'b0};
                readAddr21  = {readAddr[12:0],  1'b0};
                readAddr20  = {readAddr[12:0],  1'b0};
                readAddr19  = {readAddr[12:0],  1'b0};
                readAddr18  = {readAddr[12:0],  1'b0};
                readAddr17  = {readAddr[12:0],  1'b0};
                readAddr16  = {readAddr[12:0],  1'b0};
                readAddr15  = {readAddr[12:0],  1'b0};
                readAddr14  = {readAddr[11:0],  2'b0};
                readAddr13  = {readAddr[11:0],  2'b0};
                readAddr12  = {readAddr[11:0],  2'b0};
                readAddr11  = {readAddr[11:0],  2'b0};
                readAddr10  = {readAddr[11:0],  2'b0};
                readAddr9  = {readAddr[11:0],  2'b0};
                readAddr8  = {readAddr[11:0],  2'b0};
                readAddr7  = {readAddr[11:0],  2'b0};
                readAddr6  = {readAddr[10:0],  3'b0};
                readAddr5  = {readAddr[10:0],  3'b0};
                readAddr4  = {readAddr[10:0],  3'b0};
                readAddr3  = {readAddr[10:0],  3'b0};
                readAddr2  = {readAddr[9:0],  4'b0};
                readAddr1  = {readAddr[9:0],  4'b0};
                readAddr0  = {readAddr[8:0],  5'b0};

                writeData62 = {17'b0, writeData[31]};
                writeData61 = {17'b0, writeData[30]};
                writeData60 = {17'b0, writeData[29]};
                writeData59 = {17'b0, writeData[28]};
                writeData58 = {17'b0, writeData[27]};
                writeData57 = {17'b0, writeData[26]};
                writeData56 = {17'b0, writeData[25]};
                writeData55 = {17'b0, writeData[24]};
                writeData54 = {17'b0, writeData[23]};
                writeData53 = {17'b0, writeData[22]};
                writeData52 = {17'b0, writeData[21]};
                writeData51 = {17'b0, writeData[20]};
                writeData50 = {17'b0, writeData[19]};
                writeData49 = {17'b0, writeData[18]};
                writeData48 = {17'b0, writeData[17]};
                writeData47 = {17'b0, writeData[16]};
                writeData46 = {17'b0, writeData[15]};
                writeData45 = {17'b0, writeData[14]};
                writeData44 = {17'b0, writeData[13]};
                writeData43 = {17'b0, writeData[12]};
                writeData42 = {17'b0, writeData[11]};
                writeData41 = {17'b0, writeData[10]};
                writeData40 = {17'b0, writeData[9]};
                writeData39 = {17'b0, writeData[8]};
                writeData38 = {17'b0, writeData[7]};
                writeData37 = {17'b0, writeData[6]};
                writeData36 = {17'b0, writeData[5]};
                writeData35 = {17'b0, writeData[4]};
                writeData34 = {17'b0, writeData[3]};
                writeData33 = {17'b0, writeData[2]};
                writeData32 = {17'b0, writeData[1]};
                writeData31 = {17'b0, writeData[0]};
                writeData30 = {16'b0, writeData[31:30]};
                writeData29 = {16'b0, writeData[29:28]};
                writeData28 = {16'b0, writeData[27:26]};
                writeData27 = {16'b0, writeData[25:24]};
                writeData26 = {16'b0, writeData[23:22]};
                writeData25 = {16'b0, writeData[21:20]};
                writeData24 = {16'b0, writeData[19:18]};
                writeData23 = {16'b0, writeData[17:16]};
                writeData22 = {16'b0, writeData[15:14]};
                writeData21 = {16'b0, writeData[13:12]};
                writeData20 = {16'b0, writeData[11:10]};
                writeData19 = {16'b0, writeData[9:8]};
                writeData18 = {16'b0, writeData[7:6]};
                writeData17 = {16'b0, writeData[5:4]};
                writeData16 = {16'b0, writeData[3:2]};
                writeData15 = {16'b0, writeData[1:0]};
                writeData14 = {14'b0, writeData[31:28]};
                writeData13 = {14'b0, writeData[27:24]};
                writeData12 = {14'b0, writeData[23:20]};
                writeData11 = {14'b0, writeData[19:16]};
                writeData10 = {14'b0, writeData[15:12]};
                writeData9 = {14'b0, writeData[11:8]};
                writeData8 = {14'b0, writeData[7:4]};
                writeData7 = {14'b0, writeData[3:0]};
                writeData6 = {10'b0, writeData[31:24]};
                writeData5 = {10'b0, writeData[23:16]};
                writeData4 = {10'b0, writeData[15:8]};
                writeData3 = {10'b0, writeData[7:0]};
                writeData2 = {1'b0, writeData[31:24], 1'b0, writeData[23:16]};
                writeData1 = {1'b0, writeData[15:8], 1'b0, writeData[7:0]};
                writeData0 = {1'b0, writeData[31:24], 1'b0, writeData[23:16], 1'b0, writeData[15:8], 1'b0, writeData[7:0]};

                case (writeAddr[14:9])
                    6'b000000, 6'b000001, 6'b000010, 6'b000011,
                    6'b000100, 6'b000101, 6'b000110, 6'b000111,
                    6'b001000, 6'b001001, 6'b001010, 6'b001011,
                    6'b001100, 6'b001101, 6'b001110, 6'b001111,
                    6'b010000, 6'b010001, 6'b010010, 6'b010011,
                    6'b010100, 6'b010101, 6'b010110, 6'b010111,
                    6'b011000, 6'b011001, 6'b011010, 6'b011011,
                    6'b011100, 6'b011101, 6'b011110, 6'b011111 : begin
                        wen_a62 = {1'b0, wen};
                        wen_a61 = {1'b0, wen};
                        wen_a60 = {1'b0, wen};
                        wen_a59 = {1'b0, wen};
                        wen_a58 = {1'b0, wen};
                        wen_a57 = {1'b0, wen};
                        wen_a56 = {1'b0, wen};
                        wen_a55 = {1'b0, wen};
                        wen_a54 = {1'b0, wen};
                        wen_a53 = {1'b0, wen};
                        wen_a52 = {1'b0, wen};
                        wen_a51 = {1'b0, wen};
                        wen_a50 = {1'b0, wen};
                        wen_a49 = {1'b0, wen};
                        wen_a48 = {1'b0, wen};
                        wen_a47 = {1'b0, wen};
                        wen_a46 = {1'b0, wen};
                        wen_a45 = {1'b0, wen};
                        wen_a44 = {1'b0, wen};
                        wen_a43 = {1'b0, wen};
                        wen_a42 = {1'b0, wen};
                        wen_a41 = {1'b0, wen};
                        wen_a40 = {1'b0, wen};
                        wen_a39 = {1'b0, wen};
                        wen_a38 = {1'b0, wen};
                        wen_a37 = {1'b0, wen};
                        wen_a36 = {1'b0, wen};
                        wen_a35 = {1'b0, wen};
                        wen_a34 = {1'b0, wen};
                        wen_a33 = {1'b0, wen};
                        wen_a32 = {1'b0, wen};
                        wen_a31 = {1'b0, wen};
                        wen_a30 = {1'b0, 1'b0};
                        wen_a29 = {1'b0, 1'b0};
                        wen_a28 = {1'b0, 1'b0};
                        wen_a27 = {1'b0, 1'b0};
                        wen_a26 = {1'b0, 1'b0};
                        wen_a25 = {1'b0, 1'b0};
                        wen_a24 = {1'b0, 1'b0};
                        wen_a23 = {1'b0, 1'b0};
                        wen_a22 = {1'b0, 1'b0};
                        wen_a21 = {1'b0, 1'b0};
                        wen_a20 = {1'b0, 1'b0};
                        wen_a19 = {1'b0, 1'b0};
                        wen_a18 = {1'b0, 1'b0};
                        wen_a17 = {1'b0, 1'b0};
                        wen_a16 = {1'b0, 1'b0};
                        wen_a15 = {1'b0, 1'b0};
                        wen_a14 = {1'b0, 1'b0};
                        wen_a13 = {1'b0, 1'b0};
                        wen_a12 = {1'b0, 1'b0};
                        wen_a11 = {1'b0, 1'b0};
                        wen_a10 = {1'b0, 1'b0};
                        wen_a9 = {1'b0, 1'b0};
                        wen_a8 = {1'b0, 1'b0};
                        wen_a7 = {1'b0, 1'b0};
                        wen_a6 = {1'b0, 1'b0};
                        wen_a5 = {1'b0, 1'b0};
                        wen_a4 = {1'b0, 1'b0};
                        wen_a3 = {1'b0, 1'b0};
                        wen_a2 = {1'b0, 1'b0};
                        wen_a1 = {1'b0, 1'b0};
                        wen_a0 = {1'b0, 1'b0};
                        wen_b0 = {1'b0, 1'b0};
                    end
                    6'b100000, 6'b100001, 6'b100010, 6'b100011,
                    6'b100100, 6'b100101, 6'b100110, 6'b100111,
                    6'b101000, 6'b101001, 6'b101010, 6'b101011,
                    6'b101100, 6'b101101, 6'b101110, 6'b101111 : begin
                        wen_a62 = {1'b0, 1'b0};
                        wen_a61 = {1'b0, 1'b0};
                        wen_a60 = {1'b0, 1'b0};
                        wen_a59 = {1'b0, 1'b0};
                        wen_a58 = {1'b0, 1'b0};
                        wen_a57 = {1'b0, 1'b0};
                        wen_a56 = {1'b0, 1'b0};
                        wen_a55 = {1'b0, 1'b0};
                        wen_a54 = {1'b0, 1'b0};
                        wen_a53 = {1'b0, 1'b0};
                        wen_a52 = {1'b0, 1'b0};
                        wen_a51 = {1'b0, 1'b0};
                        wen_a50 = {1'b0, 1'b0};
                        wen_a49 = {1'b0, 1'b0};
                        wen_a48 = {1'b0, 1'b0};
                        wen_a47 = {1'b0, 1'b0};
                        wen_a46 = {1'b0, 1'b0};
                        wen_a45 = {1'b0, 1'b0};
                        wen_a44 = {1'b0, 1'b0};
                        wen_a43 = {1'b0, 1'b0};
                        wen_a42 = {1'b0, 1'b0};
                        wen_a41 = {1'b0, 1'b0};
                        wen_a40 = {1'b0, 1'b0};
                        wen_a39 = {1'b0, 1'b0};
                        wen_a38 = {1'b0, 1'b0};
                        wen_a37 = {1'b0, 1'b0};
                        wen_a36 = {1'b0, 1'b0};
                        wen_a35 = {1'b0, 1'b0};
                        wen_a34 = {1'b0, 1'b0};
                        wen_a33 = {1'b0, 1'b0};
                        wen_a32 = {1'b0, 1'b0};
                        wen_a31 = {1'b0, 1'b0};
                        wen_a30 = {1'b0, wen};
                        wen_a29 = {1'b0, wen};
                        wen_a28 = {1'b0, wen};
                        wen_a27 = {1'b0, wen};
                        wen_a26 = {1'b0, wen};
                        wen_a25 = {1'b0, wen};
                        wen_a24 = {1'b0, wen};
                        wen_a23 = {1'b0, wen};
                        wen_a22 = {1'b0, wen};
                        wen_a21 = {1'b0, wen};
                        wen_a20 = {1'b0, wen};
                        wen_a19 = {1'b0, wen};
                        wen_a18 = {1'b0, wen};
                        wen_a17 = {1'b0, wen};
                        wen_a16 = {1'b0, wen};
                        wen_a15 = {1'b0, wen};
                        wen_a14 = {1'b0, 1'b0};
                        wen_a13 = {1'b0, 1'b0};
                        wen_a12 = {1'b0, 1'b0};
                        wen_a11 = {1'b0, 1'b0};
                        wen_a10 = {1'b0, 1'b0};
                        wen_a9 = {1'b0, 1'b0};
                        wen_a8 = {1'b0, 1'b0};
                        wen_a7 = {1'b0, 1'b0};
                        wen_a6 = {1'b0, 1'b0};
                        wen_a5 = {1'b0, 1'b0};
                        wen_a4 = {1'b0, 1'b0};
                        wen_a3 = {1'b0, 1'b0};
                        wen_a2 = {1'b0, 1'b0};
                        wen_a1 = {1'b0, 1'b0};
                        wen_a0 = {1'b0, 1'b0};
                        wen_b0 = {1'b0, 1'b0};
                    end
                    6'b110000, 6'b110001, 6'b110010, 6'b110011,
                    6'b110100, 6'b110101, 6'b110110, 6'b110111 : begin
                        wen_a62 = {1'b0, 1'b0};
                        wen_a61 = {1'b0, 1'b0};
                        wen_a60 = {1'b0, 1'b0};
                        wen_a59 = {1'b0, 1'b0};
                        wen_a58 = {1'b0, 1'b0};
                        wen_a57 = {1'b0, 1'b0};
                        wen_a56 = {1'b0, 1'b0};
                        wen_a55 = {1'b0, 1'b0};
                        wen_a54 = {1'b0, 1'b0};
                        wen_a53 = {1'b0, 1'b0};
                        wen_a52 = {1'b0, 1'b0};
                        wen_a51 = {1'b0, 1'b0};
                        wen_a50 = {1'b0, 1'b0};
                        wen_a49 = {1'b0, 1'b0};
                        wen_a48 = {1'b0, 1'b0};
                        wen_a47 = {1'b0, 1'b0};
                        wen_a46 = {1'b0, 1'b0};
                        wen_a45 = {1'b0, 1'b0};
                        wen_a44 = {1'b0, 1'b0};
                        wen_a43 = {1'b0, 1'b0};
                        wen_a42 = {1'b0, 1'b0};
                        wen_a41 = {1'b0, 1'b0};
                        wen_a40 = {1'b0, 1'b0};
                        wen_a39 = {1'b0, 1'b0};
                        wen_a38 = {1'b0, 1'b0};
                        wen_a37 = {1'b0, 1'b0};
                        wen_a36 = {1'b0, 1'b0};
                        wen_a35 = {1'b0, 1'b0};
                        wen_a34 = {1'b0, 1'b0};
                        wen_a33 = {1'b0, 1'b0};
                        wen_a32 = {1'b0, 1'b0};
                        wen_a31 = {1'b0, 1'b0};
                        wen_a30 = {1'b0, 1'b0};
                        wen_a29 = {1'b0, 1'b0};
                        wen_a28 = {1'b0, 1'b0};
                        wen_a27 = {1'b0, 1'b0};
                        wen_a26 = {1'b0, 1'b0};
                        wen_a25 = {1'b0, 1'b0};
                        wen_a24 = {1'b0, 1'b0};
                        wen_a23 = {1'b0, 1'b0};
                        wen_a22 = {1'b0, 1'b0};
                        wen_a21 = {1'b0, 1'b0};
                        wen_a20 = {1'b0, 1'b0};
                        wen_a19 = {1'b0, 1'b0};
                        wen_a18 = {1'b0, 1'b0};
                        wen_a17 = {1'b0, 1'b0};
                        wen_a16 = {1'b0, 1'b0};
                        wen_a15 = {1'b0, 1'b0};
                        wen_a14 = {1'b0, wen};
                        wen_a13 = {1'b0, wen};
                        wen_a12 = {1'b0, wen};
                        wen_a11 = {1'b0, wen};
                        wen_a10 = {1'b0, wen};
                        wen_a9 = {1'b0, wen};
                        wen_a8 = {1'b0, wen};
                        wen_a7 = {1'b0, wen};
                        wen_a6 = {1'b0, 1'b0};
                        wen_a5 = {1'b0, 1'b0};
                        wen_a4 = {1'b0, 1'b0};
                        wen_a3 = {1'b0, 1'b0};
                        wen_a2 = {1'b0, 1'b0};
                        wen_a1 = {1'b0, 1'b0};
                        wen_a0 = {1'b0, 1'b0};
                        wen_b0 = {1'b0, 1'b0};
                    end
                    6'b111000, 6'b111001, 6'b111010, 6'b111011 : begin
                        wen_a62 = {1'b0, 1'b0};
                        wen_a61 = {1'b0, 1'b0};
                        wen_a60 = {1'b0, 1'b0};
                        wen_a59 = {1'b0, 1'b0};
                        wen_a58 = {1'b0, 1'b0};
                        wen_a57 = {1'b0, 1'b0};
                        wen_a56 = {1'b0, 1'b0};
                        wen_a55 = {1'b0, 1'b0};
                        wen_a54 = {1'b0, 1'b0};
                        wen_a53 = {1'b0, 1'b0};
                        wen_a52 = {1'b0, 1'b0};
                        wen_a51 = {1'b0, 1'b0};
                        wen_a50 = {1'b0, 1'b0};
                        wen_a49 = {1'b0, 1'b0};
                        wen_a48 = {1'b0, 1'b0};
                        wen_a47 = {1'b0, 1'b0};
                        wen_a46 = {1'b0, 1'b0};
                        wen_a45 = {1'b0, 1'b0};
                        wen_a44 = {1'b0, 1'b0};
                        wen_a43 = {1'b0, 1'b0};
                        wen_a42 = {1'b0, 1'b0};
                        wen_a41 = {1'b0, 1'b0};
                        wen_a40 = {1'b0, 1'b0};
                        wen_a39 = {1'b0, 1'b0};
                        wen_a38 = {1'b0, 1'b0};
                        wen_a37 = {1'b0, 1'b0};
                        wen_a36 = {1'b0, 1'b0};
                        wen_a35 = {1'b0, 1'b0};
                        wen_a34 = {1'b0, 1'b0};
                        wen_a33 = {1'b0, 1'b0};
                        wen_a32 = {1'b0, 1'b0};
                        wen_a31 = {1'b0, 1'b0};
                        wen_a30 = {1'b0, 1'b0};
                        wen_a29 = {1'b0, 1'b0};
                        wen_a28 = {1'b0, 1'b0};
                        wen_a27 = {1'b0, 1'b0};
                        wen_a26 = {1'b0, 1'b0};
                        wen_a25 = {1'b0, 1'b0};
                        wen_a24 = {1'b0, 1'b0};
                        wen_a23 = {1'b0, 1'b0};
                        wen_a22 = {1'b0, 1'b0};
                        wen_a21 = {1'b0, 1'b0};
                        wen_a20 = {1'b0, 1'b0};
                        wen_a19 = {1'b0, 1'b0};
                        wen_a18 = {1'b0, 1'b0};
                        wen_a17 = {1'b0, 1'b0};
                        wen_a16 = {1'b0, 1'b0};
                        wen_a15 = {1'b0, 1'b0};
                        wen_a14 = {1'b0, 1'b0};
                        wen_a13 = {1'b0, 1'b0};
                        wen_a12 = {1'b0, 1'b0};
                        wen_a11 = {1'b0, 1'b0};
                        wen_a10 = {1'b0, 1'b0};
                        wen_a9 = {1'b0, 1'b0};
                        wen_a8 = {1'b0, 1'b0};
                        wen_a7 = {1'b0, 1'b0};
                        wen_a6 = {1'b0, wen};
                        wen_a5 = {1'b0, wen};
                        wen_a4 = {1'b0, wen};
                        wen_a3 = {1'b0, wen};
                        wen_a2 = {1'b0, 1'b0};
                        wen_a1 = {1'b0, 1'b0};
                        wen_a0 = {1'b0, 1'b0};
                        wen_b0 = {1'b0, 1'b0};
                    end
                    6'b111100, 6'b111101 : begin
                        wen_a62 = {1'b0, 1'b0};
                        wen_a61 = {1'b0, 1'b0};
                        wen_a60 = {1'b0, 1'b0};
                        wen_a59 = {1'b0, 1'b0};
                        wen_a58 = {1'b0, 1'b0};
                        wen_a57 = {1'b0, 1'b0};
                        wen_a56 = {1'b0, 1'b0};
                        wen_a55 = {1'b0, 1'b0};
                        wen_a54 = {1'b0, 1'b0};
                        wen_a53 = {1'b0, 1'b0};
                        wen_a52 = {1'b0, 1'b0};
                        wen_a51 = {1'b0, 1'b0};
                        wen_a50 = {1'b0, 1'b0};
                        wen_a49 = {1'b0, 1'b0};
                        wen_a48 = {1'b0, 1'b0};
                        wen_a47 = {1'b0, 1'b0};
                        wen_a46 = {1'b0, 1'b0};
                        wen_a45 = {1'b0, 1'b0};
                        wen_a44 = {1'b0, 1'b0};
                        wen_a43 = {1'b0, 1'b0};
                        wen_a42 = {1'b0, 1'b0};
                        wen_a41 = {1'b0, 1'b0};
                        wen_a40 = {1'b0, 1'b0};
                        wen_a39 = {1'b0, 1'b0};
                        wen_a38 = {1'b0, 1'b0};
                        wen_a37 = {1'b0, 1'b0};
                        wen_a36 = {1'b0, 1'b0};
                        wen_a35 = {1'b0, 1'b0};
                        wen_a34 = {1'b0, 1'b0};
                        wen_a33 = {1'b0, 1'b0};
                        wen_a32 = {1'b0, 1'b0};
                        wen_a31 = {1'b0, 1'b0};
                        wen_a30 = {1'b0, 1'b0};
                        wen_a29 = {1'b0, 1'b0};
                        wen_a28 = {1'b0, 1'b0};
                        wen_a27 = {1'b0, 1'b0};
                        wen_a26 = {1'b0, 1'b0};
                        wen_a25 = {1'b0, 1'b0};
                        wen_a24 = {1'b0, 1'b0};
                        wen_a23 = {1'b0, 1'b0};
                        wen_a22 = {1'b0, 1'b0};
                        wen_a21 = {1'b0, 1'b0};
                        wen_a20 = {1'b0, 1'b0};
                        wen_a19 = {1'b0, 1'b0};
                        wen_a18 = {1'b0, 1'b0};
                        wen_a17 = {1'b0, 1'b0};
                        wen_a16 = {1'b0, 1'b0};
                        wen_a15 = {1'b0, 1'b0};
                        wen_a14 = {1'b0, 1'b0};
                        wen_a13 = {1'b0, 1'b0};
                        wen_a12 = {1'b0, 1'b0};
                        wen_a11 = {1'b0, 1'b0};
                        wen_a10 = {1'b0, 1'b0};
                        wen_a9 = {1'b0, 1'b0};
                        wen_a8 = {1'b0, 1'b0};
                        wen_a7 = {1'b0, 1'b0};
                        wen_a6 = {1'b0, 1'b0};
                        wen_a5 = {1'b0, 1'b0};
                        wen_a4 = {1'b0, 1'b0};
                        wen_a3 = {1'b0, 1'b0};
                        wen_a2 = {wen, wen};
                        wen_a1 = {wen, wen};
                        wen_a0 = {1'b0, 1'b0};
                        wen_b0 = {1'b0, 1'b0};
                    end
                    6'b111110 : begin
                        wen_a62 = {1'b0, 1'b0};
                        wen_a61 = {1'b0, 1'b0};
                        wen_a60 = {1'b0, 1'b0};
                        wen_a59 = {1'b0, 1'b0};
                        wen_a58 = {1'b0, 1'b0};
                        wen_a57 = {1'b0, 1'b0};
                        wen_a56 = {1'b0, 1'b0};
                        wen_a55 = {1'b0, 1'b0};
                        wen_a54 = {1'b0, 1'b0};
                        wen_a53 = {1'b0, 1'b0};
                        wen_a52 = {1'b0, 1'b0};
                        wen_a51 = {1'b0, 1'b0};
                        wen_a50 = {1'b0, 1'b0};
                        wen_a49 = {1'b0, 1'b0};
                        wen_a48 = {1'b0, 1'b0};
                        wen_a47 = {1'b0, 1'b0};
                        wen_a46 = {1'b0, 1'b0};
                        wen_a45 = {1'b0, 1'b0};
                        wen_a44 = {1'b0, 1'b0};
                        wen_a43 = {1'b0, 1'b0};
                        wen_a42 = {1'b0, 1'b0};
                        wen_a41 = {1'b0, 1'b0};
                        wen_a40 = {1'b0, 1'b0};
                        wen_a39 = {1'b0, 1'b0};
                        wen_a38 = {1'b0, 1'b0};
                        wen_a37 = {1'b0, 1'b0};
                        wen_a36 = {1'b0, 1'b0};
                        wen_a35 = {1'b0, 1'b0};
                        wen_a34 = {1'b0, 1'b0};
                        wen_a33 = {1'b0, 1'b0};
                        wen_a32 = {1'b0, 1'b0};
                        wen_a31 = {1'b0, 1'b0};
                        wen_a30 = {1'b0, 1'b0};
                        wen_a29 = {1'b0, 1'b0};
                        wen_a28 = {1'b0, 1'b0};
                        wen_a27 = {1'b0, 1'b0};
                        wen_a26 = {1'b0, 1'b0};
                        wen_a25 = {1'b0, 1'b0};
                        wen_a24 = {1'b0, 1'b0};
                        wen_a23 = {1'b0, 1'b0};
                        wen_a22 = {1'b0, 1'b0};
                        wen_a21 = {1'b0, 1'b0};
                        wen_a20 = {1'b0, 1'b0};
                        wen_a19 = {1'b0, 1'b0};
                        wen_a18 = {1'b0, 1'b0};
                        wen_a17 = {1'b0, 1'b0};
                        wen_a16 = {1'b0, 1'b0};
                        wen_a15 = {1'b0, 1'b0};
                        wen_a14 = {1'b0, 1'b0};
                        wen_a13 = {1'b0, 1'b0};
                        wen_a12 = {1'b0, 1'b0};
                        wen_a11 = {1'b0, 1'b0};
                        wen_a10 = {1'b0, 1'b0};
                        wen_a9 = {1'b0, 1'b0};
                        wen_a8 = {1'b0, 1'b0};
                        wen_a7 = {1'b0, 1'b0};
                        wen_a6 = {1'b0, 1'b0};
                        wen_a5 = {1'b0, 1'b0};
                        wen_a4 = {1'b0, 1'b0};
                        wen_a3 = {1'b0, 1'b0};
                        wen_a2 = {1'b0, 1'b0};
                        wen_a1 = {1'b0, 1'b0};
                        wen_a0 = {wen, wen};
                        wen_b0 = {wen, wen};
                    end
                    default : begin
                        wen_a62 = {1'b0, 1'b0};
                        wen_a61 = {1'b0, 1'b0};
                        wen_a60 = {1'b0, 1'b0};
                        wen_a59 = {1'b0, 1'b0};
                        wen_a58 = {1'b0, 1'b0};
                        wen_a57 = {1'b0, 1'b0};
                        wen_a56 = {1'b0, 1'b0};
                        wen_a55 = {1'b0, 1'b0};
                        wen_a54 = {1'b0, 1'b0};
                        wen_a53 = {1'b0, 1'b0};
                        wen_a52 = {1'b0, 1'b0};
                        wen_a51 = {1'b0, 1'b0};
                        wen_a50 = {1'b0, 1'b0};
                        wen_a49 = {1'b0, 1'b0};
                        wen_a48 = {1'b0, 1'b0};
                        wen_a47 = {1'b0, 1'b0};
                        wen_a46 = {1'b0, 1'b0};
                        wen_a45 = {1'b0, 1'b0};
                        wen_a44 = {1'b0, 1'b0};
                        wen_a43 = {1'b0, 1'b0};
                        wen_a42 = {1'b0, 1'b0};
                        wen_a41 = {1'b0, 1'b0};
                        wen_a40 = {1'b0, 1'b0};
                        wen_a39 = {1'b0, 1'b0};
                        wen_a38 = {1'b0, 1'b0};
                        wen_a37 = {1'b0, 1'b0};
                        wen_a36 = {1'b0, 1'b0};
                        wen_a35 = {1'b0, 1'b0};
                        wen_a34 = {1'b0, 1'b0};
                        wen_a33 = {1'b0, 1'b0};
                        wen_a32 = {1'b0, 1'b0};
                        wen_a31 = {1'b0, 1'b0};
                        wen_a30 = {1'b0, 1'b0};
                        wen_a29 = {1'b0, 1'b0};
                        wen_a28 = {1'b0, 1'b0};
                        wen_a27 = {1'b0, 1'b0};
                        wen_a26 = {1'b0, 1'b0};
                        wen_a25 = {1'b0, 1'b0};
                        wen_a24 = {1'b0, 1'b0};
                        wen_a23 = {1'b0, 1'b0};
                        wen_a22 = {1'b0, 1'b0};
                        wen_a21 = {1'b0, 1'b0};
                        wen_a20 = {1'b0, 1'b0};
                        wen_a19 = {1'b0, 1'b0};
                        wen_a18 = {1'b0, 1'b0};
                        wen_a17 = {1'b0, 1'b0};
                        wen_a16 = {1'b0, 1'b0};
                        wen_a15 = {1'b0, 1'b0};
                        wen_a14 = {1'b0, 1'b0};
                        wen_a13 = {1'b0, 1'b0};
                        wen_a12 = {1'b0, 1'b0};
                        wen_a11 = {1'b0, 1'b0};
                        wen_a10 = {1'b0, 1'b0};
                        wen_a9 = {1'b0, 1'b0};
                        wen_a8 = {1'b0, 1'b0};
                        wen_a7 = {1'b0, 1'b0};
                        wen_a6 = {1'b0, 1'b0};
                        wen_a5 = {1'b0, 1'b0};
                        wen_a4 = {1'b0, 1'b0};
                        wen_a3 = {1'b0, 1'b0};
                        wen_a2 = {1'b0, 1'b0};
                        wen_a1 = {1'b0, 1'b0};
                        wen_a0 = {1'b0, 1'b0};
                        wen_b0 = {1'b0, 1'b0};
                    end
                endcase

                case (ckRdAddr[14:9])
                    6'b000000, 6'b000001, 6'b000010, 6'b000011,
                    6'b000100, 6'b000101, 6'b000110, 6'b000111,
                    6'b001000, 6'b001001, 6'b001010, 6'b001011,
                    6'b001100, 6'b001101, 6'b001110, 6'b001111,
                    6'b010000, 6'b010001, 6'b010010, 6'b010011,
                    6'b010100, 6'b010101, 6'b010110, 6'b010111,
                    6'b011000, 6'b011001, 6'b011010, 6'b011011,
                    6'b011100, 6'b011101, 6'b011110, 6'b011111 : begin
                        readData = {
                                        readData62[0],
                                        readData61[0],
                                        readData60[0],
                                        readData59[0],
                                        readData58[0],
                                        readData57[0],
                                        readData56[0],
                                        readData55[0],
                                        readData54[0],
                                        readData53[0],
                                        readData52[0],
                                        readData51[0],
                                        readData50[0],
                                        readData49[0],
                                        readData48[0],
                                        readData47[0],
                                        readData46[0],
                                        readData45[0],
                                        readData44[0],
                                        readData43[0],
                                        readData42[0],
                                        readData41[0],
                                        readData40[0],
                                        readData39[0],
                                        readData38[0],
                                        readData37[0],
                                        readData36[0],
                                        readData35[0],
                                        readData34[0],
                                        readData33[0],
                                        readData32[0],
                                        readData31[0]
                        };
                    end
                    6'b100000, 6'b100001, 6'b100010, 6'b100011,
                    6'b100100, 6'b100101, 6'b100110, 6'b100111,
                    6'b101000, 6'b101001, 6'b101010, 6'b101011,
                    6'b101100, 6'b101101, 6'b101110, 6'b101111 : begin
                        readData = {
                                        readData30[1:0],
                                        readData29[1:0],
                                        readData28[1:0],
                                        readData27[1:0],
                                        readData26[1:0],
                                        readData25[1:0],
                                        readData24[1:0],
                                        readData23[1:0],
                                        readData22[1:0],
                                        readData21[1:0],
                                        readData20[1:0],
                                        readData19[1:0],
                                        readData18[1:0],
                                        readData17[1:0],
                                        readData16[1:0],
                                        readData15[1:0]
                        };
                    end
                    6'b110000, 6'b110001, 6'b110010, 6'b110011,
                    6'b110100, 6'b110101, 6'b110110, 6'b110111 : begin
                        readData = {
                                        readData14[3:0],
                                        readData13[3:0],
                                        readData12[3:0],
                                        readData11[3:0],
                                        readData10[3:0],
                                        readData9[3:0],
                                        readData8[3:0],
                                        readData7[3:0]
                        };
                    end
                    6'b111000, 6'b111001, 6'b111010, 6'b111011 : begin
                        readData = {readData6[7:0],readData5[7:0],readData4[7:0],readData3[7:0]};
                    end
                    6'b111100, 6'b111101 : begin
                        readData = {readData2[16:9],readData2[7:0],readData1[16:9],readData1[7:0]};
                    end
                    6'b111110 : begin
                        readData = {readData0[34:27],readData0[25:18],readData0[16:9],readData0[7:0]};
                    end
                    default : begin
                        readData = 32'b0;
                    end
                endcase
            end        
            32768: begin
                width64 = 3'b000;
                width63 = 3'b000;
                width62 = 3'b000;
                width61 = 3'b000;
                width60 = 3'b000;
                width59 = 3'b000;
                width58 = 3'b000;
                width57 = 3'b000;
                width56 = 3'b000;
                width55 = 3'b000;
                width54 = 3'b000;
                width53 = 3'b000;
                width52 = 3'b000;
                width51 = 3'b000;
                width50 = 3'b000;
                width49 = 3'b000;
                width48 = 3'b000;
                width47 = 3'b000;
                width46 = 3'b000;
                width45 = 3'b000;
                width44 = 3'b000;
                width43 = 3'b000;
                width42 = 3'b000;
                width41 = 3'b000;
                width40 = 3'b000;
                width39 = 3'b000;
                width38 = 3'b000;
                width37 = 3'b000;
                width36 = 3'b000;
                width35 = 3'b000;
                width34 = 3'b000;
                width33 = 3'b000;
                width32 = 3'b000;
                width31 = 3'b000;
                width30 = 3'b000;
                width29 = 3'b000;
                width28 = 3'b000;
                width27 = 3'b000;
                width26 = 3'b000;
                width25 = 3'b000;
                width24 = 3'b000;
                width23 = 3'b000;
                width22 = 3'b000;
                width21 = 3'b000;
                width20 = 3'b000;
                width19 = 3'b000;
                width18 = 3'b000;
                width17 = 3'b000;
                width16 = 3'b000;
                width15 = 3'b000;
                width14 = 3'b000;
                width13 = 3'b000;
                width12 = 3'b000;
                width11 = 3'b000;
                width10 = 3'b000;
                width9 = 3'b000;
                width8 = 3'b000;
                width7 = 3'b000;
                width6 = 3'b000;
                width5 = 3'b000;
                width4 = 3'b000;
                width3 = 3'b000;
                width2 = 3'b000;
                width1 = 3'b000;

                writeAddr64 = {writeAddr[13:0]};
                writeAddr63 = {writeAddr[13:0]};
                writeAddr62 = {writeAddr[13:0]};
                writeAddr61 = {writeAddr[13:0]};
                writeAddr60 = {writeAddr[13:0]};
                writeAddr59 = {writeAddr[13:0]};
                writeAddr58 = {writeAddr[13:0]};
                writeAddr57 = {writeAddr[13:0]};
                writeAddr56 = {writeAddr[13:0]};
                writeAddr55 = {writeAddr[13:0]};
                writeAddr54 = {writeAddr[13:0]};
                writeAddr53 = {writeAddr[13:0]};
                writeAddr52 = {writeAddr[13:0]};
                writeAddr51 = {writeAddr[13:0]};
                writeAddr50 = {writeAddr[13:0]};
                writeAddr49 = {writeAddr[13:0]};
                writeAddr48 = {writeAddr[13:0]};
                writeAddr47 = {writeAddr[13:0]};
                writeAddr46 = {writeAddr[13:0]};
                writeAddr45 = {writeAddr[13:0]};
                writeAddr44 = {writeAddr[13:0]};
                writeAddr43 = {writeAddr[13:0]};
                writeAddr42 = {writeAddr[13:0]};
                writeAddr41 = {writeAddr[13:0]};
                writeAddr40 = {writeAddr[13:0]};
                writeAddr39 = {writeAddr[13:0]};
                writeAddr38 = {writeAddr[13:0]};
                writeAddr37 = {writeAddr[13:0]};
                writeAddr36 = {writeAddr[13:0]};
                writeAddr35 = {writeAddr[13:0]};
                writeAddr34 = {writeAddr[13:0]};
                writeAddr33 = {writeAddr[13:0]};
                writeAddr32 = {writeAddr[13:0]};
                writeAddr31 = {writeAddr[13:0]};
                writeAddr30 = {writeAddr[13:0]};
                writeAddr29 = {writeAddr[13:0]};
                writeAddr28 = {writeAddr[13:0]};
                writeAddr27 = {writeAddr[13:0]};
                writeAddr26 = {writeAddr[13:0]};
                writeAddr25 = {writeAddr[13:0]};
                writeAddr24 = {writeAddr[13:0]};
                writeAddr23 = {writeAddr[13:0]};
                writeAddr22 = {writeAddr[13:0]};
                writeAddr21 = {writeAddr[13:0]};
                writeAddr20 = {writeAddr[13:0]};
                writeAddr19 = {writeAddr[13:0]};
                writeAddr18 = {writeAddr[13:0]};
                writeAddr17 = {writeAddr[13:0]};
                writeAddr16 = {writeAddr[13:0]};
                writeAddr15 = {writeAddr[13:0]};
                writeAddr14 = {writeAddr[13:0]};
                writeAddr13 = {writeAddr[13:0]};
                writeAddr12 = {writeAddr[13:0]};
                writeAddr11 = {writeAddr[13:0]};
                writeAddr10 = {writeAddr[13:0]};
                writeAddr9 = {writeAddr[13:0]};
                writeAddr8 = {writeAddr[13:0]};
                writeAddr7 = {writeAddr[13:0]};
                writeAddr6 = {writeAddr[13:0]};
                writeAddr5 = {writeAddr[13:0]};
                writeAddr4 = {writeAddr[13:0]};
                writeAddr3 = {writeAddr[13:0]};
                writeAddr2 = {writeAddr[13:0]};
                writeAddr1 = {writeAddr[13:0]};

                readAddr64 = {readAddr[13:0]};
                readAddr63 = {readAddr[13:0]};
                readAddr62 = {readAddr[13:0]};
                readAddr61 = {readAddr[13:0]};
                readAddr60 = {readAddr[13:0]};
                readAddr59 = {readAddr[13:0]};
                readAddr58 = {readAddr[13:0]};
                readAddr57 = {readAddr[13:0]};
                readAddr56 = {readAddr[13:0]};
                readAddr55 = {readAddr[13:0]};
                readAddr54 = {readAddr[13:0]};
                readAddr53 = {readAddr[13:0]};
                readAddr52 = {readAddr[13:0]};
                readAddr51 = {readAddr[13:0]};
                readAddr50 = {readAddr[13:0]};
                readAddr49 = {readAddr[13:0]};
                readAddr48 = {readAddr[13:0]};
                readAddr47 = {readAddr[13:0]};
                readAddr46 = {readAddr[13:0]};
                readAddr45 = {readAddr[13:0]};
                readAddr44 = {readAddr[13:0]};
                readAddr43 = {readAddr[13:0]};
                readAddr42 = {readAddr[13:0]};
                readAddr41 = {readAddr[13:0]};
                readAddr40 = {readAddr[13:0]};
                readAddr39 = {readAddr[13:0]};
                readAddr38 = {readAddr[13:0]};
                readAddr37 = {readAddr[13:0]};
                readAddr36 = {readAddr[13:0]};
                readAddr35 = {readAddr[13:0]};
                readAddr34 = {readAddr[13:0]};
                readAddr33 = {readAddr[13:0]};
                readAddr32 = {readAddr[13:0]};
                readAddr31 = {readAddr[13:0]};
                readAddr30 = {readAddr[13:0]};
                readAddr29 = {readAddr[13:0]};
                readAddr28 = {readAddr[13:0]};
                readAddr27 = {readAddr[13:0]};
                readAddr26 = {readAddr[13:0]};
                readAddr25 = {readAddr[13:0]};
                readAddr24 = {readAddr[13:0]};
                readAddr23 = {readAddr[13:0]};
                readAddr22 = {readAddr[13:0]};
                readAddr21 = {readAddr[13:0]};
                readAddr20 = {readAddr[13:0]};
                readAddr19 = {readAddr[13:0]};
                readAddr18 = {readAddr[13:0]};
                readAddr17 = {readAddr[13:0]};
                readAddr16 = {readAddr[13:0]};
                readAddr15 = {readAddr[13:0]};
                readAddr14 = {readAddr[13:0]};
                readAddr13 = {readAddr[13:0]};
                readAddr12 = {readAddr[13:0]};
                readAddr11 = {readAddr[13:0]};
                readAddr10 = {readAddr[13:0]};
                readAddr9 = {readAddr[13:0]};
                readAddr8 = {readAddr[13:0]};
                readAddr7 = {readAddr[13:0]};
                readAddr6 = {readAddr[13:0]};
                readAddr5 = {readAddr[13:0]};
                readAddr4 = {readAddr[13:0]};
                readAddr3 = {readAddr[13:0]};
                readAddr2 = {readAddr[13:0]};
                readAddr1 = {readAddr[13:0]};

                writeData64 = {17'b0, writeData[31]};
                writeData63 = {17'b0, writeData[30]};
                writeData62 = {17'b0, writeData[29]};
                writeData61 = {17'b0, writeData[28]};
                writeData60 = {17'b0, writeData[27]};
                writeData59 = {17'b0, writeData[26]};
                writeData58 = {17'b0, writeData[25]};
                writeData57 = {17'b0, writeData[24]};
                writeData56 = {17'b0, writeData[23]};
                writeData55 = {17'b0, writeData[22]};
                writeData54 = {17'b0, writeData[21]};
                writeData53 = {17'b0, writeData[20]};
                writeData52 = {17'b0, writeData[19]};
                writeData51 = {17'b0, writeData[18]};
                writeData50 = {17'b0, writeData[17]};
                writeData49 = {17'b0, writeData[16]};
                writeData48 = {17'b0, writeData[15]};
                writeData47 = {17'b0, writeData[14]};
                writeData46 = {17'b0, writeData[13]};
                writeData45 = {17'b0, writeData[12]};
                writeData44 = {17'b0, writeData[11]};
                writeData43 = {17'b0, writeData[10]};
                writeData42 = {17'b0, writeData[9]};
                writeData41 = {17'b0, writeData[8]};
                writeData40 = {17'b0, writeData[7]};
                writeData39 = {17'b0, writeData[6]};
                writeData38 = {17'b0, writeData[5]};
                writeData37 = {17'b0, writeData[4]};
                writeData36 = {17'b0, writeData[3]};
                writeData35 = {17'b0, writeData[2]};
                writeData34 = {17'b0, writeData[1]};
                writeData33 = {17'b0, writeData[0]};
                writeData32 = {17'b0, writeData[31]};
                writeData31 = {17'b0, writeData[30]};
                writeData30 = {17'b0, writeData[29]};
                writeData29 = {17'b0, writeData[28]};
                writeData28 = {17'b0, writeData[27]};
                writeData27 = {17'b0, writeData[26]};
                writeData26 = {17'b0, writeData[25]};
                writeData25 = {17'b0, writeData[24]};
                writeData24 = {17'b0, writeData[23]};
                writeData23 = {17'b0, writeData[22]};
                writeData22 = {17'b0, writeData[21]};
                writeData21 = {17'b0, writeData[20]};
                writeData20 = {17'b0, writeData[19]};
                writeData19 = {17'b0, writeData[18]};
                writeData18 = {17'b0, writeData[17]};
                writeData17 = {17'b0, writeData[16]};
                writeData16 = {17'b0, writeData[15]};
                writeData15 = {17'b0, writeData[14]};
                writeData14 = {17'b0, writeData[13]};
                writeData13 = {17'b0, writeData[12]};
                writeData12 = {17'b0, writeData[11]};
                writeData11 = {17'b0, writeData[10]};
                writeData10 = {17'b0, writeData[9]};
                writeData9 = {17'b0, writeData[8]};
                writeData8 = {17'b0, writeData[7]};
                writeData7 = {17'b0, writeData[6]};
                writeData6 = {17'b0, writeData[5]};
                writeData5 = {17'b0, writeData[4]};
                writeData4 = {17'b0, writeData[3]};
                writeData3 = {17'b0, writeData[2]};
                writeData2 = {17'b0, writeData[1]};
                writeData1 = {17'b0, writeData[0]};

                case (writeAddr[14:9])
                    6'b000000, 6'b000001, 6'b000010, 6'b000011,
                    6'b000100, 6'b000101, 6'b000110, 6'b000111,
                    6'b001000, 6'b001001, 6'b001010, 6'b001011,
                    6'b001100, 6'b001101, 6'b001110, 6'b001111,
                    6'b010000, 6'b010001, 6'b010010, 6'b010011,
                    6'b010100, 6'b010101, 6'b010110, 6'b010111,
                    6'b011000, 6'b011001, 6'b011010, 6'b011011,
                    6'b011100, 6'b011101, 6'b011110, 6'b011111 : begin
                        wen_a64 = {1'b0, wen};
                        wen_a63 = {1'b0, wen};
                        wen_a62 = {1'b0, wen};
                        wen_a61 = {1'b0, wen};
                        wen_a60 = {1'b0, wen};
                        wen_a59 = {1'b0, wen};
                        wen_a58 = {1'b0, wen};
                        wen_a57 = {1'b0, wen};
                        wen_a56 = {1'b0, wen};
                        wen_a55 = {1'b0, wen};
                        wen_a54 = {1'b0, wen};
                        wen_a53 = {1'b0, wen};
                        wen_a52 = {1'b0, wen};
                        wen_a51 = {1'b0, wen};
                        wen_a50 = {1'b0, wen};
                        wen_a49 = {1'b0, wen};
                        wen_a48 = {1'b0, wen};
                        wen_a47 = {1'b0, wen};
                        wen_a46 = {1'b0, wen};
                        wen_a45 = {1'b0, wen};
                        wen_a44 = {1'b0, wen};
                        wen_a43 = {1'b0, wen};
                        wen_a42 = {1'b0, wen};
                        wen_a41 = {1'b0, wen};
                        wen_a40 = {1'b0, wen};
                        wen_a39 = {1'b0, wen};
                        wen_a38 = {1'b0, wen};
                        wen_a37 = {1'b0, wen};
                        wen_a36 = {1'b0, wen};
                        wen_a35 = {1'b0, wen};
                        wen_a34 = {1'b0, wen};
                        wen_a33 = {1'b0, wen};
                        wen_a32 = {1'b0, 1'b0};
                        wen_a31 = {1'b0, 1'b0};
                        wen_a30 = {1'b0, 1'b0};
                        wen_a29 = {1'b0, 1'b0};
                        wen_a28 = {1'b0, 1'b0};
                        wen_a27 = {1'b0, 1'b0};
                        wen_a26 = {1'b0, 1'b0};
                        wen_a25 = {1'b0, 1'b0};
                        wen_a24 = {1'b0, 1'b0};
                        wen_a23 = {1'b0, 1'b0};
                        wen_a22 = {1'b0, 1'b0};
                        wen_a21 = {1'b0, 1'b0};
                        wen_a20 = {1'b0, 1'b0};
                        wen_a19 = {1'b0, 1'b0};
                        wen_a18 = {1'b0, 1'b0};
                        wen_a17 = {1'b0, 1'b0};
                        wen_a16 = {1'b0, 1'b0};
                        wen_a15 = {1'b0, 1'b0};
                        wen_a14 = {1'b0, 1'b0};
                        wen_a13 = {1'b0, 1'b0};
                        wen_a12 = {1'b0, 1'b0};
                        wen_a11 = {1'b0, 1'b0};
                        wen_a10 = {1'b0, 1'b0};
                        wen_a9 = {1'b0, 1'b0};
                        wen_a8 = {1'b0, 1'b0};
                        wen_a7 = {1'b0, 1'b0};
                        wen_a6 = {1'b0, 1'b0};
                        wen_a5 = {1'b0, 1'b0};
                        wen_a4 = {1'b0, 1'b0};
                        wen_a3 = {1'b0, 1'b0};
                        wen_a2 = {1'b0, 1'b0};
                        wen_a1 = {1'b0, 1'b0};
                    end
                    6'b100000, 6'b100001, 6'b100010, 6'b100011,
                    6'b100100, 6'b100101, 6'b100110, 6'b100111,
                    6'b101000, 6'b101001, 6'b101010, 6'b101011,
                    6'b101100, 6'b101101, 6'b101110, 6'b101111,
                    6'b110000, 6'b110001, 6'b110010, 6'b110011,
                    6'b110100, 6'b110101, 6'b110110, 6'b110111,
                    6'b111000, 6'b111001, 6'b111010, 6'b111011,
                    6'b111100, 6'b111101, 6'b111110, 6'b111111 : begin
                        wen_a64 = {1'b0, 1'b0};
                        wen_a63 = {1'b0, 1'b0};
                        wen_a62 = {1'b0, 1'b0};
                        wen_a61 = {1'b0, 1'b0};
                        wen_a60 = {1'b0, 1'b0};
                        wen_a59 = {1'b0, 1'b0};
                        wen_a58 = {1'b0, 1'b0};
                        wen_a57 = {1'b0, 1'b0};
                        wen_a56 = {1'b0, 1'b0};
                        wen_a55 = {1'b0, 1'b0};
                        wen_a54 = {1'b0, 1'b0};
                        wen_a53 = {1'b0, 1'b0};
                        wen_a52 = {1'b0, 1'b0};
                        wen_a51 = {1'b0, 1'b0};
                        wen_a50 = {1'b0, 1'b0};
                        wen_a49 = {1'b0, 1'b0};
                        wen_a48 = {1'b0, 1'b0};
                        wen_a47 = {1'b0, 1'b0};
                        wen_a46 = {1'b0, 1'b0};
                        wen_a45 = {1'b0, 1'b0};
                        wen_a44 = {1'b0, 1'b0};
                        wen_a43 = {1'b0, 1'b0};
                        wen_a42 = {1'b0, 1'b0};
                        wen_a41 = {1'b0, 1'b0};
                        wen_a40 = {1'b0, 1'b0};
                        wen_a39 = {1'b0, 1'b0};
                        wen_a38 = {1'b0, 1'b0};
                        wen_a37 = {1'b0, 1'b0};
                        wen_a36 = {1'b0, 1'b0};
                        wen_a35 = {1'b0, 1'b0};
                        wen_a34 = {1'b0, 1'b0};
                        wen_a33 = {1'b0, 1'b0};
                        wen_a32 = {1'b0, wen};
                        wen_a31 = {1'b0, wen};
                        wen_a30 = {1'b0, wen};
                        wen_a29 = {1'b0, wen};
                        wen_a28 = {1'b0, wen};
                        wen_a27 = {1'b0, wen};
                        wen_a26 = {1'b0, wen};
                        wen_a25 = {1'b0, wen};
                        wen_a24 = {1'b0, wen};
                        wen_a23 = {1'b0, wen};
                        wen_a22 = {1'b0, wen};
                        wen_a21 = {1'b0, wen};
                        wen_a20 = {1'b0, wen};
                        wen_a19 = {1'b0, wen};
                        wen_a18 = {1'b0, wen};
                        wen_a17 = {1'b0, wen};
                        wen_a16 = {1'b0, wen};
                        wen_a15 = {1'b0, wen};
                        wen_a14 = {1'b0, wen};
                        wen_a13 = {1'b0, wen};
                        wen_a12 = {1'b0, wen};
                        wen_a11 = {1'b0, wen};
                        wen_a10 = {1'b0, wen};
                        wen_a9 = {1'b0, wen};
                        wen_a8 = {1'b0, wen};
                        wen_a7 = {1'b0, wen};
                        wen_a6 = {1'b0, wen};
                        wen_a5 = {1'b0, wen};
                        wen_a4 = {1'b0, wen};
                        wen_a3 = {1'b0, wen};
                        wen_a2 = {1'b0, wen};
                        wen_a1 = {1'b0, wen};
                    end
                endcase

                case (ckRdAddr[14:9])
                    6'b000000, 6'b000001, 6'b000010, 6'b000011,
                    6'b000100, 6'b000101, 6'b000110, 6'b000111,
                    6'b001000, 6'b001001, 6'b001010, 6'b001011,
                    6'b001100, 6'b001101, 6'b001110, 6'b001111,
                    6'b010000, 6'b010001, 6'b010010, 6'b010011,
                    6'b010100, 6'b010101, 6'b010110, 6'b010111,
                    6'b011000, 6'b011001, 6'b011010, 6'b011011,
                    6'b011100, 6'b011101, 6'b011110, 6'b011111 : begin
                        readData = {
                                        readData64[0],
                                        readData63[0],
                                        readData62[0],
                                        readData61[0],
                                        readData60[0],
                                        readData59[0],
                                        readData58[0],
                                        readData57[0],
                                        readData56[0],
                                        readData55[0],
                                        readData54[0],
                                        readData53[0],
                                        readData52[0],
                                        readData51[0],
                                        readData50[0],
                                        readData49[0],
                                        readData48[0],
                                        readData47[0],
                                        readData46[0],
                                        readData45[0],
                                        readData44[0],
                                        readData43[0],
                                        readData42[0],
                                        readData41[0],
                                        readData40[0],
                                        readData39[0],
                                        readData38[0],
                                        readData37[0],
                                        readData36[0],
                                        readData35[0],
                                        readData34[0],
                                        readData33[0]
                        };
                    end
                    6'b100000, 6'b100001, 6'b100010, 6'b100011,
                    6'b100100, 6'b100101, 6'b100110, 6'b100111,
                    6'b101000, 6'b101001, 6'b101010, 6'b101011,
                    6'b101100, 6'b101101, 6'b101110, 6'b101111,
                    6'b110000, 6'b110001, 6'b110010, 6'b110011,
                    6'b110100, 6'b110101, 6'b110110, 6'b110111,
                    6'b111000, 6'b111001, 6'b111010, 6'b111011,
                    6'b111100, 6'b111101, 6'b111110, 6'b111111 : begin
                        readData = {
                                        readData32[0],
                                        readData31[0],
                                        readData30[0],
                                        readData29[0],
                                        readData28[0],
                                        readData27[0],
                                        readData26[0],
                                        readData25[0],
                                        readData24[0],
                                        readData23[0],
                                        readData22[0],
                                        readData21[0],
                                        readData20[0],
                                        readData19[0],
                                        readData18[0],
                                        readData17[0],
                                        readData16[0],
                                        readData15[0],
                                        readData14[0],
                                        readData13[0],
                                        readData12[0],
                                        readData11[0],
                                        readData10[0],
                                        readData9[0],
                                        readData8[0],
                                        readData7[0],
                                        readData6[0],
                                        readData5[0],
                                        readData4[0],
                                        readData3[0],
                                        readData2[0],
                                        readData1[0]
                        };
                    end
                endcase
            end        
          33280: begin
                     width64 = 3'b000;
                     width63 = 3'b000;
                     width62 = 3'b000;
                     width61 = 3'b000;
                     width60 = 3'b000;
                     width59 = 3'b000;
                     width58 = 3'b000;
                     width57 = 3'b000;
                     width56 = 3'b000;
                     width55 = 3'b000;
                     width54 = 3'b000;
                     width53 = 3'b000;
                     width52 = 3'b000;
                     width51 = 3'b000;
                     width50 = 3'b000;
                     width49 = 3'b000;
                     width48 = 3'b000;
                     width47 = 3'b000;
                     width46 = 3'b000;
                     width45 = 3'b000;
                     width44 = 3'b000;
                     width43 = 3'b000;
                     width42 = 3'b000;
                     width41 = 3'b000;
                     width40 = 3'b000;
                     width39 = 3'b000;
                     width38 = 3'b000;
                     width37 = 3'b000;
                     width36 = 3'b000;
                     width35 = 3'b000;
                     width34 = 3'b000;
                     width33 = 3'b000;
                     width32 = 3'b000;
                     width31 = 3'b000;
                     width30 = 3'b000;
                     width29 = 3'b000;
                     width28 = 3'b000;
                     width27 = 3'b000;
                     width26 = 3'b000;
                     width25 = 3'b000;
                     width24 = 3'b000;
                     width23 = 3'b000;
                     width22 = 3'b000;
                     width21 = 3'b000;
                     width20 = 3'b000;
                     width19 = 3'b000;
                     width18 = 3'b000;
                     width17 = 3'b000;
                     width16 = 3'b000;
                     width15 = 3'b000;
                     width14 = 3'b000;
                     width13 = 3'b000;
                     width12 = 3'b000;
                     width11 = 3'b000;
                     width10 = 3'b000;
                     width9 = 3'b000;
                     width8 = 3'b000;
                     width7 = 3'b000;
                     width6 = 3'b000;
                     width5 = 3'b000;
                     width4 = 3'b000;
                     width3 = 3'b000;
                     width2 = 3'b000;
                     width1 = 3'b000;
                     width0 = 3'b101;

                    writeAddr64 = {writeAddr[13:0]};
                    writeAddr63 = {writeAddr[13:0]};
                    writeAddr62 = {writeAddr[13:0]};
                    writeAddr61 = {writeAddr[13:0]};
                    writeAddr60 = {writeAddr[13:0]};
                    writeAddr59 = {writeAddr[13:0]};
                    writeAddr58 = {writeAddr[13:0]};
                    writeAddr57 = {writeAddr[13:0]};
                    writeAddr56 = {writeAddr[13:0]};
                    writeAddr55 = {writeAddr[13:0]};
                    writeAddr54 = {writeAddr[13:0]};
                    writeAddr53 = {writeAddr[13:0]};
                    writeAddr52 = {writeAddr[13:0]};
                    writeAddr51 = {writeAddr[13:0]};
                    writeAddr50 = {writeAddr[13:0]};
                    writeAddr49 = {writeAddr[13:0]};
                    writeAddr48 = {writeAddr[13:0]};
                    writeAddr47 = {writeAddr[13:0]};
                    writeAddr46 = {writeAddr[13:0]};
                    writeAddr45 = {writeAddr[13:0]};
                    writeAddr44 = {writeAddr[13:0]};
                    writeAddr43 = {writeAddr[13:0]};
                    writeAddr42 = {writeAddr[13:0]};
                    writeAddr41 = {writeAddr[13:0]};
                    writeAddr40 = {writeAddr[13:0]};
                    writeAddr39 = {writeAddr[13:0]};
                    writeAddr38 = {writeAddr[13:0]};
                    writeAddr37 = {writeAddr[13:0]};
                    writeAddr36 = {writeAddr[13:0]};
                    writeAddr35 = {writeAddr[13:0]};
                    writeAddr34 = {writeAddr[13:0]};
                    writeAddr33 = {writeAddr[13:0]};
                    writeAddr32 = {writeAddr[13:0]};
                    writeAddr31 = {writeAddr[13:0]};
                    writeAddr30 = {writeAddr[13:0]};
                    writeAddr29 = {writeAddr[13:0]};
                    writeAddr28 = {writeAddr[13:0]};
                    writeAddr27 = {writeAddr[13:0]};
                    writeAddr26 = {writeAddr[13:0]};
                    writeAddr25 = {writeAddr[13:0]};
                    writeAddr24 = {writeAddr[13:0]};
                    writeAddr23 = {writeAddr[13:0]};
                    writeAddr22 = {writeAddr[13:0]};
                    writeAddr21 = {writeAddr[13:0]};
                    writeAddr20 = {writeAddr[13:0]};
                    writeAddr19 = {writeAddr[13:0]};
                    writeAddr18 = {writeAddr[13:0]};
                    writeAddr17 = {writeAddr[13:0]};
                    writeAddr16 = {writeAddr[13:0]};
                    writeAddr15 = {writeAddr[13:0]};
                    writeAddr14 = {writeAddr[13:0]};
                    writeAddr13 = {writeAddr[13:0]};
                    writeAddr12 = {writeAddr[13:0]};
                    writeAddr11 = {writeAddr[13:0]};
                    writeAddr10 = {writeAddr[13:0]};
                    writeAddr9 = {writeAddr[13:0]};
                    writeAddr8 = {writeAddr[13:0]};
                    writeAddr7 = {writeAddr[13:0]};
                    writeAddr6 = {writeAddr[13:0]};
                    writeAddr5 = {writeAddr[13:0]};
                    writeAddr4 = {writeAddr[13:0]};
                    writeAddr3 = {writeAddr[13:0]};
                     writeAddr2 = {writeAddr[13:0]};
                     writeAddr1 = {writeAddr[13:0]};
                     writeAddr0 = {writeAddr[8:0], 5'b0};
                         
                    readAddr64 = {readAddr[13:0]};
                    readAddr63 = {readAddr[13:0]};
                    readAddr62 = {readAddr[13:0]};
                    readAddr61 = {readAddr[13:0]};
                    readAddr60 = {readAddr[13:0]};
                    readAddr59 = {readAddr[13:0]};
                    readAddr58 = {readAddr[13:0]};
                    readAddr57 = {readAddr[13:0]};
                    readAddr56 = {readAddr[13:0]};
                    readAddr55 = {readAddr[13:0]};
                    readAddr54 = {readAddr[13:0]};
                    readAddr53 = {readAddr[13:0]};
                    readAddr52 = {readAddr[13:0]};
                    readAddr51 = {readAddr[13:0]};
                    readAddr50 = {readAddr[13:0]};
                    readAddr49 = {readAddr[13:0]};
                    readAddr48 = {readAddr[13:0]};
                    readAddr47 = {readAddr[13:0]};
                    readAddr46 = {readAddr[13:0]};
                    readAddr45 = {readAddr[13:0]};
                    readAddr44 = {readAddr[13:0]};
                    readAddr43 = {readAddr[13:0]};
                    readAddr42 = {readAddr[13:0]};
                    readAddr41 = {readAddr[13:0]};
                    readAddr40 = {readAddr[13:0]};
                    readAddr39 = {readAddr[13:0]};
                    readAddr38 = {readAddr[13:0]};
                    readAddr37 = {readAddr[13:0]};
                    readAddr36 = {readAddr[13:0]};
                    readAddr35 = {readAddr[13:0]};
                    readAddr34 = {readAddr[13:0]};
                    readAddr33 = {readAddr[13:0]};
                    readAddr32 = {readAddr[13:0]};
                    readAddr31 = {readAddr[13:0]};
                    readAddr30 = {readAddr[13:0]};
                    readAddr29 = {readAddr[13:0]};
                    readAddr28 = {readAddr[13:0]};
                    readAddr27 = {readAddr[13:0]};
                    readAddr26 = {readAddr[13:0]};
                    readAddr25 = {readAddr[13:0]};
                    readAddr24 = {readAddr[13:0]};
                    readAddr23 = {readAddr[13:0]};
                    readAddr22 = {readAddr[13:0]};
                    readAddr21 = {readAddr[13:0]};
                    readAddr20 = {readAddr[13:0]};
                    readAddr19 = {readAddr[13:0]};
                    readAddr18 = {readAddr[13:0]};
                    readAddr17 = {readAddr[13:0]};
                    readAddr16 = {readAddr[13:0]};
                    readAddr15 = {readAddr[13:0]};
                    readAddr14 = {readAddr[13:0]};
                    readAddr13 = {readAddr[13:0]};
                    readAddr12 = {readAddr[13:0]};
                    readAddr11 = {readAddr[13:0]};
                    readAddr10 = {readAddr[13:0]};
                    readAddr9 = {readAddr[13:0]};
                    readAddr8 = {readAddr[13:0]};
                    readAddr7 = {readAddr[13:0]};
                    readAddr6 = {readAddr[13:0]};
                    readAddr5 = {readAddr[13:0]};
                    readAddr4 = {readAddr[13:0]};
                    readAddr3 = {readAddr[13:0]};
                     readAddr2 = {readAddr[13:0]};
                     readAddr1 = {readAddr[13:0]};
                     readAddr0 = {readAddr[8:0], 5'b0};
                     
                     writeData64 = {17'b0, writeData[31]};
                     writeData63 = {17'b0, writeData[30]};
                     writeData62 = {17'b0, writeData[29]};
                     writeData61 = {17'b0, writeData[28]};
                     writeData60 = {17'b0, writeData[27]};
                     writeData59 = {17'b0, writeData[26]};
                     writeData58 = {17'b0, writeData[25]};
                     writeData57 = {17'b0, writeData[24]};
                     writeData56 = {17'b0, writeData[23]};
                     writeData55 = {17'b0, writeData[22]};
                     writeData54 = {17'b0, writeData[21]};
                     writeData53 = {17'b0, writeData[20]};
                     writeData52 = {17'b0, writeData[19]};
                     writeData51 = {17'b0, writeData[18]};
                     writeData50 = {17'b0, writeData[17]};
                     writeData49 = {17'b0, writeData[16]};
                     writeData48 = {17'b0, writeData[15]};
                     writeData47 = {17'b0, writeData[14]};
                     writeData46 = {17'b0, writeData[13]};
                     writeData45 = {17'b0, writeData[12]};
                     writeData44 = {17'b0, writeData[11]};
                     writeData43 = {17'b0, writeData[10]};
                     writeData42 = {17'b0, writeData[9]};
                     writeData41 = {17'b0, writeData[8]};
                     writeData40 = {17'b0, writeData[7]};
                     writeData39 = {17'b0, writeData[6]};
                     writeData38 = {17'b0, writeData[5]};
                     writeData37 = {17'b0, writeData[4]};
                     writeData36 = {17'b0, writeData[3]};
                     writeData35 = {17'b0, writeData[2]};
                     writeData34 = {17'b0, writeData[1]};
                     writeData33 = {17'b0, writeData[0]};
                     writeData32 = {17'b0, writeData[31]};
                     writeData31 = {17'b0, writeData[30]};
                     writeData30 = {17'b0, writeData[29]};
                     writeData29 = {17'b0, writeData[28]};
                     writeData28 = {17'b0, writeData[27]};
                     writeData27 = {17'b0, writeData[26]};
                     writeData26 = {17'b0, writeData[25]};
                     writeData25 = {17'b0, writeData[24]};
                     writeData24 = {17'b0, writeData[23]};
                     writeData23 = {17'b0, writeData[22]};
                     writeData22 = {17'b0, writeData[21]};
                     writeData21 = {17'b0, writeData[20]};
                     writeData20 = {17'b0, writeData[19]};
                     writeData19 = {17'b0, writeData[18]};
                     writeData18 = {17'b0, writeData[17]};
                     writeData17 = {17'b0, writeData[16]};
                     writeData16 = {17'b0, writeData[15]};
                     writeData15 = {17'b0, writeData[14]};
                     writeData14 = {17'b0, writeData[13]};
                     writeData13 = {17'b0, writeData[12]};
                     writeData12 = {17'b0, writeData[11]};
                     writeData11 = {17'b0, writeData[10]};
                     writeData10 = {17'b0, writeData[9]};
                     writeData9 = {17'b0, writeData[8]};
                     writeData8 = {17'b0, writeData[7]};
                     writeData7 = {17'b0, writeData[6]};
                     writeData6 = {17'b0, writeData[5]};
                     writeData5 = {17'b0, writeData[4]};
                     writeData4 = {17'b0, writeData[3]};
                     writeData3 = {17'b0, writeData[2]};
                     writeData2 = {17'b0, writeData[1]};
                     writeData1 = {17'b0, writeData[0]};
                     writeData0 = {1'b0, writeData[31:24], 1'b0, writeData[23:16], 1'b0, writeData[15:8], 1'b0, writeData[7:0]};


                     case (writeAddr[15:9])
                       7'b0000000, 7'b0000001, 7'b0000010, 7'b0000011,
                         7'b0000100, 7'b0000101, 7'b0000110, 7'b0000111,
                         7'b0001000, 7'b0001001, 7'b0001010, 7'b0001011,
                         7'b0001100, 7'b0001101, 7'b0001110, 7'b0001111,
                         7'b0010000, 7'b0010001, 7'b0010010, 7'b0010011,
                         7'b0010100, 7'b0010101, 7'b0010110, 7'b0010111,
                         7'b0011000, 7'b0011001, 7'b0011010, 7'b0011011,
                         7'b0011100, 7'b0011101, 7'b0011110, 7'b0011111 : begin
                            wen_a64 = {1'b0, wen};
                            wen_a63 = {1'b0, wen};
                            wen_a62 = {1'b0, wen};
                            wen_a61 = {1'b0, wen};
                            wen_a60 = {1'b0, wen};
                            wen_a59 = {1'b0, wen};
                            wen_a58 = {1'b0, wen};
                            wen_a57 = {1'b0, wen};
                            wen_a56 = {1'b0, wen};
                            wen_a55 = {1'b0, wen};
                            wen_a54 = {1'b0, wen};
                            wen_a53 = {1'b0, wen};
                            wen_a52 = {1'b0, wen};
                            wen_a51 = {1'b0, wen};
                            wen_a50 = {1'b0, wen};
                            wen_a49 = {1'b0, wen};
                            wen_a48 = {1'b0, wen};
                            wen_a47 = {1'b0, wen};
                            wen_a46 = {1'b0, wen};
                            wen_a45 = {1'b0, wen};
                            wen_a44 = {1'b0, wen};
                            wen_a43 = {1'b0, wen};
                            wen_a42 = {1'b0, wen};
                            wen_a41 = {1'b0, wen};
                            wen_a40 = {1'b0, wen};
                            wen_a39 = {1'b0, wen};
                            wen_a38 = {1'b0, wen};
                            wen_a37 = {1'b0, wen};
                            wen_a36 = {1'b0, wen};
                            wen_a35 = {1'b0, wen};
                            wen_a34 = {1'b0, wen};
                            wen_a33 = {1'b0, wen};
                            wen_a32 = {1'b0, 1'b0};
                            wen_a31 = {1'b0, 1'b0};
                            wen_a30 = {1'b0, 1'b0};
                            wen_a29 = {1'b0, 1'b0};
                            wen_a28 = {1'b0, 1'b0};
                            wen_a27 = {1'b0, 1'b0};
                            wen_a26 = {1'b0, 1'b0};
                            wen_a25 = {1'b0, 1'b0};
                            wen_a24 = {1'b0, 1'b0};
                            wen_a23 = {1'b0, 1'b0};
                            wen_a22 = {1'b0, 1'b0};
                            wen_a21 = {1'b0, 1'b0};
                            wen_a20 = {1'b0, 1'b0};
                            wen_a19 = {1'b0, 1'b0};
                            wen_a18 = {1'b0, 1'b0};
                            wen_a17 = {1'b0, 1'b0};
                            wen_a16 = {1'b0, 1'b0};
                            wen_a15 = {1'b0, 1'b0};
                            wen_a14 = {1'b0, 1'b0};
                            wen_a13 = {1'b0, 1'b0};
                            wen_a12 = {1'b0, 1'b0};
                            wen_a11 = {1'b0, 1'b0};
                            wen_a10 = {1'b0, 1'b0};
                            wen_a9  = {1'b0, 1'b0};
                            wen_a8  = {1'b0, 1'b0};
                            wen_a7  = {1'b0, 1'b0};
                            wen_a6  = {1'b0, 1'b0};
                            wen_a5  = {1'b0, 1'b0};
                            wen_a4  = {1'b0, 1'b0};
                            wen_a3  = {1'b0, 1'b0};
                            wen_a2  = {1'b0, 1'b0};
                            wen_a1  = {1'b0, 1'b0};
                            wen_a0  = {1'b0, 1'b0};
                            wen_b0  = {1'b0, 1'b0};
                         end
                         7'b0100000, 7'b0100001, 7'b0100010, 7'b0100011,
                         7'b0100100, 7'b0100101, 7'b0100110, 7'b0100111,
                         7'b0101000, 7'b0101001, 7'b0101010, 7'b0101011,
                         7'b0101100, 7'b0101101, 7'b0101110, 7'b0101111,
                         7'b0110000, 7'b0110001, 7'b0110010, 7'b0110011,
                         7'b0110100, 7'b0110101, 7'b0110110, 7'b0110111,             
                         7'b0111000, 7'b0111001, 7'b0111010, 7'b0111011,
                         7'b0111100, 7'b0111101, 7'b0111110, 7'b0111111  : begin
                            wen_a64 = {1'b0, 1'b0};
                            wen_a63 = {1'b0, 1'b0};
                            wen_a62 = {1'b0, 1'b0};
                            wen_a61 = {1'b0, 1'b0};
                            wen_a60 = {1'b0, 1'b0};
                            wen_a59 = {1'b0, 1'b0};
                            wen_a58 = {1'b0, 1'b0};
                            wen_a57 = {1'b0, 1'b0};
                            wen_a56 = {1'b0, 1'b0};
                            wen_a55 = {1'b0, 1'b0};
                            wen_a54 = {1'b0, 1'b0};
                            wen_a53 = {1'b0, 1'b0};
                            wen_a52 = {1'b0, 1'b0};
                            wen_a51 = {1'b0, 1'b0};
                            wen_a50 = {1'b0, 1'b0};
                            wen_a49 = {1'b0, 1'b0};
                            wen_a48 = {1'b0, 1'b0};
                            wen_a47 = {1'b0, 1'b0};
                            wen_a46 = {1'b0, 1'b0};
                            wen_a45 = {1'b0, 1'b0};
                            wen_a44 = {1'b0, 1'b0};
                            wen_a43 = {1'b0, 1'b0};
                            wen_a42 = {1'b0, 1'b0};
                            wen_a41 = {1'b0, 1'b0};
                            wen_a40 = {1'b0, 1'b0};
                            wen_a39 = {1'b0, 1'b0};
                            wen_a38 = {1'b0, 1'b0};
                            wen_a37 = {1'b0, 1'b0};
                            wen_a36 = {1'b0, 1'b0};
                            wen_a35 = {1'b0, 1'b0};
                            wen_a34 = {1'b0, 1'b0};
                            wen_a33 = {1'b0, 1'b0};
                            wen_a32 = {1'b0, wen};
                            wen_a31 = {1'b0, wen};
                            wen_a30 = {1'b0, wen};
                            wen_a29 = {1'b0, wen};
                            wen_a28 = {1'b0, wen};
                            wen_a27 = {1'b0, wen};
                            wen_a26 = {1'b0, wen};
                            wen_a25 = {1'b0, wen};
                            wen_a24 = {1'b0, wen};
                            wen_a23 = {1'b0, wen};
                            wen_a22 = {1'b0, wen};
                            wen_a21 = {1'b0, wen};
                            wen_a20 = {1'b0, wen};
                            wen_a19 = {1'b0, wen};
                            wen_a18 = {1'b0, wen};
                            wen_a17 = {1'b0, wen};
                            wen_a16 = {1'b0, wen};
                            wen_a15 = {1'b0, wen};
                            wen_a14 = {1'b0, wen};
                            wen_a13 = {1'b0, wen};
                            wen_a12 = {1'b0, wen};
                            wen_a11 = {1'b0, wen};
                            wen_a10 = {1'b0, wen};
                            wen_a9 = {1'b0, wen};
                            wen_a8 = {1'b0, wen};
                            wen_a7 = {1'b0, wen};
                            wen_a6 = {1'b0, wen};
                            wen_a5 = {1'b0, wen};
                            wen_a4 = {1'b0, wen};
                            wen_a3 = {1'b0, wen};
                            wen_a2 = {1'b0, wen};
                            wen_a1 = {1'b0, wen};
                            wen_a0 = {1'b0, 1'b0};
                            wen_b0 = {1'b0, 1'b0};

                         end
                       7'b1000000 : begin
                        wen_a64 = {1'b0, 1'b0};
                        wen_a63 = {1'b0, 1'b0};
                        wen_a62 = {1'b0, 1'b0};
                        wen_a61 = {1'b0, 1'b0};
                        wen_a60 = {1'b0, 1'b0};
                        wen_a59 = {1'b0, 1'b0};
                        wen_a58 = {1'b0, 1'b0};
                        wen_a57 = {1'b0, 1'b0};
                        wen_a56 = {1'b0, 1'b0};
                        wen_a55 = {1'b0, 1'b0};
                        wen_a54 = {1'b0, 1'b0};
                        wen_a53 = {1'b0, 1'b0};
                        wen_a52 = {1'b0, 1'b0};
                        wen_a51 = {1'b0, 1'b0};
                        wen_a50 = {1'b0, 1'b0};
                        wen_a49 = {1'b0, 1'b0};
                        wen_a48 = {1'b0, 1'b0};
                        wen_a47 = {1'b0, 1'b0};
                        wen_a46 = {1'b0, 1'b0};
                        wen_a45 = {1'b0, 1'b0};
                        wen_a44 = {1'b0, 1'b0};
                        wen_a43 = {1'b0, 1'b0};
                        wen_a42 = {1'b0, 1'b0};
                        wen_a41 = {1'b0, 1'b0};
                        wen_a40 = {1'b0, 1'b0};
                        wen_a39 = {1'b0, 1'b0};
                        wen_a38 = {1'b0, 1'b0};
                        wen_a37 = {1'b0, 1'b0};
                        wen_a36 = {1'b0, 1'b0};
                        wen_a35 = {1'b0, 1'b0};
                        wen_a34 = {1'b0, 1'b0};
                        wen_a33 = {1'b0, 1'b0};
                        wen_a32 = {1'b0, 1'b0};
                        wen_a31 = {1'b0, 1'b0};
                        wen_a30 = {1'b0, 1'b0};
                        wen_a29 = {1'b0, 1'b0};
                        wen_a28 = {1'b0, 1'b0};
                        wen_a27 = {1'b0, 1'b0};
                        wen_a26 = {1'b0, 1'b0};
                        wen_a25 = {1'b0, 1'b0};
                        wen_a24 = {1'b0, 1'b0};
                        wen_a23 = {1'b0, 1'b0};
                        wen_a22 = {1'b0, 1'b0};
                        wen_a21 = {1'b0, 1'b0};
                        wen_a20 = {1'b0, 1'b0};
                        wen_a19 = {1'b0, 1'b0};
                        wen_a18 = {1'b0, 1'b0};
                        wen_a17 = {1'b0, 1'b0};
                        wen_a16 = {1'b0, 1'b0};
                        wen_a15 = {1'b0, 1'b0};
                        wen_a14 = {1'b0, 1'b0};
                        wen_a13 = {1'b0, 1'b0};
                        wen_a12 = {1'b0, 1'b0};
                        wen_a11 = {1'b0, 1'b0};
                        wen_a10 = {1'b0, 1'b0};
                        wen_a9 =  {1'b0, 1'b0};
                        wen_a8 =  {1'b0, 1'b0};
                        wen_a7 =  {1'b0, 1'b0};
                        wen_a6 =  {1'b0, 1'b0};
                        wen_a5 =  {1'b0, 1'b0};
                        wen_a4 =  {1'b0, 1'b0};
                        wen_a3 = {1'b0, 1'b0};
                        wen_a2 = {1'b0, 1'b0};
                        wen_a1 = {1'b0, 1'b0};
                        wen_a0 = {wen, wen};
                        wen_b0 = {wen, wen};
                    end
                       default : begin
                        wen_a64 = {1'b0, 1'b0};
                        wen_a63 = {1'b0, 1'b0};
                        wen_a62 = {1'b0, 1'b0};
                        wen_a61 = {1'b0, 1'b0};
                        wen_a60 = {1'b0, 1'b0};
                        wen_a59 = {1'b0, 1'b0};
                        wen_a58 = {1'b0, 1'b0};
                        wen_a57 = {1'b0, 1'b0};
                        wen_a56 = {1'b0, 1'b0};
                        wen_a55 = {1'b0, 1'b0};
                        wen_a54 = {1'b0, 1'b0};
                        wen_a53 = {1'b0, 1'b0};
                        wen_a52 = {1'b0, 1'b0};
                        wen_a51 = {1'b0, 1'b0};
                        wen_a50 = {1'b0, 1'b0};
                        wen_a49 = {1'b0, 1'b0};
                        wen_a48 = {1'b0, 1'b0};
                        wen_a47 = {1'b0, 1'b0};
                        wen_a46 = {1'b0, 1'b0};
                        wen_a45 = {1'b0, 1'b0};
                        wen_a44 = {1'b0, 1'b0};
                        wen_a43 = {1'b0, 1'b0};
                        wen_a42 = {1'b0, 1'b0};
                        wen_a41 = {1'b0, 1'b0};
                        wen_a40 = {1'b0, 1'b0};
                        wen_a39 = {1'b0, 1'b0};
                        wen_a38 = {1'b0, 1'b0};
                        wen_a37 = {1'b0, 1'b0};
                        wen_a36 = {1'b0, 1'b0};
                        wen_a35 = {1'b0, 1'b0};
                        wen_a34 = {1'b0, 1'b0};
                        wen_a33 = {1'b0, 1'b0};
                        wen_a32 = {1'b0, 1'b0};
                        wen_a31 = {1'b0, 1'b0};
                        wen_a30 = {1'b0, 1'b0};
                        wen_a29 = {1'b0, 1'b0};
                        wen_a28 = {1'b0, 1'b0};
                        wen_a27 = {1'b0, 1'b0};
                        wen_a26 = {1'b0, 1'b0};
                        wen_a25 = {1'b0, 1'b0};
                        wen_a24 = {1'b0, 1'b0};
                        wen_a23 = {1'b0, 1'b0};
                        wen_a22 = {1'b0, 1'b0};
                        wen_a21 = {1'b0, 1'b0};
                        wen_a20 = {1'b0, 1'b0};
                        wen_a19 = {1'b0, 1'b0};
                        wen_a18 = {1'b0, 1'b0};
                        wen_a17 = {1'b0, 1'b0};
                        wen_a16 = {1'b0, 1'b0};
                        wen_a15 = {1'b0, 1'b0};
                        wen_a14 = {1'b0, 1'b0};
                        wen_a13 = {1'b0, 1'b0};
                        wen_a12 = {1'b0, 1'b0};
                        wen_a11 = {1'b0, 1'b0};
                        wen_a10 = {1'b0, 1'b0};
                        wen_a9 =  {1'b0, 1'b0};
                        wen_a8 =  {1'b0, 1'b0};
                        wen_a7 =  {1'b0, 1'b0};
                        wen_a6 =  {1'b0, 1'b0};
                        wen_a5 =  {1'b0, 1'b0};
                        wen_a4 =  {1'b0, 1'b0};
                        wen_a3 = {1'b0, 1'b0};
                        wen_a2 = {1'b0, 1'b0};
                        wen_a1 = {1'b0, 1'b0};
                        wen_a0 = {1'b0, 1'b0};
                        wen_b0 = {1'b0, 1'b0};
                       end
                     endcase // case (writeAddr[14:9])
                     

                     case (ckRdAddr[15:9])
                       7'b0000000, 7'b0000001, 7'b0000010, 7'b0000011,
                         7'b0000100, 7'b0000101, 7'b0000110, 7'b0000111,
                         7'b0001000, 7'b0001001, 7'b0001010, 7'b0001011,
                         7'b0001100, 7'b0001101, 7'b0001110, 7'b0001111,
                         7'b0010000, 7'b0010001, 7'b0010010, 7'b0010011,
                         7'b0010100, 7'b0010101, 7'b0010110, 7'b0010111,
                         7'b0011000, 7'b0011001, 7'b0011010, 7'b0011011,
                         7'b0011100, 7'b0011101, 7'b0011110, 7'b0011111  : begin

                            readData = {
                                        readData64[0],
                                        readData63[0],
                                        readData62[0],
                                        readData61[0],
                                        readData60[0],
                                        readData59[0],
                                        readData58[0],
                                        readData57[0],
                                        readData56[0],
                                        readData55[0], 
                                        readData54[0],
                                        readData53[0],
                                        readData52[0],
                                        readData51[0],
                                        readData50[0],
                                        readData49[0],
                                        readData48[0],
                                        readData47[0],
                                        readData46[0],
                                        readData45[0],
                                        readData44[0],
                                        readData43[0],
                                        readData42[0],
                                        readData41[0],
                                        readData40[0],
                                        readData39[0],
                                        readData38[0],
                                        readData37[0],
                                        readData36[0],
                                        readData35[0],
                                        readData34[0],
                                        readData33[0]                                        
                                        };
                         end // case: 7'b0000000, 7'b0000001, 7'b0000010, 7'b0000011,...
                       7'b0100000, 7'b0100001, 7'b0100010, 7'b0100011,
                         7'b0100100, 7'b0100101, 7'b0100110, 7'b0100111,
                         7'b0101000, 7'b0101001, 7'b0101010, 7'b0101011,
                         7'b0101100, 7'b0101101, 7'b0101110, 7'b0101111,
                         7'b0110000, 7'b0110001, 7'b0110010, 7'b0110011,
                         7'b0110100, 7'b0110101, 7'b0110110, 7'b0110111,             
                         7'b0111000, 7'b0111001, 7'b0111010, 7'b0111011,
                         7'b0111100, 7'b0111101, 7'b0111110, 7'b0111111 : begin
                            readData = {
                                        readData32[0],                
                                        readData31[0],
                                        readData30[0],
                                        readData29[0],
                                        readData28[0],
                                        readData27[0],
                                        readData26[0],
                                        readData25[0],
                                        readData24[0],
                                        readData23[0],
                                        readData22[0],
                                        readData21[0],
                                        readData20[0],
                                        readData19[0],
                                        readData18[0],
                                        readData17[0],
                                        readData16[0],
                                        readData15[0],
                                        readData14[0],
                                        readData13[0],
                                        readData12[0],
                                        readData11[0],
                                        readData10[0],
                                        readData9[0],
                                        readData8[0],
                                        readData7[0],
                                        readData6[0],
                                        readData5[0],
                                        readData4[0],
                                        readData3[0],
                                        readData2[0],
                                        readData1[0]};
                       end
                       7'b1000000 : begin
                          readData = {readData0[34:27],readData0[25:18],readData0[16:9],readData0[7:0]};
                       end
                       default : begin
                          readData = 32'b0;
                       end
                     endcase // case (ckRdAddr[14:9])                     
          end // case: 33280

          33792: begin
                     width66 = 3'b000;
                     width65 = 3'b000;
                     width64 = 3'b000;
                     width63 = 3'b000;
                     width62 = 3'b000;
                     width61 = 3'b000;
                     width60 = 3'b000;
                     width59 = 3'b000;
                     width58 = 3'b000;
                     width57 = 3'b000;
                     width56 = 3'b000;
                     width55 = 3'b000;
                     width54 = 3'b000;
                     width53 = 3'b000;
                     width52 = 3'b000;
                     width51 = 3'b000;
                     width50 = 3'b000;
                     width49 = 3'b000;
                     width48 = 3'b000;
                     width47 = 3'b000;
                     width46 = 3'b000;
                     width45 = 3'b000;
                     width44 = 3'b000;
                     width43 = 3'b000;
                     width42 = 3'b000;
                     width41 = 3'b000;
                     width40 = 3'b000;
                     width39 = 3'b000;
                     width38 = 3'b000;
                     width37 = 3'b000;
                     width36 = 3'b000;
                     width35 = 3'b000;
                     width34 = 3'b000;
                     width33 = 3'b000;
                     width32 = 3'b000;
                     width31 = 3'b000;
                     width30 = 3'b000;
                     width29 = 3'b000;
                     width28 = 3'b000;
                     width27 = 3'b000;
                     width26 = 3'b000;
                     width25 = 3'b000;
                     width24 = 3'b000;
                     width23 = 3'b000;
                     width22 = 3'b000;
                     width21 = 3'b000;
                     width20 = 3'b000;
                     width19 = 3'b000;
                     width18 = 3'b000;
                     width17 = 3'b000;
                     width16 = 3'b000;
                     width15 = 3'b000;
                     width14 = 3'b000;
                     width13 = 3'b000;
                     width12 = 3'b000;
                     width11 = 3'b000;
                     width10 = 3'b000;
                     width9 = 3'b000;
                     width8 = 3'b000;
                     width7 = 3'b000;
                     width6 = 3'b000;
                     width5 = 3'b000;
                     width4 = 3'b000;
                     width3 = 3'b000;
                     width2 = 3'b100;
                     width1 = 3'b100;


                    writeAddr66 = {writeAddr[13:0]};
                    writeAddr65 = {writeAddr[13:0]};
                    writeAddr64 = {writeAddr[13:0]};
                    writeAddr63 = {writeAddr[13:0]};
                    writeAddr62 = {writeAddr[13:0]};
                    writeAddr61 = {writeAddr[13:0]};
                    writeAddr60 = {writeAddr[13:0]};
                    writeAddr59 = {writeAddr[13:0]};
                    writeAddr58 = {writeAddr[13:0]};
                    writeAddr57 = {writeAddr[13:0]};
                    writeAddr56 = {writeAddr[13:0]};
                    writeAddr55 = {writeAddr[13:0]};
                    writeAddr54 = {writeAddr[13:0]};
                    writeAddr53 = {writeAddr[13:0]};
                    writeAddr52 = {writeAddr[13:0]};
                    writeAddr51 = {writeAddr[13:0]};
                    writeAddr50 = {writeAddr[13:0]};
                    writeAddr49 = {writeAddr[13:0]};
                    writeAddr48 = {writeAddr[13:0]};
                    writeAddr47 = {writeAddr[13:0]};
                    writeAddr46 = {writeAddr[13:0]};
                    writeAddr45 = {writeAddr[13:0]};
                    writeAddr44 = {writeAddr[13:0]};
                    writeAddr43 = {writeAddr[13:0]};
                    writeAddr42 = {writeAddr[13:0]};
                    writeAddr41 = {writeAddr[13:0]};
                    writeAddr40 = {writeAddr[13:0]};
                    writeAddr39 = {writeAddr[13:0]};
                    writeAddr38 = {writeAddr[13:0]};
                    writeAddr37 = {writeAddr[13:0]};
                    writeAddr36 = {writeAddr[13:0]};
                    writeAddr35 = {writeAddr[13:0]};
                    writeAddr34 = {writeAddr[13:0]};
                    writeAddr33 = {writeAddr[13:0]};
                    writeAddr32 = {writeAddr[13:0]};
                    writeAddr31 = {writeAddr[13:0]};
                    writeAddr30 = {writeAddr[13:0]};
                    writeAddr29 = {writeAddr[13:0]};
                    writeAddr28 = {writeAddr[13:0]};
                    writeAddr27 = {writeAddr[13:0]};
                    writeAddr26 = {writeAddr[13:0]};
                    writeAddr25 = {writeAddr[13:0]};
                    writeAddr24 = {writeAddr[13:0]};
                    writeAddr23 = {writeAddr[13:0]};
                    writeAddr22 = {writeAddr[13:0]};
                    writeAddr21 = {writeAddr[13:0]};
                    writeAddr20 = {writeAddr[13:0]};
                    writeAddr19 = {writeAddr[13:0]};
                    writeAddr18 = {writeAddr[13:0]};
                    writeAddr17 = {writeAddr[13:0]};
                    writeAddr16 = {writeAddr[13:0]};
                    writeAddr15 = {writeAddr[13:0]};
                    writeAddr14 = {writeAddr[13:0]};
                    writeAddr13 = {writeAddr[13:0]};
                    writeAddr12 = {writeAddr[13:0]};
                    writeAddr11 = {writeAddr[13:0]};
                    writeAddr10 = {writeAddr[13:0]};
                    writeAddr9 = {writeAddr[13:0]};
                    writeAddr8 = {writeAddr[13:0]};
                    writeAddr7 = {writeAddr[13:0]};
                    writeAddr6 = {writeAddr[13:0]};
                    writeAddr5 = {writeAddr[13:0]};
                    writeAddr4 = {writeAddr[13:0]};
             writeAddr3 = {writeAddr[13:0]};
             writeAddr2 = {writeAddr[9:0], 4'b0};
             writeAddr1 = {writeAddr[9:0], 4'b0};

                    readAddr66 = {readAddr[13:0]};                         
                    readAddr65 = {readAddr[13:0]};
                    readAddr64 = {readAddr[13:0]};
                    readAddr63 = {readAddr[13:0]};
                    readAddr62 = {readAddr[13:0]};
                    readAddr61 = {readAddr[13:0]};
                    readAddr60 = {readAddr[13:0]};
                    readAddr59 = {readAddr[13:0]};
                    readAddr58 = {readAddr[13:0]};
                    readAddr57 = {readAddr[13:0]};
                    readAddr56 = {readAddr[13:0]};
                    readAddr55 = {readAddr[13:0]};
                    readAddr54 = {readAddr[13:0]};
                    readAddr53 = {readAddr[13:0]};
                    readAddr52 = {readAddr[13:0]};
                    readAddr51 = {readAddr[13:0]};
                    readAddr50 = {readAddr[13:0]};
                    readAddr49 = {readAddr[13:0]};
                    readAddr48 = {readAddr[13:0]};
                    readAddr47 = {readAddr[13:0]};
                    readAddr46 = {readAddr[13:0]};
                    readAddr45 = {readAddr[13:0]};
                    readAddr44 = {readAddr[13:0]};
                    readAddr43 = {readAddr[13:0]};
                    readAddr42 = {readAddr[13:0]};
                    readAddr41 = {readAddr[13:0]};
                    readAddr40 = {readAddr[13:0]};
                    readAddr39 = {readAddr[13:0]};
                    readAddr38 = {readAddr[13:0]};
                    readAddr37 = {readAddr[13:0]};
                    readAddr36 = {readAddr[13:0]};
                    readAddr35 = {readAddr[13:0]};
                    readAddr34 = {readAddr[13:0]};
                    readAddr33 = {readAddr[13:0]};
                    readAddr32 = {readAddr[13:0]};
                    readAddr31 = {readAddr[13:0]};
                    readAddr30 = {readAddr[13:0]};
                    readAddr29 = {readAddr[13:0]};
                    readAddr28 = {readAddr[13:0]};
                    readAddr27 = {readAddr[13:0]};
                    readAddr26 = {readAddr[13:0]};
                    readAddr25 = {readAddr[13:0]};
                    readAddr24 = {readAddr[13:0]};
                    readAddr23 = {readAddr[13:0]};
                    readAddr22 = {readAddr[13:0]};
                    readAddr21 = {readAddr[13:0]};
                    readAddr20 = {readAddr[13:0]};
                    readAddr19 = {readAddr[13:0]};
                    readAddr18 = {readAddr[13:0]};
                    readAddr17 = {readAddr[13:0]};
                    readAddr16 = {readAddr[13:0]};
                    readAddr15 = {readAddr[13:0]};
                    readAddr14 = {readAddr[13:0]};
                    readAddr13 = {readAddr[13:0]};
                    readAddr12 = {readAddr[13:0]};
                    readAddr11 = {readAddr[13:0]};
                    readAddr10 = {readAddr[13:0]};
                    readAddr9 = {readAddr[13:0]};
                    readAddr8 = {readAddr[13:0]};
                    readAddr7 = {readAddr[13:0]};
                    readAddr6 = {readAddr[13:0]};
                    readAddr5 = {readAddr[13:0]};
                    readAddr4 = {readAddr[13:0]};
                    readAddr3 = {readAddr[13:0]};
                    readAddr2  = {readAddr[9:0],  4'b0};
                    readAddr1  = {readAddr[9:0],  4'b0};
                     
                     writeData66 = {17'b0, writeData[31]};
                     writeData65 = {17'b0, writeData[30]};
                     writeData64 = {17'b0, writeData[29]};
                     writeData63 = {17'b0, writeData[28]};
                     writeData62 = {17'b0, writeData[27]};
                     writeData61 = {17'b0, writeData[26]};
                     writeData60 = {17'b0, writeData[25]};
                     writeData59 = {17'b0, writeData[24]};
                     writeData58 = {17'b0, writeData[23]};
                     writeData57 = {17'b0, writeData[22]};
                     writeData56 = {17'b0, writeData[21]};
                     writeData55 = {17'b0, writeData[20]};
                     writeData54 = {17'b0, writeData[19]};
                     writeData53 = {17'b0, writeData[18]};
                     writeData52 = {17'b0, writeData[17]};
                     writeData51 = {17'b0, writeData[16]};
                     writeData50 = {17'b0, writeData[15]};
                     writeData49 = {17'b0, writeData[14]};
                     writeData48 = {17'b0, writeData[13]};
                     writeData47 = {17'b0, writeData[12]};
                     writeData46 = {17'b0, writeData[11]};
                     writeData45 = {17'b0, writeData[10]};
                     writeData44 = {17'b0, writeData[9]};
                     writeData43 = {17'b0, writeData[8]};
                     writeData42 = {17'b0, writeData[7]};
                     writeData41 = {17'b0, writeData[6]};
                     writeData40 = {17'b0, writeData[5]};
                     writeData39 = {17'b0, writeData[4]};
                     writeData38 = {17'b0, writeData[3]};
                     writeData37 = {17'b0, writeData[2]};
                     writeData36 = {17'b0, writeData[1]};
                     writeData35 = {17'b0, writeData[0]};
                     writeData34 = {17'b0, writeData[31]};
                     writeData33 = {17'b0, writeData[30]};
                     writeData32 = {17'b0, writeData[29]};
                     writeData31 = {17'b0, writeData[28]};
                     writeData30 = {17'b0, writeData[27]};
                     writeData29 = {17'b0, writeData[26]};
                     writeData28 = {17'b0, writeData[25]};
                     writeData27 = {17'b0, writeData[24]};
                     writeData26 = {17'b0, writeData[23]};
                     writeData25 = {17'b0, writeData[22]};
                     writeData24 = {17'b0, writeData[21]};
                     writeData23 = {17'b0, writeData[20]};
                     writeData22 = {17'b0, writeData[19]};
                     writeData21 = {17'b0, writeData[18]};
                     writeData20 = {17'b0, writeData[17]};
                     writeData19 = {17'b0, writeData[16]};
                     writeData18 = {17'b0, writeData[15]};
                     writeData17 = {17'b0, writeData[14]};
                     writeData16 = {17'b0, writeData[13]};
                     writeData15 = {17'b0, writeData[12]};
                     writeData14 = {17'b0, writeData[11]};
                     writeData13 = {17'b0, writeData[10]};
                     writeData12 = {17'b0, writeData[9]};
                     writeData11 = {17'b0, writeData[8]};
                     writeData10 = {17'b0, writeData[7]};
                     writeData9 = {17'b0, writeData[6]};
                     writeData8 = {17'b0, writeData[5]};
                     writeData7 = {17'b0, writeData[4]};
                     writeData6 = {17'b0, writeData[3]};
                     writeData5 = {17'b0, writeData[2]};
                     writeData4 = {17'b0, writeData[1]};
                     writeData3 = {17'b0, writeData[0]};
                     writeData2 = {1'b0, writeData[31:24], 1'b0, writeData[23:16]};
                     writeData1 = {1'b0, writeData[15:8], 1'b0, writeData[7:0]};


                case (writeAddr[15:9])
                       7'b0000000, 7'b0000001, 7'b0000010, 7'b0000011,
                         7'b0000100, 7'b0000101, 7'b0000110, 7'b0000111,
                         7'b0001000, 7'b0001001, 7'b0001010, 7'b0001011,
                         7'b0001100, 7'b0001101, 7'b0001110, 7'b0001111,
                         7'b0010000, 7'b0010001, 7'b0010010, 7'b0010011,
                         7'b0010100, 7'b0010101, 7'b0010110, 7'b0010111,
                         7'b0011000, 7'b0011001, 7'b0011010, 7'b0011011,
                         7'b0011100, 7'b0011101, 7'b0011110, 7'b0011111 : begin
                            wen_a66 = {1'b0, wen};
                            wen_a65 = {1'b0, wen};
                            wen_a64 = {1'b0, wen};
                            wen_a63 = {1'b0, wen};
                            wen_a62 = {1'b0, wen};
                            wen_a61 = {1'b0, wen};
                            wen_a60 = {1'b0, wen};
                            wen_a59 = {1'b0, wen};
                            wen_a58 = {1'b0, wen};
                            wen_a57 = {1'b0, wen};
                            wen_a56 = {1'b0, wen};
                            wen_a55 = {1'b0, wen};
                            wen_a54 = {1'b0, wen};
                            wen_a53 = {1'b0, wen};
                            wen_a52 = {1'b0, wen};
                            wen_a51 = {1'b0, wen};
                            wen_a50 = {1'b0, wen};
                            wen_a49 = {1'b0, wen};
                            wen_a48 = {1'b0, wen};
                            wen_a47 = {1'b0, wen};
                            wen_a46 = {1'b0, wen};
                            wen_a45 = {1'b0, wen};
                            wen_a44 = {1'b0, wen};
                            wen_a43 = {1'b0, wen};
                            wen_a42 = {1'b0, wen};
                            wen_a41 = {1'b0, wen};
                            wen_a40 = {1'b0, wen};
                            wen_a39 = {1'b0, wen};
                            wen_a38 = {1'b0, wen};
                            wen_a37 = {1'b0, wen};
                            wen_a36 = {1'b0, wen};
                            wen_a35 = {1'b0, wen};
                            wen_a34 = {1'b0, 1'b0};
                            wen_a33 = {1'b0, 1'b0};
                            wen_a32 = {1'b0, 1'b0};
                            wen_a31 = {1'b0, 1'b0};
                            wen_a30 = {1'b0, 1'b0};
                            wen_a29 = {1'b0, 1'b0};
                            wen_a28 = {1'b0, 1'b0};
                            wen_a27 = {1'b0, 1'b0};
                            wen_a26 = {1'b0, 1'b0};
                            wen_a25 = {1'b0, 1'b0};
                            wen_a24 = {1'b0, 1'b0};
                            wen_a23 = {1'b0, 1'b0};
                            wen_a22 = {1'b0, 1'b0};
                            wen_a21 = {1'b0, 1'b0};
                            wen_a20 = {1'b0, 1'b0};
                            wen_a19 = {1'b0, 1'b0};
                            wen_a18 = {1'b0, 1'b0};
                            wen_a17 = {1'b0, 1'b0};
                            wen_a16 = {1'b0, 1'b0};
                            wen_a15 = {1'b0, 1'b0};
                            wen_a14 = {1'b0, 1'b0};
                            wen_a13 = {1'b0, 1'b0};
                            wen_a12 = {1'b0, 1'b0};
                            wen_a11 = {1'b0, 1'b0};
                            wen_a10 = {1'b0, 1'b0};
                            wen_a9  = {1'b0, 1'b0};
                            wen_a8  = {1'b0, 1'b0};
                            wen_a7  = {1'b0, 1'b0};
                            wen_a6  = {1'b0, 1'b0};
                            wen_a5  = {1'b0, 1'b0};
                            wen_a4  = {1'b0, 1'b0};
                            wen_a3  = {1'b0, 1'b0};    
                            wen_a2  = {1'b0, 1'b0};
                            wen_a1  = {1'b0, 1'b0};
                    end
                         7'b0100000, 7'b0100001, 7'b0100010, 7'b0100011,
                         7'b0100100, 7'b0100101, 7'b0100110, 7'b0100111,
                         7'b0101000, 7'b0101001, 7'b0101010, 7'b0101011,
                         7'b0101100, 7'b0101101, 7'b0101110, 7'b0101111,
                         7'b0110000, 7'b0110001, 7'b0110010, 7'b0110011,
                         7'b0110100, 7'b0110101, 7'b0110110, 7'b0110111,             
                         7'b0111000, 7'b0111001, 7'b0111010, 7'b0111011,
                         7'b0111100, 7'b0111101, 7'b0111110, 7'b0111111  : begin
                            wen_a66 = {1'b0, 1'b0};
                            wen_a65 = {1'b0, 1'b0};
                            wen_a64 = {1'b0, 1'b0};
                            wen_a63 = {1'b0, 1'b0};
                            wen_a62 = {1'b0, 1'b0};
                            wen_a61 = {1'b0, 1'b0};
                            wen_a60 = {1'b0, 1'b0};
                            wen_a59 = {1'b0, 1'b0};
                            wen_a58 = {1'b0, 1'b0};
                            wen_a57 = {1'b0, 1'b0};
                            wen_a56 = {1'b0, 1'b0};
                            wen_a55 = {1'b0, 1'b0};
                            wen_a54 = {1'b0, 1'b0};
                            wen_a53 = {1'b0, 1'b0};
                            wen_a52 = {1'b0, 1'b0};
                            wen_a51 = {1'b0, 1'b0};
                            wen_a50 = {1'b0, 1'b0};
                            wen_a49 = {1'b0, 1'b0};
                            wen_a48 = {1'b0, 1'b0};
                            wen_a47 = {1'b0, 1'b0};
                            wen_a46 = {1'b0, 1'b0};
                            wen_a45 = {1'b0, 1'b0};
                            wen_a44 = {1'b0, 1'b0};
                            wen_a43 = {1'b0, 1'b0};
                            wen_a42 = {1'b0, 1'b0};
                            wen_a41 = {1'b0, 1'b0};
                            wen_a40 = {1'b0, 1'b0};
                            wen_a39 = {1'b0, 1'b0};
                            wen_a38 = {1'b0, 1'b0};
                            wen_a37 = {1'b0, 1'b0};
                            wen_a36 = {1'b0, 1'b0};
                            wen_a35 = {1'b0, 1'b0};
                            wen_a34 = {1'b0, wen};
                            wen_a33 = {1'b0, wen};
                            wen_a32 = {1'b0, wen};
                            wen_a31 = {1'b0, wen};
                            wen_a30 = {1'b0, wen};
                            wen_a29 = {1'b0, wen};
                            wen_a28 = {1'b0, wen};
                            wen_a27 = {1'b0, wen};
                            wen_a26 = {1'b0, wen};
                            wen_a25 = {1'b0, wen};
                            wen_a24 = {1'b0, wen};
                            wen_a23 = {1'b0, wen};
                            wen_a22 = {1'b0, wen};
                            wen_a21 = {1'b0, wen};
                            wen_a20 = {1'b0, wen};
                            wen_a19 = {1'b0, wen};
                            wen_a18 = {1'b0, wen};
                            wen_a17 = {1'b0, wen};
                            wen_a16 = {1'b0, wen};
                            wen_a15 = {1'b0, wen};
                            wen_a14 = {1'b0, wen};
                            wen_a13 = {1'b0, wen};
                            wen_a12 = {1'b0, wen};
                            wen_a11 = {1'b0, wen};
                            wen_a10 = {1'b0, wen};
                            wen_a9  = {1'b0, wen};
                            wen_a8  = {1'b0, wen};
                            wen_a7  = {1'b0, wen};
                            wen_a6  = {1'b0, wen};
                            wen_a5  = {1'b0, wen};
                            wen_a4  = {1'b0, wen};
                            wen_a3  = {1'b0, wen};
                            wen_a2  = {1'b0, 1'b0};
                            wen_a1  = {1'b0, 1'b0};
                    end
                    7'b1000000, 7'b1000001 : begin
                        wen_a66 = {1'b0, 1'b0};
                        wen_a65 = {1'b0, 1'b0};
                        wen_a64 = {1'b0, 1'b0};
                        wen_a63 = {1'b0, 1'b0};
                        wen_a62 = {1'b0, 1'b0};
                        wen_a61 = {1'b0, 1'b0};
                        wen_a60 = {1'b0, 1'b0};
                        wen_a59 = {1'b0, 1'b0};
                        wen_a58 = {1'b0, 1'b0};
                        wen_a57 = {1'b0, 1'b0};
                        wen_a56 = {1'b0, 1'b0};
                        wen_a55 = {1'b0, 1'b0};
                        wen_a54 = {1'b0, 1'b0};
                        wen_a53 = {1'b0, 1'b0};
                        wen_a52 = {1'b0, 1'b0};
                        wen_a51 = {1'b0, 1'b0};
                        wen_a50 = {1'b0, 1'b0};
                        wen_a49 = {1'b0, 1'b0};
                        wen_a48 = {1'b0, 1'b0};
                        wen_a47 = {1'b0, 1'b0};
                        wen_a46 = {1'b0, 1'b0};
                        wen_a45 = {1'b0, 1'b0};
                        wen_a44 = {1'b0, 1'b0};
                        wen_a43 = {1'b0, 1'b0};
                        wen_a42 = {1'b0, 1'b0};
                        wen_a41 = {1'b0, 1'b0};
                        wen_a40 = {1'b0, 1'b0};
                        wen_a39 = {1'b0, 1'b0};
                        wen_a38 = {1'b0, 1'b0};
                        wen_a37 = {1'b0, 1'b0};
                        wen_a36 = {1'b0, 1'b0};
                        wen_a35 = {1'b0, 1'b0};
                        wen_a34 = {1'b0, 1'b0};
                        wen_a33 = {1'b0, 1'b0};
                        wen_a32 = {1'b0, 1'b0};
                        wen_a31 = {1'b0, 1'b0};
                        wen_a30 = {1'b0, 1'b0};
                        wen_a29 = {1'b0, 1'b0};
                        wen_a28 = {1'b0, 1'b0};
                        wen_a27 = {1'b0, 1'b0};
                        wen_a26 = {1'b0, 1'b0};
                        wen_a25 = {1'b0, 1'b0};
                        wen_a24 = {1'b0, 1'b0};
                        wen_a23 = {1'b0, 1'b0};
                        wen_a22 = {1'b0, 1'b0};
                        wen_a21 = {1'b0, 1'b0};
                        wen_a20 = {1'b0, 1'b0};
                        wen_a19 = {1'b0, 1'b0};
                        wen_a18 = {1'b0, 1'b0};
                        wen_a17 = {1'b0, 1'b0};
                        wen_a16 = {1'b0, 1'b0};
                        wen_a15 = {1'b0, 1'b0};
                        wen_a14 = {1'b0, 1'b0};
                        wen_a13 = {1'b0, 1'b0};
                        wen_a12 = {1'b0, 1'b0};
                        wen_a11 = {1'b0, 1'b0};
                        wen_a10 = {1'b0, 1'b0};
                        wen_a9 = {1'b0, 1'b0};
                        wen_a8 = {1'b0, 1'b0};
                        wen_a7 = {1'b0, 1'b0};
                        wen_a6 = {1'b0, 1'b0};
                        wen_a5 = {1'b0, 1'b0};
                        wen_a4 = {1'b0, 1'b0};
                        wen_a3 = {1'b0, 1'b0};
                        wen_a2 = {wen, wen};
                        wen_a1 = {wen, wen};
                    end
                    default : begin
                        wen_a66 = {1'b0, 1'b0};
                        wen_a65 = {1'b0, 1'b0};
                        wen_a64 = {1'b0, 1'b0};
                        wen_a63 = {1'b0, 1'b0};
                        wen_a62 = {1'b0, 1'b0};
                        wen_a61 = {1'b0, 1'b0};
                        wen_a60 = {1'b0, 1'b0};
                        wen_a59 = {1'b0, 1'b0};
                        wen_a58 = {1'b0, 1'b0};
                        wen_a57 = {1'b0, 1'b0};
                        wen_a56 = {1'b0, 1'b0};
                        wen_a55 = {1'b0, 1'b0};
                        wen_a54 = {1'b0, 1'b0};
                        wen_a53 = {1'b0, 1'b0};
                        wen_a52 = {1'b0, 1'b0};
                        wen_a51 = {1'b0, 1'b0};
                        wen_a50 = {1'b0, 1'b0};
                        wen_a49 = {1'b0, 1'b0};
                        wen_a48 = {1'b0, 1'b0};
                        wen_a47 = {1'b0, 1'b0};
                        wen_a46 = {1'b0, 1'b0};
                        wen_a45 = {1'b0, 1'b0};
                        wen_a44 = {1'b0, 1'b0};
                        wen_a43 = {1'b0, 1'b0};
                        wen_a42 = {1'b0, 1'b0};
                        wen_a41 = {1'b0, 1'b0};
                        wen_a40 = {1'b0, 1'b0};
                        wen_a39 = {1'b0, 1'b0};
                        wen_a38 = {1'b0, 1'b0};
                        wen_a37 = {1'b0, 1'b0};
                        wen_a36 = {1'b0, 1'b0};
                        wen_a35 = {1'b0, 1'b0};
                        wen_a34 = {1'b0, 1'b0};
                        wen_a33 = {1'b0, 1'b0};
                        wen_a32 = {1'b0, 1'b0};
                        wen_a31 = {1'b0, 1'b0};
                        wen_a30 = {1'b0, 1'b0};
                        wen_a29 = {1'b0, 1'b0};
                        wen_a28 = {1'b0, 1'b0};
                        wen_a27 = {1'b0, 1'b0};
                        wen_a26 = {1'b0, 1'b0};
                        wen_a25 = {1'b0, 1'b0};
                        wen_a24 = {1'b0, 1'b0};
                        wen_a23 = {1'b0, 1'b0};
                        wen_a22 = {1'b0, 1'b0};
                        wen_a21 = {1'b0, 1'b0};
                        wen_a20 = {1'b0, 1'b0};
                        wen_a19 = {1'b0, 1'b0};
                        wen_a18 = {1'b0, 1'b0};
                        wen_a17 = {1'b0, 1'b0};
                        wen_a16 = {1'b0, 1'b0};
                        wen_a15 = {1'b0, 1'b0};
                        wen_a14 = {1'b0, 1'b0};
                        wen_a13 = {1'b0, 1'b0};
                        wen_a12 = {1'b0, 1'b0};
                        wen_a11 = {1'b0, 1'b0};
                        wen_a10 = {1'b0, 1'b0};
                        wen_a9 = {1'b0, 1'b0};
                        wen_a8 = {1'b0, 1'b0};
                        wen_a7 = {1'b0, 1'b0};
                        wen_a6 = {1'b0, 1'b0};
                        wen_a5 = {1'b0, 1'b0};
                        wen_a4 = {1'b0, 1'b0};
                        wen_a3 = {1'b0, 1'b0};
                        wen_a2 = {1'b0, 1'b0};
                        wen_a1 = {1'b0, 1'b0};
                    end
               endcase // case (writeAddr[15:9])

                case (ckRdAddr[15:9])

                       7'b0000000, 7'b0000001, 7'b0000010, 7'b0000011,
                         7'b0000100, 7'b0000101, 7'b0000110, 7'b0000111,
                         7'b0001000, 7'b0001001, 7'b0001010, 7'b0001011,
                         7'b0001100, 7'b0001101, 7'b0001110, 7'b0001111,
                         7'b0010000, 7'b0010001, 7'b0010010, 7'b0010011,
                         7'b0010100, 7'b0010101, 7'b0010110, 7'b0010111,
                         7'b0011000, 7'b0011001, 7'b0011010, 7'b0011011,
                         7'b0011100, 7'b0011101, 7'b0011110, 7'b0011111 : begin

                        readData = {
                                        readData66[0],
                                        readData65[0],
                                        readData64[0],
                                        readData63[0],
                                        readData62[0],
                                        readData61[0],
                                        readData60[0],
                                        readData59[0],
                                        readData58[0],
                                        readData57[0],
                                        readData56[0],
                                        readData55[0], 
                                        readData54[0],
                                        readData53[0],
                                        readData52[0],
                                        readData51[0],
                                        readData50[0],
                                        readData49[0],
                                        readData48[0],
                                        readData47[0],
                                        readData46[0],
                                        readData45[0],
                                        readData44[0],
                                        readData43[0],
                                        readData42[0],
                                        readData41[0],
                                        readData40[0],
                                        readData39[0],
                                        readData38[0],
                                        readData37[0],
                                        readData36[0],
                                        readData35[0]
                        };
                    end
                  7'b0100000, 7'b0100001, 7'b0100010, 7'b0100011,
                    7'b0100100, 7'b0100101, 7'b0100110, 7'b0100111,
                    7'b0101000, 7'b0101001, 7'b0101010, 7'b0101011,
                    7'b0101100, 7'b0101101, 7'b0101110, 7'b0101111,
                    7'b0110000, 7'b0110001, 7'b0110010, 7'b0110011,
                    7'b0110100, 7'b0110101, 7'b0110110, 7'b0110111,             
                    7'b0111000, 7'b0111001, 7'b0111010, 7'b0111011,
                    7'b0111100, 7'b0111101, 7'b0111110, 7'b0111111  : begin
                        readData = {
                                        readData34[0],
                                        readData33[0],
                                        readData32[0],
                                        readData31[0],
                                        readData30[0],
                                        readData29[0],
                                        readData28[0],
                                        readData27[0],
                                        readData26[0],
                                        readData25[0],
                                        readData24[0],
                                        readData23[0],
                                        readData22[0],
                                        readData21[0],
                                        readData20[0],
                                        readData19[0],
                                        readData18[0],
                                        readData17[0],
                                        readData16[0],
                                        readData15[0],
                                        readData14[0],
                                        readData13[0],
                                        readData12[0],
                                        readData11[0],
                                        readData10[0],
                                        readData9[0],
                                        readData8[0],
                                        readData7[0],
                                        readData6[0],
                                        readData5[0],
                                        readData4[0],
                                        readData3[0]
                                    };                       
                    end                            
                    7'b1000000, 7'b1000001 : begin
                        readData = {readData2[16:9],readData2[7:0],readData1[16:9],readData1[7:0]};
                    end
                    default : begin
                        readData = 32'b0;
                    end
                endcase
          end // case: 33792
          34304: begin
                     width66 = 3'b000;
                     width65 = 3'b000;
                     width64 = 3'b000;
                     width63 = 3'b000;
                     width62 = 3'b000;
                     width61 = 3'b000;
                     width60 = 3'b000;
                     width59 = 3'b000;
                     width58 = 3'b000;
                     width57 = 3'b000;
                     width56 = 3'b000;
                     width55 = 3'b000;
                     width54 = 3'b000;
                     width53 = 3'b000;
                     width52 = 3'b000;
                     width51 = 3'b000;
                     width50 = 3'b000;
                     width49 = 3'b000;
                     width48 = 3'b000;
                     width47 = 3'b000;
                     width46 = 3'b000;
                     width45 = 3'b000;
                     width44 = 3'b000;
                     width43 = 3'b000;
                     width42 = 3'b000;
                     width41 = 3'b000;
                     width40 = 3'b000;
                     width39 = 3'b000;
                     width38 = 3'b000;
                     width37 = 3'b000;
                     width36 = 3'b000;
                     width35 = 3'b000;
                     width34 = 3'b000;
                     width33 = 3'b000;
                     width32 = 3'b000;
                     width31 = 3'b000;
                     width30 = 3'b000;
                     width29 = 3'b000;
                     width28 = 3'b000;
                     width27 = 3'b000;
                     width26 = 3'b000;
                     width25 = 3'b000;
                     width24 = 3'b000;
                     width23 = 3'b000;
                     width22 = 3'b000;
                     width21 = 3'b000;
                     width20 = 3'b000;
                     width19 = 3'b000;
                     width18 = 3'b000;
                     width17 = 3'b000;
                     width16 = 3'b000;
                     width15 = 3'b000;
                     width14 = 3'b000;
                     width13 = 3'b000;
                     width12 = 3'b000;
                     width11 = 3'b000;
                     width10 = 3'b000;
                     width9 = 3'b000;
                     width8 = 3'b000;
                     width7 = 3'b000;
                     width6 = 3'b000;
                     width5 = 3'b000;
                     width4 = 3'b000;
                     width3 = 3'b000;
                     width2 = 3'b100;
                     width1 = 3'b100;
                     width0 = 3'b101;
                                    
                    writeAddr66 = {writeAddr[13:0]};
                    writeAddr65 = {writeAddr[13:0]};
                    writeAddr64 = {writeAddr[13:0]};
                    writeAddr63 = {writeAddr[13:0]};
                    writeAddr62 = {writeAddr[13:0]};
                    writeAddr61 = {writeAddr[13:0]};
                    writeAddr60 = {writeAddr[13:0]};
                    writeAddr59 = {writeAddr[13:0]};
                    writeAddr58 = {writeAddr[13:0]};
                    writeAddr57 = {writeAddr[13:0]};
                    writeAddr56 = {writeAddr[13:0]};
                    writeAddr55 = {writeAddr[13:0]};
                    writeAddr54 = {writeAddr[13:0]};
                    writeAddr53 = {writeAddr[13:0]};
                    writeAddr52 = {writeAddr[13:0]};
                    writeAddr51 = {writeAddr[13:0]};
                    writeAddr50 = {writeAddr[13:0]};
                    writeAddr49 = {writeAddr[13:0]};
                    writeAddr48 = {writeAddr[13:0]};
                    writeAddr47 = {writeAddr[13:0]};
                    writeAddr46 = {writeAddr[13:0]};
                    writeAddr45 = {writeAddr[13:0]};
                    writeAddr44 = {writeAddr[13:0]};
                    writeAddr43 = {writeAddr[13:0]};
                    writeAddr42 = {writeAddr[13:0]};
                    writeAddr41 = {writeAddr[13:0]};
                    writeAddr40 = {writeAddr[13:0]};
                    writeAddr39 = {writeAddr[13:0]};
                    writeAddr38 = {writeAddr[13:0]};
                    writeAddr37 = {writeAddr[13:0]};
                    writeAddr36 = {writeAddr[13:0]};
                    writeAddr35 = {writeAddr[13:0]};
                    writeAddr34 = {writeAddr[13:0]};
                    writeAddr33 = {writeAddr[13:0]};
                    writeAddr32 = {writeAddr[13:0]};
                    writeAddr31 = {writeAddr[13:0]};
                    writeAddr30 = {writeAddr[13:0]};
                    writeAddr29 = {writeAddr[13:0]};
                    writeAddr28 = {writeAddr[13:0]};
                    writeAddr27 = {writeAddr[13:0]};
                    writeAddr26 = {writeAddr[13:0]};
                    writeAddr25 = {writeAddr[13:0]};
                    writeAddr24 = {writeAddr[13:0]};
                    writeAddr23 = {writeAddr[13:0]};
                    writeAddr22 = {writeAddr[13:0]};
                    writeAddr21 = {writeAddr[13:0]};
                    writeAddr20 = {writeAddr[13:0]};
                    writeAddr19 = {writeAddr[13:0]};
                    writeAddr18 = {writeAddr[13:0]};
                    writeAddr17 = {writeAddr[13:0]};
                    writeAddr16 = {writeAddr[13:0]};
                    writeAddr15 = {writeAddr[13:0]};
                    writeAddr14 = {writeAddr[13:0]};
                    writeAddr13 = {writeAddr[13:0]};
                    writeAddr12 = {writeAddr[13:0]};
                    writeAddr11 = {writeAddr[13:0]};
                    writeAddr10 = {writeAddr[13:0]};
                    writeAddr9 = {writeAddr[13:0]};
                    writeAddr8 = {writeAddr[13:0]};
                    writeAddr7 = {writeAddr[13:0]};
                    writeAddr6 = {writeAddr[13:0]};
                    writeAddr5 = {writeAddr[13:0]};
                    writeAddr4 = {writeAddr[13:0]};
             writeAddr3 = {writeAddr[13:0]};
             writeAddr2 = {writeAddr[9:0], 4'b0};
             writeAddr1 = {writeAddr[9:0], 4'b0};
             writeAddr0 = {writeAddr[8:0], 5'b0};

                    readAddr66 = {readAddr[13:0]};                         
                    readAddr65 = {readAddr[13:0]};
                    readAddr64 = {readAddr[13:0]};
                    readAddr63 = {readAddr[13:0]};
                    readAddr62 = {readAddr[13:0]};
                    readAddr61 = {readAddr[13:0]};
                    readAddr60 = {readAddr[13:0]};
                    readAddr59 = {readAddr[13:0]};
                    readAddr58 = {readAddr[13:0]};
                    readAddr57 = {readAddr[13:0]};
                    readAddr56 = {readAddr[13:0]};
                    readAddr55 = {readAddr[13:0]};
                    readAddr54 = {readAddr[13:0]};
                    readAddr53 = {readAddr[13:0]};
                    readAddr52 = {readAddr[13:0]};
                    readAddr51 = {readAddr[13:0]};
                    readAddr50 = {readAddr[13:0]};
                    readAddr49 = {readAddr[13:0]};
                    readAddr48 = {readAddr[13:0]};
                    readAddr47 = {readAddr[13:0]};
                    readAddr46 = {readAddr[13:0]};
                    readAddr45 = {readAddr[13:0]};
                    readAddr44 = {readAddr[13:0]};
                    readAddr43 = {readAddr[13:0]};
                    readAddr42 = {readAddr[13:0]};
                    readAddr41 = {readAddr[13:0]};
                    readAddr40 = {readAddr[13:0]};
                    readAddr39 = {readAddr[13:0]};
                    readAddr38 = {readAddr[13:0]};
                    readAddr37 = {readAddr[13:0]};
                    readAddr36 = {readAddr[13:0]};
                    readAddr35 = {readAddr[13:0]};
                    readAddr34 = {readAddr[13:0]};
                    readAddr33 = {readAddr[13:0]};
                    readAddr32 = {readAddr[13:0]};
                    readAddr31 = {readAddr[13:0]};
                    readAddr30 = {readAddr[13:0]};
                    readAddr29 = {readAddr[13:0]};
                    readAddr28 = {readAddr[13:0]};
                    readAddr27 = {readAddr[13:0]};
                    readAddr26 = {readAddr[13:0]};
                    readAddr25 = {readAddr[13:0]};
                    readAddr24 = {readAddr[13:0]};
                    readAddr23 = {readAddr[13:0]};
                    readAddr22 = {readAddr[13:0]};
                    readAddr21 = {readAddr[13:0]};
                    readAddr20 = {readAddr[13:0]};
                    readAddr19 = {readAddr[13:0]};
                    readAddr18 = {readAddr[13:0]};
                    readAddr17 = {readAddr[13:0]};
                    readAddr16 = {readAddr[13:0]};
                    readAddr15 = {readAddr[13:0]};
                    readAddr14 = {readAddr[13:0]};
                    readAddr13 = {readAddr[13:0]};
                    readAddr12 = {readAddr[13:0]};
                    readAddr11 = {readAddr[13:0]};
                    readAddr10 = {readAddr[13:0]};
                    readAddr9 = {readAddr[13:0]};
                    readAddr8 = {readAddr[13:0]};
                    readAddr7 = {readAddr[13:0]};
                    readAddr6 = {readAddr[13:0]};
                    readAddr5 = {readAddr[13:0]};
                    readAddr4 = {readAddr[13:0]};
                    readAddr3 = {readAddr[13:0]};
                    readAddr2  = {readAddr[9:0],  4'b0};
                    readAddr1  = {readAddr[9:0],  4'b0};
                    readAddr0  = {readAddr[8:0],  5'b0};
                     

                     writeData66 = {17'b0, writeData[31]};
                     writeData65 = {17'b0, writeData[30]};
                     writeData64 = {17'b0, writeData[29]};
                     writeData63 = {17'b0, writeData[28]};
                     writeData62 = {17'b0, writeData[27]};
                     writeData61 = {17'b0, writeData[26]};
                     writeData60 = {17'b0, writeData[25]};
                     writeData59 = {17'b0, writeData[24]};
                     writeData58 = {17'b0, writeData[23]};
                     writeData57 = {17'b0, writeData[22]};
                     writeData56 = {17'b0, writeData[21]};
                     writeData55 = {17'b0, writeData[20]};
                     writeData54 = {17'b0, writeData[19]};
                     writeData53 = {17'b0, writeData[18]};
                     writeData52 = {17'b0, writeData[17]};
                     writeData51 = {17'b0, writeData[16]};
                     writeData50 = {17'b0, writeData[15]};
                     writeData49 = {17'b0, writeData[14]};
                     writeData48 = {17'b0, writeData[13]};
                     writeData47 = {17'b0, writeData[12]};
                     writeData46 = {17'b0, writeData[11]};
                     writeData45 = {17'b0, writeData[10]};
                     writeData44 = {17'b0, writeData[9]};
                     writeData43 = {17'b0, writeData[8]};
                     writeData42 = {17'b0, writeData[7]};
                     writeData41 = {17'b0, writeData[6]};
                     writeData40 = {17'b0, writeData[5]};
                     writeData39 = {17'b0, writeData[4]};
                     writeData38 = {17'b0, writeData[3]};
                     writeData37 = {17'b0, writeData[2]};
                     writeData36 = {17'b0, writeData[1]};
                     writeData35 = {17'b0, writeData[0]};
                     writeData34 = {17'b0, writeData[31]};
                     writeData33 = {17'b0, writeData[30]};
                     writeData32 = {17'b0, writeData[29]};
                     writeData31 = {17'b0, writeData[28]};
                     writeData30 = {17'b0, writeData[27]};
                     writeData29 = {17'b0, writeData[26]};
                     writeData28 = {17'b0, writeData[25]};
                     writeData27 = {17'b0, writeData[24]};
                     writeData26 = {17'b0, writeData[23]};
                     writeData25 = {17'b0, writeData[22]};
                     writeData24 = {17'b0, writeData[21]};
                     writeData23 = {17'b0, writeData[20]};
                     writeData22 = {17'b0, writeData[19]};
                     writeData21 = {17'b0, writeData[18]};
                     writeData20 = {17'b0, writeData[17]};
                     writeData19 = {17'b0, writeData[16]};
                     writeData18 = {17'b0, writeData[15]};
                     writeData17 = {17'b0, writeData[14]};
                     writeData16 = {17'b0, writeData[13]};
                     writeData15 = {17'b0, writeData[12]};
                     writeData14 = {17'b0, writeData[11]};
                     writeData13 = {17'b0, writeData[10]};
                     writeData12 = {17'b0, writeData[9]};
                     writeData11 = {17'b0, writeData[8]};
                     writeData10 = {17'b0, writeData[7]};
                     writeData9 = {17'b0, writeData[6]};
                     writeData8 = {17'b0, writeData[5]};
                     writeData7 = {17'b0, writeData[4]};
                     writeData6 = {17'b0, writeData[3]};
                     writeData5 = {17'b0, writeData[2]};
                     writeData4 = {17'b0, writeData[1]};
                     writeData3 = {17'b0, writeData[0]};
                writeData2 = {1'b0, writeData[31:24], 1'b0, writeData[23:16]};
                writeData1 = {1'b0, writeData[15:8], 1'b0, writeData[7:0]};
                writeData0 = {1'b0, writeData[31:24], 1'b0, writeData[23:16], 1'b0, writeData[15:8], 1'b0, writeData[7:0]};


                case (writeAddr[15:9])
                       7'b0000000, 7'b0000001, 7'b0000010, 7'b0000011,
                         7'b0000100, 7'b0000101, 7'b0000110, 7'b0000111,
                         7'b0001000, 7'b0001001, 7'b0001010, 7'b0001011,
                         7'b0001100, 7'b0001101, 7'b0001110, 7'b0001111,
                         7'b0010000, 7'b0010001, 7'b0010010, 7'b0010011,
                         7'b0010100, 7'b0010101, 7'b0010110, 7'b0010111,
                         7'b0011000, 7'b0011001, 7'b0011010, 7'b0011011,
                         7'b0011100, 7'b0011101, 7'b0011110, 7'b0011111 : begin
                            wen_a66 = {1'b0, wen};
                            wen_a65 = {1'b0, wen};
                            wen_a64 = {1'b0, wen};
                            wen_a63 = {1'b0, wen};
                            wen_a62 = {1'b0, wen};
                            wen_a61 = {1'b0, wen};
                            wen_a60 = {1'b0, wen};
                            wen_a59 = {1'b0, wen};
                            wen_a58 = {1'b0, wen};
                            wen_a57 = {1'b0, wen};
                            wen_a56 = {1'b0, wen};
                            wen_a55 = {1'b0, wen};
                            wen_a54 = {1'b0, wen};
                            wen_a53 = {1'b0, wen};
                            wen_a52 = {1'b0, wen};
                            wen_a51 = {1'b0, wen};
                            wen_a50 = {1'b0, wen};
                            wen_a49 = {1'b0, wen};
                            wen_a48 = {1'b0, wen};
                            wen_a47 = {1'b0, wen};
                            wen_a46 = {1'b0, wen};
                            wen_a45 = {1'b0, wen};
                            wen_a44 = {1'b0, wen};
                            wen_a43 = {1'b0, wen};
                            wen_a42 = {1'b0, wen};
                            wen_a41 = {1'b0, wen};
                            wen_a40 = {1'b0, wen};
                            wen_a39 = {1'b0, wen};
                            wen_a38 = {1'b0, wen};
                            wen_a37 = {1'b0, wen};
                            wen_a36 = {1'b0, wen};
                            wen_a35 = {1'b0, wen};
                            wen_a34 = {1'b0, 1'b0};
                            wen_a33 = {1'b0, 1'b0};
                            wen_a32 = {1'b0, 1'b0};
                            wen_a31 = {1'b0, 1'b0};
                            wen_a30 = {1'b0, 1'b0};
                            wen_a29 = {1'b0, 1'b0};
                            wen_a28 = {1'b0, 1'b0};
                            wen_a27 = {1'b0, 1'b0};
                            wen_a26 = {1'b0, 1'b0};
                            wen_a25 = {1'b0, 1'b0};
                            wen_a24 = {1'b0, 1'b0};
                            wen_a23 = {1'b0, 1'b0};
                            wen_a22 = {1'b0, 1'b0};
                            wen_a21 = {1'b0, 1'b0};
                            wen_a20 = {1'b0, 1'b0};
                            wen_a19 = {1'b0, 1'b0};
                            wen_a18 = {1'b0, 1'b0};
                            wen_a17 = {1'b0, 1'b0};
                            wen_a16 = {1'b0, 1'b0};
                            wen_a15 = {1'b0, 1'b0};
                            wen_a14 = {1'b0, 1'b0};
                            wen_a13 = {1'b0, 1'b0};
                            wen_a12 = {1'b0, 1'b0};
                            wen_a11 = {1'b0, 1'b0};
                            wen_a10 = {1'b0, 1'b0};
                            wen_a9  = {1'b0, 1'b0};
                            wen_a8  = {1'b0, 1'b0};
                            wen_a7  = {1'b0, 1'b0};
                            wen_a6  = {1'b0, 1'b0};
                            wen_a5  = {1'b0, 1'b0};
                            wen_a4  = {1'b0, 1'b0};
                            wen_a3  = {1'b0, 1'b0};
                            wen_a2  = {1'b0, 1'b0};
                            wen_a1  = {1'b0, 1'b0};
                            wen_a0  = {1'b0, 1'b0};
                            wen_b0  = {1'b0, 1'b0};

                    end
                         7'b0100000, 7'b0100001, 7'b0100010, 7'b0100011,
                         7'b0100100, 7'b0100101, 7'b0100110, 7'b0100111,
                         7'b0101000, 7'b0101001, 7'b0101010, 7'b0101011,
                         7'b0101100, 7'b0101101, 7'b0101110, 7'b0101111,
                         7'b0110000, 7'b0110001, 7'b0110010, 7'b0110011,
                         7'b0110100, 7'b0110101, 7'b0110110, 7'b0110111,             
                         7'b0111000, 7'b0111001, 7'b0111010, 7'b0111011,
                         7'b0111100, 7'b0111101, 7'b0111110, 7'b0111111  : begin
                            wen_a66 = {1'b0, 1'b0};
                            wen_a65 = {1'b0, 1'b0};
                            wen_a64 = {1'b0, 1'b0};
                            wen_a63 = {1'b0, 1'b0};
                            wen_a62 = {1'b0, 1'b0};
                            wen_a61 = {1'b0, 1'b0};
                            wen_a60 = {1'b0, 1'b0};
                            wen_a59 = {1'b0, 1'b0};
                            wen_a58 = {1'b0, 1'b0};
                            wen_a57 = {1'b0, 1'b0};
                            wen_a56 = {1'b0, 1'b0};
                            wen_a55 = {1'b0, 1'b0};
                            wen_a54 = {1'b0, 1'b0};
                            wen_a53 = {1'b0, 1'b0};
                            wen_a52 = {1'b0, 1'b0};
                            wen_a51 = {1'b0, 1'b0};
                            wen_a50 = {1'b0, 1'b0};
                            wen_a49 = {1'b0, 1'b0};
                            wen_a48 = {1'b0, 1'b0};
                            wen_a47 = {1'b0, 1'b0};
                            wen_a46 = {1'b0, 1'b0};
                            wen_a45 = {1'b0, 1'b0};
                            wen_a44 = {1'b0, 1'b0};
                            wen_a43 = {1'b0, 1'b0};
                            wen_a42 = {1'b0, 1'b0};
                            wen_a41 = {1'b0, 1'b0};
                            wen_a40 = {1'b0, 1'b0};
                            wen_a39 = {1'b0, 1'b0};
                            wen_a38 = {1'b0, 1'b0};
                            wen_a37 = {1'b0, 1'b0};
                            wen_a36 = {1'b0, 1'b0};
                            wen_a35 = {1'b0, 1'b0};
                            wen_a34 = {1'b0, wen};
                            wen_a33 = {1'b0, wen};
                            wen_a32 = {1'b0, wen};
                            wen_a31 = {1'b0, wen};
                            wen_a30 = {1'b0, wen};
                            wen_a29 = {1'b0, wen};
                            wen_a28 = {1'b0, wen};
                            wen_a27 = {1'b0, wen};
                            wen_a26 = {1'b0, wen};
                            wen_a25 = {1'b0, wen};
                            wen_a24 = {1'b0, wen};
                            wen_a23 = {1'b0, wen};
                            wen_a22 = {1'b0, wen};
                            wen_a21 = {1'b0, wen};
                            wen_a20 = {1'b0, wen};
                            wen_a19 = {1'b0, wen};
                            wen_a18 = {1'b0, wen};
                            wen_a17 = {1'b0, wen};
                            wen_a16 = {1'b0, wen};
                            wen_a15 = {1'b0, wen};
                            wen_a14 = {1'b0, wen};
                            wen_a13 = {1'b0, wen};
                            wen_a12 = {1'b0, wen};
                            wen_a11 = {1'b0, wen};
                            wen_a10 = {1'b0, wen};
                            wen_a9  = {1'b0, wen};
                            wen_a8  = {1'b0, wen};
                            wen_a7  = {1'b0, wen};
                            wen_a6  = {1'b0, wen};
                            wen_a5  = {1'b0, wen};
                            wen_a4  = {1'b0, wen};
                            wen_a3  = {1'b0, wen};
                            wen_a2  = {1'b0, 1'b0};
                            wen_a1  = {1'b0, 1'b0};
                            wen_a0  = {1'b0, 1'b0};
                            wen_b0  = {1'b0, 1'b0};

                    end

                    7'b1000000, 7'b1000001 : begin
                        wen_a66 = {1'b0, 1'b0};
                        wen_a65 = {1'b0, 1'b0};
                        wen_a64 = {1'b0, 1'b0};
                        wen_a63 = {1'b0, 1'b0};
                        wen_a62 = {1'b0, 1'b0};
                        wen_a61 = {1'b0, 1'b0};
                        wen_a60 = {1'b0, 1'b0};
                        wen_a59 = {1'b0, 1'b0};
                        wen_a58 = {1'b0, 1'b0};
                        wen_a57 = {1'b0, 1'b0};
                        wen_a56 = {1'b0, 1'b0};
                        wen_a55 = {1'b0, 1'b0};
                        wen_a54 = {1'b0, 1'b0};
                        wen_a53 = {1'b0, 1'b0};
                        wen_a52 = {1'b0, 1'b0};
                        wen_a51 = {1'b0, 1'b0};
                        wen_a50 = {1'b0, 1'b0};
                        wen_a49 = {1'b0, 1'b0};
                        wen_a48 = {1'b0, 1'b0};
                        wen_a47 = {1'b0, 1'b0};
                        wen_a46 = {1'b0, 1'b0};
                        wen_a45 = {1'b0, 1'b0};
                        wen_a44 = {1'b0, 1'b0};
                        wen_a43 = {1'b0, 1'b0};
                        wen_a42 = {1'b0, 1'b0};
                        wen_a41 = {1'b0, 1'b0};
                        wen_a40 = {1'b0, 1'b0};
                        wen_a39 = {1'b0, 1'b0};
                        wen_a38 = {1'b0, 1'b0};
                        wen_a37 = {1'b0, 1'b0};
                        wen_a36 = {1'b0, 1'b0};
                        wen_a35 = {1'b0, 1'b0};
                        wen_a34 = {1'b0, 1'b0};
                        wen_a33 = {1'b0, 1'b0};
                        wen_a32 = {1'b0, 1'b0};
                        wen_a31 = {1'b0, 1'b0};
                        wen_a30 = {1'b0, 1'b0};
                        wen_a29 = {1'b0, 1'b0};
                        wen_a28 = {1'b0, 1'b0};
                        wen_a27 = {1'b0, 1'b0};
                        wen_a26 = {1'b0, 1'b0};
                        wen_a25 = {1'b0, 1'b0};
                        wen_a24 = {1'b0, 1'b0};
                        wen_a23 = {1'b0, 1'b0};
                        wen_a22 = {1'b0, 1'b0};
                        wen_a21 = {1'b0, 1'b0};
                        wen_a20 = {1'b0, 1'b0};
                        wen_a19 = {1'b0, 1'b0};
                        wen_a18 = {1'b0, 1'b0};
                        wen_a17 = {1'b0, 1'b0};
                        wen_a16 = {1'b0, 1'b0};
                        wen_a15 = {1'b0, 1'b0};
                        wen_a14 = {1'b0, 1'b0};
                        wen_a13 = {1'b0, 1'b0};
                        wen_a12 = {1'b0, 1'b0};
                        wen_a11 = {1'b0, 1'b0};
                        wen_a10 = {1'b0, 1'b0};
                        wen_a9 = {1'b0, 1'b0};
                        wen_a8 = {1'b0, 1'b0};
                        wen_a7 = {1'b0, 1'b0};
                        wen_a6 = {1'b0, 1'b0};
                        wen_a5 = {1'b0, 1'b0};
                        wen_a4 = {1'b0, 1'b0};
                        wen_a3 = {1'b0, 1'b0};
                        wen_a2 = {wen, wen};
                        wen_a1 = {wen, wen};
                        wen_a0 = {1'b0, 1'b0};
                        wen_b0 = {1'b0, 1'b0};
                    end
                    7'b1000010 : begin
                        wen_a66 = {1'b0, 1'b0};
                        wen_a65 = {1'b0, 1'b0};
                        wen_a64 = {1'b0, 1'b0};
                        wen_a63 = {1'b0, 1'b0};
                        wen_a62 = {1'b0, 1'b0};
                        wen_a61 = {1'b0, 1'b0};
                        wen_a60 = {1'b0, 1'b0};
                        wen_a59 = {1'b0, 1'b0};
                        wen_a58 = {1'b0, 1'b0};
                        wen_a57 = {1'b0, 1'b0};
                        wen_a56 = {1'b0, 1'b0};
                        wen_a55 = {1'b0, 1'b0};
                        wen_a54 = {1'b0, 1'b0};
                        wen_a53 = {1'b0, 1'b0};
                        wen_a52 = {1'b0, 1'b0};
                        wen_a51 = {1'b0, 1'b0};
                        wen_a50 = {1'b0, 1'b0};
                        wen_a49 = {1'b0, 1'b0};
                        wen_a48 = {1'b0, 1'b0};
                        wen_a47 = {1'b0, 1'b0};
                        wen_a46 = {1'b0, 1'b0};
                        wen_a45 = {1'b0, 1'b0};
                        wen_a44 = {1'b0, 1'b0};
                        wen_a43 = {1'b0, 1'b0};
                        wen_a42 = {1'b0, 1'b0};
                        wen_a41 = {1'b0, 1'b0};
                        wen_a40 = {1'b0, 1'b0};
                        wen_a39 = {1'b0, 1'b0};
                        wen_a38 = {1'b0, 1'b0};
                        wen_a37 = {1'b0, 1'b0};
                        wen_a36 = {1'b0, 1'b0};
                        wen_a35 = {1'b0, 1'b0};
                        wen_a34 = {1'b0, 1'b0};
                        wen_a33 = {1'b0, 1'b0};
                        wen_a32 = {1'b0, 1'b0};
                        wen_a31 = {1'b0, 1'b0};
                        wen_a30 = {1'b0, 1'b0};
                        wen_a29 = {1'b0, 1'b0};
                        wen_a28 = {1'b0, 1'b0};
                        wen_a27 = {1'b0, 1'b0};
                        wen_a26 = {1'b0, 1'b0};
                        wen_a25 = {1'b0, 1'b0};
                        wen_a24 = {1'b0, 1'b0};
                        wen_a23 = {1'b0, 1'b0};
                        wen_a22 = {1'b0, 1'b0};
                        wen_a21 = {1'b0, 1'b0};
                        wen_a20 = {1'b0, 1'b0};
                        wen_a19 = {1'b0, 1'b0};
                        wen_a18 = {1'b0, 1'b0};
                        wen_a17 = {1'b0, 1'b0};
                        wen_a16 = {1'b0, 1'b0};
                        wen_a15 = {1'b0, 1'b0};
                        wen_a14 = {1'b0, 1'b0};
                        wen_a13 = {1'b0, 1'b0};
                        wen_a12 = {1'b0, 1'b0};
                        wen_a11 = {1'b0, 1'b0};
                        wen_a10 = {1'b0, 1'b0};
                        wen_a9 = {1'b0, 1'b0};
                        wen_a8 = {1'b0, 1'b0};
                        wen_a7 = {1'b0, 1'b0};
                        wen_a6 = {1'b0, 1'b0};
                        wen_a5 = {1'b0, 1'b0};
                        wen_a4 = {1'b0, 1'b0};
                        wen_a3 = {1'b0, 1'b0};
                        wen_a2 = {1'b0, 1'b0};
                        wen_a1 = {1'b0, 1'b0};
                        wen_a0 = {wen, wen};
                        wen_b0 = {wen, wen};

                    end
                    default : begin
                        wen_a66 = {1'b0, 1'b0};
                        wen_a65 = {1'b0, 1'b0};
                        wen_a64 = {1'b0, 1'b0};
                        wen_a63 = {1'b0, 1'b0};
                        wen_a62 = {1'b0, 1'b0};
                        wen_a61 = {1'b0, 1'b0};
                        wen_a60 = {1'b0, 1'b0};
                        wen_a59 = {1'b0, 1'b0};
                        wen_a58 = {1'b0, 1'b0};
                        wen_a57 = {1'b0, 1'b0};
                        wen_a56 = {1'b0, 1'b0};
                        wen_a55 = {1'b0, 1'b0};
                        wen_a54 = {1'b0, 1'b0};
                        wen_a53 = {1'b0, 1'b0};
                        wen_a52 = {1'b0, 1'b0};
                        wen_a51 = {1'b0, 1'b0};
                        wen_a50 = {1'b0, 1'b0};
                        wen_a49 = {1'b0, 1'b0};
                        wen_a48 = {1'b0, 1'b0};
                        wen_a47 = {1'b0, 1'b0};
                        wen_a46 = {1'b0, 1'b0};
                        wen_a45 = {1'b0, 1'b0};
                        wen_a44 = {1'b0, 1'b0};
                        wen_a43 = {1'b0, 1'b0};
                        wen_a42 = {1'b0, 1'b0};
                        wen_a41 = {1'b0, 1'b0};
                        wen_a40 = {1'b0, 1'b0};
                        wen_a39 = {1'b0, 1'b0};
                        wen_a38 = {1'b0, 1'b0};
                        wen_a37 = {1'b0, 1'b0};
                        wen_a36 = {1'b0, 1'b0};
                        wen_a35 = {1'b0, 1'b0};
                        wen_a34 = {1'b0, 1'b0};
                        wen_a33 = {1'b0, 1'b0};
                        wen_a32 = {1'b0, 1'b0};
                        wen_a31 = {1'b0, 1'b0};
                        wen_a30 = {1'b0, 1'b0};
                        wen_a29 = {1'b0, 1'b0};
                        wen_a28 = {1'b0, 1'b0};
                        wen_a27 = {1'b0, 1'b0};
                        wen_a26 = {1'b0, 1'b0};
                        wen_a25 = {1'b0, 1'b0};
                        wen_a24 = {1'b0, 1'b0};
                        wen_a23 = {1'b0, 1'b0};
                        wen_a22 = {1'b0, 1'b0};
                        wen_a21 = {1'b0, 1'b0};
                        wen_a20 = {1'b0, 1'b0};
                        wen_a19 = {1'b0, 1'b0};
                        wen_a18 = {1'b0, 1'b0};
                        wen_a17 = {1'b0, 1'b0};
                        wen_a16 = {1'b0, 1'b0};
                        wen_a15 = {1'b0, 1'b0};
                        wen_a14 = {1'b0, 1'b0};
                        wen_a13 = {1'b0, 1'b0};
                        wen_a12 = {1'b0, 1'b0};
                        wen_a11 = {1'b0, 1'b0};
                        wen_a10 = {1'b0, 1'b0};
                        wen_a9 = {1'b0, 1'b0};
                        wen_a8 = {1'b0, 1'b0};
                        wen_a7 = {1'b0, 1'b0};
                        wen_a6 = {1'b0, 1'b0};
                        wen_a5 = {1'b0, 1'b0};
                        wen_a4 = {1'b0, 1'b0};
                        wen_a3 = {1'b0, 1'b0};
                        wen_a2 = {1'b0, 1'b0};
                        wen_a1 = {1'b0, 1'b0};
                        wen_a0 = {1'b0, 1'b0};
                        wen_b0 = {1'b0, 1'b0};
                    end
               endcase // case (writeAddr[15:9])

                case (ckRdAddr[15:9])

                       7'b0000000, 7'b0000001, 7'b0000010, 7'b0000011,
                         7'b0000100, 7'b0000101, 7'b0000110, 7'b0000111,
                         7'b0001000, 7'b0001001, 7'b0001010, 7'b0001011,
                         7'b0001100, 7'b0001101, 7'b0001110, 7'b0001111,
                         7'b0010000, 7'b0010001, 7'b0010010, 7'b0010011,
                         7'b0010100, 7'b0010101, 7'b0010110, 7'b0010111,
                         7'b0011000, 7'b0011001, 7'b0011010, 7'b0011011,
                         7'b0011100, 7'b0011101, 7'b0011110, 7'b0011111 : begin

                        readData = {
                                        readData66[0],
                                        readData65[0],
                                        readData64[0],
                                        readData63[0],
                                        readData62[0],
                                        readData61[0],
                                        readData60[0],
                                        readData59[0],
                                        readData58[0],
                                        readData57[0],
                                        readData56[0],
                                        readData55[0], 
                                        readData54[0],
                                        readData53[0],
                                        readData52[0],
                                        readData51[0],
                                        readData50[0],
                                        readData49[0],
                                        readData48[0],
                                        readData47[0],
                                        readData46[0],
                                        readData45[0],
                                        readData44[0],
                                        readData43[0],
                                        readData42[0],
                                        readData41[0],
                                        readData40[0],
                                        readData39[0],
                                        readData38[0],
                                        readData37[0],
                                        readData36[0],
                                        readData35[0]
                        };
                    end
                    7'b0100000, 7'b0100001, 7'b0100010, 7'b0100011,
                    7'b0100100, 7'b0100101, 7'b0100110, 7'b0100111,
                    7'b0101000, 7'b0101001, 7'b0101010, 7'b0101011,
                    7'b0101100, 7'b0101101, 7'b0101110, 7'b0101111,
                    7'b0110000, 7'b0110001, 7'b0110010, 7'b0110011,
                    7'b0110100, 7'b0110101, 7'b0110110, 7'b0110111,             
                    7'b0111000, 7'b0111001, 7'b0111010, 7'b0111011,
                    7'b0111100, 7'b0111101, 7'b0111110, 7'b0111111  : begin
                        readData = {
                                        readData34[0],
                                        readData33[0],
                                        readData32[0],
                                        readData31[0],
                                        readData30[0],
                                        readData29[0],
                                        readData28[0],
                                        readData27[0],
                                        readData26[0],
                                        readData25[0],
                                        readData24[0],
                                        readData23[0],
                                        readData22[0],
                                        readData21[0],
                                        readData20[0],
                                        readData19[0],
                                        readData18[0],
                                        readData17[0],
                                        readData16[0],
                                        readData15[0],
                                        readData14[0],
                                        readData13[0],
                                        readData12[0],
                                        readData11[0],
                                        readData10[0],
                                        readData9[0],
                                        readData8[0],
                                        readData7[0],
                                        readData6[0],
                                        readData5[0],
                                        readData4[0],
                                        readData3[0]
                                    };                       
                    end                            
                    7'b1000000, 7'b1000001 : begin
                        readData = {readData2[16:9],readData2[7:0],readData1[16:9],readData1[7:0]};
                    end
                    7'b1000010 : begin
                        readData = {readData0[34:27],readData0[25:18],readData0[16:9],readData0[7:0]};
                    end
                    default : begin
                       readData = 32'b0;
                    end
               endcase // case (ckRdAddr[15:9])                                    
            end // case: 34304
          34816: begin
                     width68 = 3'b000;
                     width67 = 3'b000;
                     width66 = 3'b000;
                     width65 = 3'b000;
                     width64 = 3'b000;
                     width63 = 3'b000;
                     width62 = 3'b000;
                     width61 = 3'b000;
                     width60 = 3'b000;
                     width59 = 3'b000;
                     width58 = 3'b000;
                     width57 = 3'b000;
                     width56 = 3'b000;
                     width55 = 3'b000;
                     width54 = 3'b000;
                     width53 = 3'b000;
                     width52 = 3'b000;
                     width51 = 3'b000;
                     width50 = 3'b000;
                     width49 = 3'b000;
                     width48 = 3'b000;
                     width47 = 3'b000;
                     width46 = 3'b000;
                     width45 = 3'b000;
                     width44 = 3'b000;
                     width43 = 3'b000;
                     width42 = 3'b000;
                     width41 = 3'b000;
                     width40 = 3'b000;
                     width39 = 3'b000;
                     width38 = 3'b000;
                     width37 = 3'b000;
                     width36 = 3'b000;
                     width35 = 3'b000;
                     width34 = 3'b000;
                     width33 = 3'b000;
                     width32 = 3'b000;
                     width31 = 3'b000;
                     width30 = 3'b000;
                     width29 = 3'b000;
                     width28 = 3'b000;
                     width27 = 3'b000;
                     width26 = 3'b000;
                     width25 = 3'b000;
                     width24 = 3'b000;
                     width23 = 3'b000;
                     width22 = 3'b000;
                     width21 = 3'b000;
                     width20 = 3'b000;
                     width19 = 3'b000;
                     width18 = 3'b000;
                     width17 = 3'b000;
                     width16 = 3'b000;
                     width15 = 3'b000;
                     width14 = 3'b000;
                     width13 = 3'b000;
                     width12 = 3'b000;
                     width11 = 3'b000;
                     width10 = 3'b000;
                     width9 = 3'b000;
                     width8 = 3'b000;
                     width7 = 3'b000;
                     width6 = 3'b000;
                     width5 = 3'b000;
                     width4 = 3'b011;
                     width3 = 3'b011;
                     width2 = 3'b011;
                     width1 = 3'b011;

                                    
                    writeAddr68 = {writeAddr[13:0]};
                    writeAddr67 = {writeAddr[13:0]};
                    writeAddr66 = {writeAddr[13:0]};
                    writeAddr65 = {writeAddr[13:0]};
                    writeAddr64 = {writeAddr[13:0]};
                    writeAddr63 = {writeAddr[13:0]};
                    writeAddr62 = {writeAddr[13:0]};
                    writeAddr61 = {writeAddr[13:0]};
                    writeAddr60 = {writeAddr[13:0]};
                    writeAddr59 = {writeAddr[13:0]};
                    writeAddr58 = {writeAddr[13:0]};
                    writeAddr57 = {writeAddr[13:0]};
                    writeAddr56 = {writeAddr[13:0]};
                    writeAddr55 = {writeAddr[13:0]};
                    writeAddr54 = {writeAddr[13:0]};
                    writeAddr53 = {writeAddr[13:0]};
                    writeAddr52 = {writeAddr[13:0]};
                    writeAddr51 = {writeAddr[13:0]};
                    writeAddr50 = {writeAddr[13:0]};
                    writeAddr49 = {writeAddr[13:0]};
                    writeAddr48 = {writeAddr[13:0]};
                    writeAddr47 = {writeAddr[13:0]};
                    writeAddr46 = {writeAddr[13:0]};
                    writeAddr45 = {writeAddr[13:0]};
                    writeAddr44 = {writeAddr[13:0]};
                    writeAddr43 = {writeAddr[13:0]};
                    writeAddr42 = {writeAddr[13:0]};
                    writeAddr41 = {writeAddr[13:0]};
                    writeAddr40 = {writeAddr[13:0]};
                    writeAddr39 = {writeAddr[13:0]};
                    writeAddr38 = {writeAddr[13:0]};
                    writeAddr37 = {writeAddr[13:0]};
                    writeAddr36 = {writeAddr[13:0]};
                    writeAddr35 = {writeAddr[13:0]};
                    writeAddr34 = {writeAddr[13:0]};
                    writeAddr33 = {writeAddr[13:0]};
                    writeAddr32 = {writeAddr[13:0]};
                    writeAddr31 = {writeAddr[13:0]};
                    writeAddr30 = {writeAddr[13:0]};
                    writeAddr29 = {writeAddr[13:0]};
                    writeAddr28 = {writeAddr[13:0]};
                    writeAddr27 = {writeAddr[13:0]};
                    writeAddr26 = {writeAddr[13:0]};
                    writeAddr25 = {writeAddr[13:0]};
                    writeAddr24 = {writeAddr[13:0]};
                    writeAddr23 = {writeAddr[13:0]};
                    writeAddr22 = {writeAddr[13:0]};
                    writeAddr21 = {writeAddr[13:0]};
                    writeAddr20 = {writeAddr[13:0]};
                    writeAddr19 = {writeAddr[13:0]};
                    writeAddr18 = {writeAddr[13:0]};
                    writeAddr17 = {writeAddr[13:0]};
                    writeAddr16 = {writeAddr[13:0]};
                    writeAddr15 = {writeAddr[13:0]};
                    writeAddr14 = {writeAddr[13:0]};
                    writeAddr13 = {writeAddr[13:0]};
                    writeAddr12 = {writeAddr[13:0]};
                    writeAddr11 = {writeAddr[13:0]};
                    writeAddr10 = {writeAddr[13:0]};
                    writeAddr9 = {writeAddr[13:0]};
                    writeAddr8 = {writeAddr[13:0]};
                    writeAddr7 = {writeAddr[13:0]};
                    writeAddr6 = {writeAddr[13:0]};
                    writeAddr5 = {writeAddr[13:0]};
                writeAddr4 = {writeAddr[10:0], 3'b0};
                writeAddr3 = {writeAddr[10:0], 3'b0};
             writeAddr2 = {writeAddr[10:0], 3'b0};
             writeAddr1 = {writeAddr[10:0], 3'b0};


                    readAddr68 = {readAddr[13:0]};
                    readAddr67 = {readAddr[13:0]};
                    readAddr66 = {readAddr[13:0]};
                    readAddr65 = {readAddr[13:0]};
                    readAddr64 = {readAddr[13:0]};
                    readAddr63 = {readAddr[13:0]};
                    readAddr62 = {readAddr[13:0]};
                    readAddr61 = {readAddr[13:0]};
                    readAddr60 = {readAddr[13:0]};
                    readAddr59 = {readAddr[13:0]};
                    readAddr58 = {readAddr[13:0]};
                    readAddr57 = {readAddr[13:0]};
                    readAddr56 = {readAddr[13:0]};
                    readAddr55 = {readAddr[13:0]};
                    readAddr54 = {readAddr[13:0]};
                    readAddr53 = {readAddr[13:0]};
                    readAddr52 = {readAddr[13:0]};
                    readAddr51 = {readAddr[13:0]};
                    readAddr50 = {readAddr[13:0]};
                    readAddr49 = {readAddr[13:0]};
                    readAddr48 = {readAddr[13:0]};
                    readAddr47 = {readAddr[13:0]};
                    readAddr46 = {readAddr[13:0]};
                    readAddr45 = {readAddr[13:0]};
                    readAddr44 = {readAddr[13:0]};
                    readAddr43 = {readAddr[13:0]};
                    readAddr42 = {readAddr[13:0]};
                    readAddr41 = {readAddr[13:0]};
                    readAddr40 = {readAddr[13:0]};
                    readAddr39 = {readAddr[13:0]};
                    readAddr38 = {readAddr[13:0]};
                    readAddr37 = {readAddr[13:0]};
                    readAddr36 = {readAddr[13:0]};
                    readAddr35 = {readAddr[13:0]};
                    readAddr34 = {readAddr[13:0]};
                    readAddr33 = {readAddr[13:0]};
                    readAddr32 = {readAddr[13:0]};
                    readAddr31 = {readAddr[13:0]};
                    readAddr30 = {readAddr[13:0]};
                    readAddr29 = {readAddr[13:0]};
                    readAddr28 = {readAddr[13:0]};
                    readAddr27 = {readAddr[13:0]};
                    readAddr26 = {readAddr[13:0]};
                    readAddr25 = {readAddr[13:0]};
                    readAddr24 = {readAddr[13:0]};
                    readAddr23 = {readAddr[13:0]};
                    readAddr22 = {readAddr[13:0]};
                    readAddr21 = {readAddr[13:0]};
                    readAddr20 = {readAddr[13:0]};
                    readAddr19 = {readAddr[13:0]};
                    readAddr18 = {readAddr[13:0]};
                    readAddr17 = {readAddr[13:0]};
                    readAddr16 = {readAddr[13:0]};
                    readAddr15 = {readAddr[13:0]};
                    readAddr14 = {readAddr[13:0]};
                    readAddr13 = {readAddr[13:0]};
                    readAddr12 = {readAddr[13:0]};
                    readAddr11 = {readAddr[13:0]};
                    readAddr10 = {readAddr[13:0]};
                    readAddr9 = {readAddr[13:0]};
                    readAddr8 = {readAddr[13:0]};
                    readAddr7 = {readAddr[13:0]};
                    readAddr6 = {readAddr[13:0]};
                    readAddr5 = {readAddr[13:0]};
                readAddr4  = {readAddr[10:0],  3'b0};
                readAddr3  = {readAddr[10:0],  3'b0};
                readAddr2  = {readAddr[10:0],  3'b0};
                readAddr1  = {readAddr[10:0],  3'b0};

                     writeData68 = {17'b0, writeData[31]};
                     writeData67 = {17'b0, writeData[30]};
                     writeData66 = {17'b0, writeData[29]};
                     writeData65 = {17'b0, writeData[28]};
                     writeData64 = {17'b0, writeData[27]};
                     writeData63 = {17'b0, writeData[26]};
                     writeData62 = {17'b0, writeData[25]};
                     writeData61 = {17'b0, writeData[24]};
                     writeData60 = {17'b0, writeData[23]};
                     writeData59 = {17'b0, writeData[22]};
                     writeData58 = {17'b0, writeData[21]};
                     writeData57 = {17'b0, writeData[20]};
                     writeData56 = {17'b0, writeData[19]};
                     writeData55 = {17'b0, writeData[18]};
                     writeData54 = {17'b0, writeData[17]};
                     writeData53 = {17'b0, writeData[16]};
                     writeData52 = {17'b0, writeData[15]};
                     writeData51 = {17'b0, writeData[14]};
                     writeData50 = {17'b0, writeData[13]};
                     writeData49 = {17'b0, writeData[12]};
                     writeData48 = {17'b0, writeData[11]};
                     writeData47 = {17'b0, writeData[10]};
                     writeData46 = {17'b0, writeData[9]};
                     writeData45 = {17'b0, writeData[8]};
                     writeData44 = {17'b0, writeData[7]};
                     writeData43 = {17'b0, writeData[6]};
                     writeData42 = {17'b0, writeData[5]};
                     writeData41 = {17'b0, writeData[4]};
                     writeData40 = {17'b0, writeData[3]};
                     writeData39 = {17'b0, writeData[2]};
                     writeData38 = {17'b0, writeData[1]};
                     writeData37 = {17'b0, writeData[0]};
                     writeData36 = {17'b0, writeData[31]};
                     writeData35 = {17'b0, writeData[30]};
                     writeData34 = {17'b0, writeData[29]};
                     writeData33 = {17'b0, writeData[28]};
                     writeData32 = {17'b0, writeData[27]};
                     writeData31 = {17'b0, writeData[26]};
                     writeData30 = {17'b0, writeData[25]};
                     writeData29 = {17'b0, writeData[24]};
                     writeData28 = {17'b0, writeData[23]};
                     writeData27 = {17'b0, writeData[22]};
                     writeData26 = {17'b0, writeData[21]};
                     writeData25 = {17'b0, writeData[20]};
                     writeData24 = {17'b0, writeData[19]};
                     writeData23 = {17'b0, writeData[18]};
                     writeData22 = {17'b0, writeData[17]};
                     writeData21 = {17'b0, writeData[16]};
                     writeData20 = {17'b0, writeData[15]};
                     writeData19 = {17'b0, writeData[14]};
                     writeData18 = {17'b0, writeData[13]};
                     writeData17 = {17'b0, writeData[12]};
                     writeData16 = {17'b0, writeData[11]};
                     writeData15 = {17'b0, writeData[10]};
                     writeData14 = {17'b0, writeData[9]};
                     writeData13 = {17'b0, writeData[8]};
                     writeData12 = {17'b0, writeData[7]};
                     writeData11 = {17'b0, writeData[6]};
                     writeData10 = {17'b0, writeData[5]};
                     writeData9 = {17'b0, writeData[4]};
                     writeData8 = {17'b0, writeData[3]};
                     writeData7 = {17'b0, writeData[2]};
                     writeData6 = {17'b0, writeData[1]};
                     writeData5 = {17'b0, writeData[0]};
                writeData4 = {10'b0, writeData[31:24]};
                writeData3 = {10'b0, writeData[23:16]};
                writeData2 = {10'b0, writeData[15:8]};
                writeData1 = {10'b0, writeData[7:0]};


                case (writeAddr[15:9])
                       7'b0000000, 7'b0000001, 7'b0000010, 7'b0000011,
                         7'b0000100, 7'b0000101, 7'b0000110, 7'b0000111,
                         7'b0001000, 7'b0001001, 7'b0001010, 7'b0001011,
                         7'b0001100, 7'b0001101, 7'b0001110, 7'b0001111,
                         7'b0010000, 7'b0010001, 7'b0010010, 7'b0010011,
                         7'b0010100, 7'b0010101, 7'b0010110, 7'b0010111,
                         7'b0011000, 7'b0011001, 7'b0011010, 7'b0011011,
                         7'b0011100, 7'b0011101, 7'b0011110, 7'b0011111 : begin
                            wen_a68 = {1'b0, wen};
                            wen_a67 = {1'b0, wen};
                            wen_a66 = {1'b0, wen};
                            wen_a65 = {1'b0, wen};
                            wen_a64 = {1'b0, wen};
                            wen_a63 = {1'b0, wen};
                            wen_a62 = {1'b0, wen};
                            wen_a61 = {1'b0, wen};
                            wen_a60 = {1'b0, wen};
                            wen_a59 = {1'b0, wen};
                            wen_a58 = {1'b0, wen};
                            wen_a57 = {1'b0, wen};
                            wen_a56 = {1'b0, wen};
                            wen_a55 = {1'b0, wen};
                            wen_a54 = {1'b0, wen};
                            wen_a53 = {1'b0, wen};
                            wen_a52 = {1'b0, wen};
                            wen_a51 = {1'b0, wen};
                            wen_a50 = {1'b0, wen};
                            wen_a49 = {1'b0, wen};
                            wen_a48 = {1'b0, wen};
                            wen_a47 = {1'b0, wen};
                            wen_a46 = {1'b0, wen};
                            wen_a45 = {1'b0, wen};
                            wen_a44 = {1'b0, wen};
                            wen_a43 = {1'b0, wen};
                            wen_a42 = {1'b0, wen};
                            wen_a41 = {1'b0, wen};
                            wen_a40 = {1'b0, wen};
                            wen_a39 = {1'b0, wen};
                            wen_a38 = {1'b0, wen};
                            wen_a37 = {1'b0, wen};
                            wen_a36 = {1'b0, 1'b0};
                            wen_a35 = {1'b0, 1'b0};
                            wen_a34 = {1'b0, 1'b0};
                            wen_a33 = {1'b0, 1'b0};
                            wen_a32 = {1'b0, 1'b0};
                            wen_a31 = {1'b0, 1'b0};
                            wen_a30 = {1'b0, 1'b0};
                            wen_a29 = {1'b0, 1'b0};
                            wen_a28 = {1'b0, 1'b0};
                            wen_a27 = {1'b0, 1'b0};
                            wen_a26 = {1'b0, 1'b0};
                            wen_a25 = {1'b0, 1'b0};
                            wen_a24 = {1'b0, 1'b0};
                            wen_a23 = {1'b0, 1'b0};
                            wen_a22 = {1'b0, 1'b0};
                            wen_a21 = {1'b0, 1'b0};
                            wen_a20 = {1'b0, 1'b0};
                            wen_a19 = {1'b0, 1'b0};
                            wen_a18 = {1'b0, 1'b0};
                            wen_a17 = {1'b0, 1'b0};
                            wen_a16 = {1'b0, 1'b0};
                            wen_a15 = {1'b0, 1'b0};
                            wen_a14 = {1'b0, 1'b0};
                            wen_a13 = {1'b0, 1'b0};
                            wen_a12 = {1'b0, 1'b0};
                            wen_a11 = {1'b0, 1'b0};
                            wen_a10 = {1'b0, 1'b0};
                            wen_a9  = {1'b0, 1'b0};
                            wen_a8  = {1'b0, 1'b0};
                            wen_a7  = {1'b0, 1'b0};
                            wen_a6  = {1'b0, 1'b0};
                            wen_a5  = {1'b0, 1'b0};
                            wen_a4  = {1'b0, 1'b0};
                            wen_a3  = {1'b0, 1'b0};
                            wen_a2  = {1'b0, 1'b0};
                            wen_a1  = {1'b0, 1'b0};
                    end        
                         7'b0100000, 7'b0100001, 7'b0100010, 7'b0100011,
                         7'b0100100, 7'b0100101, 7'b0100110, 7'b0100111,
                         7'b0101000, 7'b0101001, 7'b0101010, 7'b0101011,
                         7'b0101100, 7'b0101101, 7'b0101110, 7'b0101111,
                         7'b0110000, 7'b0110001, 7'b0110010, 7'b0110011,
                         7'b0110100, 7'b0110101, 7'b0110110, 7'b0110111,             
                         7'b0111000, 7'b0111001, 7'b0111010, 7'b0111011,
                         7'b0111100, 7'b0111101, 7'b0111110, 7'b0111111  : begin
                            wen_a68 = {1'b0, 1'b0};
                            wen_a67 = {1'b0, 1'b0};
                            wen_a66 = {1'b0, 1'b0};
                            wen_a65 = {1'b0, 1'b0};
                            wen_a64 = {1'b0, 1'b0};
                            wen_a63 = {1'b0, 1'b0};
                            wen_a62 = {1'b0, 1'b0};
                            wen_a61 = {1'b0, 1'b0};
                            wen_a60 = {1'b0, 1'b0};
                            wen_a59 = {1'b0, 1'b0};
                            wen_a58 = {1'b0, 1'b0};
                            wen_a57 = {1'b0, 1'b0};
                            wen_a56 = {1'b0, 1'b0};
                            wen_a55 = {1'b0, 1'b0};
                            wen_a54 = {1'b0, 1'b0};
                            wen_a53 = {1'b0, 1'b0};
                            wen_a52 = {1'b0, 1'b0};
                            wen_a51 = {1'b0, 1'b0};
                            wen_a50 = {1'b0, 1'b0};
                            wen_a49 = {1'b0, 1'b0};
                            wen_a48 = {1'b0, 1'b0};
                            wen_a47 = {1'b0, 1'b0};
                            wen_a46 = {1'b0, 1'b0};
                            wen_a45 = {1'b0, 1'b0};
                            wen_a44 = {1'b0, 1'b0};
                            wen_a43 = {1'b0, 1'b0};
                            wen_a42 = {1'b0, 1'b0};
                            wen_a41 = {1'b0, 1'b0};
                            wen_a40 = {1'b0, 1'b0};
                            wen_a39 = {1'b0, 1'b0};
                            wen_a38 = {1'b0, 1'b0};
                            wen_a37 = {1'b0, 1'b0};
                            wen_a36 = {1'b0, wen};
                            wen_a35 = {1'b0, wen};
                            wen_a34 = {1'b0, wen};
                            wen_a33 = {1'b0, wen};
                            wen_a32 = {1'b0, wen};
                            wen_a31 = {1'b0, wen};
                            wen_a30 = {1'b0, wen};
                            wen_a29 = {1'b0, wen};
                            wen_a28 = {1'b0, wen};
                            wen_a27 = {1'b0, wen};
                            wen_a26 = {1'b0, wen};
                            wen_a25 = {1'b0, wen};
                            wen_a24 = {1'b0, wen};
                            wen_a23 = {1'b0, wen};
                            wen_a22 = {1'b0, wen};
                            wen_a21 = {1'b0, wen};
                            wen_a20 = {1'b0, wen};
                            wen_a19 = {1'b0, wen};
                            wen_a18 = {1'b0, wen};
                            wen_a17 = {1'b0, wen};
                            wen_a16 = {1'b0, wen};
                            wen_a15 = {1'b0, wen};
                            wen_a14 = {1'b0, wen};
                            wen_a13 = {1'b0, wen};
                            wen_a12 = {1'b0, wen};
                            wen_a11 = {1'b0, wen};
                            wen_a10 = {1'b0, wen};
                            wen_a9  = {1'b0, wen};
                            wen_a8  = {1'b0, wen};
                            wen_a7  = {1'b0, wen};
                            wen_a6  = {1'b0, wen};
                            wen_a5  = {1'b0, wen};
                            wen_a4  = {1'b0, 1'b0};
                            wen_a3  = {1'b0, 1'b0};
                            wen_a2  = {1'b0, 1'b0};
                            wen_a1  = {1'b0, 1'b0};

                    end        

                     7'b1000000, 7'b1000001, 7'b1000010, 7'b1000011 : begin
                        wen_a68 = {1'b0, 1'b0};
                        wen_a67 = {1'b0, 1'b0};
                        wen_a66 = {1'b0, 1'b0};
                        wen_a65 = {1'b0, 1'b0};
                        wen_a64 = {1'b0, 1'b0};
                        wen_a63 = {1'b0, 1'b0};
                        wen_a62 = {1'b0, 1'b0};
                        wen_a61 = {1'b0, 1'b0};
                        wen_a60 = {1'b0, 1'b0};
                        wen_a59 = {1'b0, 1'b0};
                        wen_a58 = {1'b0, 1'b0};
                        wen_a57 = {1'b0, 1'b0};
                        wen_a56 = {1'b0, 1'b0};
                        wen_a55 = {1'b0, 1'b0};
                        wen_a54 = {1'b0, 1'b0};
                        wen_a53 = {1'b0, 1'b0};
                        wen_a52 = {1'b0, 1'b0};
                        wen_a51 = {1'b0, 1'b0};
                        wen_a50 = {1'b0, 1'b0};
                        wen_a49 = {1'b0, 1'b0};
                        wen_a48 = {1'b0, 1'b0};
                        wen_a47 = {1'b0, 1'b0};
                        wen_a46 = {1'b0, 1'b0};
                        wen_a45 = {1'b0, 1'b0};
                        wen_a44 = {1'b0, 1'b0};
                        wen_a43 = {1'b0, 1'b0};
                        wen_a42 = {1'b0, 1'b0};
                        wen_a41 = {1'b0, 1'b0};
                        wen_a40 = {1'b0, 1'b0};
                        wen_a39 = {1'b0, 1'b0};
                        wen_a38 = {1'b0, 1'b0};
                        wen_a37 = {1'b0, 1'b0};
                        wen_a36 = {1'b0, 1'b0};
                        wen_a35 = {1'b0, 1'b0};
                        wen_a34 = {1'b0, 1'b0};
                        wen_a33 = {1'b0, 1'b0};
                        wen_a32 = {1'b0, 1'b0};
                        wen_a31 = {1'b0, 1'b0};
                        wen_a30 = {1'b0, 1'b0};
                        wen_a29 = {1'b0, 1'b0};
                        wen_a28 = {1'b0, 1'b0};
                        wen_a27 = {1'b0, 1'b0};
                        wen_a26 = {1'b0, 1'b0};
                        wen_a25 = {1'b0, 1'b0};
                        wen_a24 = {1'b0, 1'b0};
                        wen_a23 = {1'b0, 1'b0};
                        wen_a22 = {1'b0, 1'b0};
                        wen_a21 = {1'b0, 1'b0};
                        wen_a20 = {1'b0, 1'b0};
                        wen_a19 = {1'b0, 1'b0};
                        wen_a18 = {1'b0, 1'b0};
                        wen_a17 = {1'b0, 1'b0};
                        wen_a16 = {1'b0, 1'b0};
                        wen_a15 = {1'b0, 1'b0};
                        wen_a14 = {1'b0, 1'b0};
                        wen_a13 = {1'b0, 1'b0};
                        wen_a12 = {1'b0, 1'b0};
                        wen_a11 = {1'b0, 1'b0};
                        wen_a10 = {1'b0, 1'b0};
                        wen_a9 = {1'b0, 1'b0};
                        wen_a8 = {1'b0, 1'b0};
                        wen_a7 = {1'b0, 1'b0};
                        wen_a6 = {1'b0, 1'b0};
                        wen_a5 = {1'b0, 1'b0};
                        wen_a4 = {1'b0, wen};
                        wen_a3 = {1'b0, wen};
                        wen_a2 = {1'b0, wen};
                        wen_a1 = {1'b0, wen};
                    end
                    default : begin
                        wen_a68 = {1'b0, 1'b0};
                        wen_a67 = {1'b0, 1'b0};
                        wen_a66 = {1'b0, 1'b0};
                        wen_a65 = {1'b0, 1'b0};
                        wen_a64 = {1'b0, 1'b0};
                        wen_a63 = {1'b0, 1'b0};
                        wen_a62 = {1'b0, 1'b0};
                        wen_a61 = {1'b0, 1'b0};
                        wen_a60 = {1'b0, 1'b0};
                        wen_a59 = {1'b0, 1'b0};
                        wen_a58 = {1'b0, 1'b0};
                        wen_a57 = {1'b0, 1'b0};
                        wen_a56 = {1'b0, 1'b0};
                        wen_a55 = {1'b0, 1'b0};
                        wen_a54 = {1'b0, 1'b0};
                        wen_a53 = {1'b0, 1'b0};
                        wen_a52 = {1'b0, 1'b0};
                        wen_a51 = {1'b0, 1'b0};
                        wen_a50 = {1'b0, 1'b0};
                        wen_a49 = {1'b0, 1'b0};
                        wen_a48 = {1'b0, 1'b0};
                        wen_a47 = {1'b0, 1'b0};
                        wen_a46 = {1'b0, 1'b0};
                        wen_a45 = {1'b0, 1'b0};
                        wen_a44 = {1'b0, 1'b0};
                        wen_a43 = {1'b0, 1'b0};
                        wen_a42 = {1'b0, 1'b0};
                        wen_a41 = {1'b0, 1'b0};
                        wen_a40 = {1'b0, 1'b0};
                        wen_a39 = {1'b0, 1'b0};
                        wen_a38 = {1'b0, 1'b0};
                        wen_a37 = {1'b0, 1'b0};
                        wen_a36 = {1'b0, 1'b0};
                        wen_a35 = {1'b0, 1'b0};
                        wen_a34 = {1'b0, 1'b0};
                        wen_a33 = {1'b0, 1'b0};
                        wen_a32 = {1'b0, 1'b0};
                        wen_a31 = {1'b0, 1'b0};
                        wen_a30 = {1'b0, 1'b0};
                        wen_a29 = {1'b0, 1'b0};
                        wen_a28 = {1'b0, 1'b0};
                        wen_a27 = {1'b0, 1'b0};
                        wen_a26 = {1'b0, 1'b0};
                        wen_a25 = {1'b0, 1'b0};
                        wen_a24 = {1'b0, 1'b0};
                        wen_a23 = {1'b0, 1'b0};
                        wen_a22 = {1'b0, 1'b0};
                        wen_a21 = {1'b0, 1'b0};
                        wen_a20 = {1'b0, 1'b0};
                        wen_a19 = {1'b0, 1'b0};
                        wen_a18 = {1'b0, 1'b0};
                        wen_a17 = {1'b0, 1'b0};
                        wen_a16 = {1'b0, 1'b0};
                        wen_a15 = {1'b0, 1'b0};
                        wen_a14 = {1'b0, 1'b0};
                        wen_a13 = {1'b0, 1'b0};
                        wen_a12 = {1'b0, 1'b0};
                        wen_a11 = {1'b0, 1'b0};
                        wen_a10 = {1'b0, 1'b0};
                        wen_a9 = {1'b0, 1'b0};
                        wen_a8 = {1'b0, 1'b0};
                        wen_a7 = {1'b0, 1'b0};
                        wen_a6 = {1'b0, 1'b0};
                        wen_a5 = {1'b0, 1'b0};
                        wen_a4 = {1'b0, 1'b0};
                        wen_a3 = {1'b0, 1'b0};
                        wen_a2 = {1'b0, 1'b0};
                        wen_a1 = {1'b0, 1'b0};
                    end
               endcase // case (writeAddr[15:9])

                case (ckRdAddr[15:9])

                       7'b0000000, 7'b0000001, 7'b0000010, 7'b0000011,
                         7'b0000100, 7'b0000101, 7'b0000110, 7'b0000111,
                         7'b0001000, 7'b0001001, 7'b0001010, 7'b0001011,
                         7'b0001100, 7'b0001101, 7'b0001110, 7'b0001111,
                         7'b0010000, 7'b0010001, 7'b0010010, 7'b0010011,
                         7'b0010100, 7'b0010101, 7'b0010110, 7'b0010111,
                         7'b0011000, 7'b0011001, 7'b0011010, 7'b0011011,
                         7'b0011100, 7'b0011101, 7'b0011110, 7'b0011111  : begin
                        readData = {
                                        readData68[0],
                                        readData67[0],
                                        readData66[0],
                                        readData65[0],
                                        readData64[0],
                                        readData63[0],
                                        readData62[0],
                                        readData61[0],
                                        readData60[0],
                                        readData59[0],
                                        readData58[0],
                                        readData57[0],
                                        readData56[0],
                                        readData55[0], 
                                        readData54[0],
                                        readData53[0],
                                        readData52[0],
                                        readData51[0],
                                        readData50[0],
                                        readData49[0],
                                        readData48[0],
                                        readData47[0],
                                        readData46[0],
                                        readData45[0],
                                        readData44[0],
                                        readData43[0],
                                        readData42[0],
                                        readData41[0],
                                        readData40[0],
                                        readData39[0],
                                        readData38[0],
                                        readData37[0]
                        };
                    end
                  7'b0100000, 7'b0100001, 7'b0100010, 7'b0100011,
                    7'b0100100, 7'b0100101, 7'b0100110, 7'b0100111,
                    7'b0101000, 7'b0101001, 7'b0101010, 7'b0101011,
                    7'b0101100, 7'b0101101, 7'b0101110, 7'b0101111,
                    7'b0110000, 7'b0110001, 7'b0110010, 7'b0110011,
                    7'b0110100, 7'b0110101, 7'b0110110, 7'b0110111,             
                    7'b0111000, 7'b0111001, 7'b0111010, 7'b0111011,
                    7'b0111100, 7'b0111101, 7'b0111110, 7'b0111111 : begin
                       readData = {
                                        readData36[0],
                                        readData35[0],
                                        readData34[0],
                                        readData33[0],
                                        readData32[0],
                                        readData31[0],
                                        readData30[0],
                                        readData29[0],
                                        readData28[0],
                                        readData27[0],
                                        readData26[0],
                                        readData25[0],
                                        readData24[0],
                                        readData23[0],
                                        readData22[0],
                                        readData21[0],
                                        readData20[0],
                                        readData19[0],
                                        readData18[0],
                                        readData17[0],
                                        readData16[0],
                                        readData15[0],
                                        readData14[0],
                                        readData13[0],
                                        readData12[0],
                                        readData11[0],
                                        readData10[0],
                                        readData9[0],
                                        readData8[0],
                                        readData7[0],
                                        readData6[0],
                                        readData5[0]
                                   };

                    end
                    7'b1000000, 7'b1000001, 7'b1000010, 7'b1000011 : begin
                        readData = {readData4[7:0],readData3[7:0],readData2[7:0],readData1[7:0]};
                    end
                    default : begin
                       readData = 32'b0;
                    end
               endcase // case (ckRdAddr[15:9])                                    
           end // case: 34816
          35328: begin
                     width68 = 3'b000;
                     width67 = 3'b000;
                     width66 = 3'b000;
                     width65 = 3'b000;
                     width64 = 3'b000;
                     width63 = 3'b000;
                     width62 = 3'b000;
                     width61 = 3'b000;
                     width60 = 3'b000;
                     width59 = 3'b000;
                     width58 = 3'b000;
                     width57 = 3'b000;
                     width56 = 3'b000;
                     width55 = 3'b000;
                     width54 = 3'b000;
                     width53 = 3'b000;
                     width52 = 3'b000;
                     width51 = 3'b000;
                     width50 = 3'b000;
                     width49 = 3'b000;
                     width48 = 3'b000;
                     width47 = 3'b000;
                     width46 = 3'b000;
                     width45 = 3'b000;
                     width44 = 3'b000;
                     width43 = 3'b000;
                     width42 = 3'b000;
                     width41 = 3'b000;
                     width40 = 3'b000;
                     width39 = 3'b000;
                     width38 = 3'b000;
                     width37 = 3'b000;
                     width36 = 3'b000;
                     width35 = 3'b000;
                     width34 = 3'b000;
                     width33 = 3'b000;
                     width32 = 3'b000;
                     width31 = 3'b000;
                     width30 = 3'b000;
                     width29 = 3'b000;
                     width28 = 3'b000;
                     width27 = 3'b000;
                     width26 = 3'b000;
                     width25 = 3'b000;
                     width24 = 3'b000;
                     width23 = 3'b000;
                     width22 = 3'b000;
                     width21 = 3'b000;
                     width20 = 3'b000;
                     width19 = 3'b000;
                     width18 = 3'b000;
                     width17 = 3'b000;
                     width16 = 3'b000;
                     width15 = 3'b000;
                     width14 = 3'b000;
                     width13 = 3'b000;
                     width12 = 3'b000;
                     width11 = 3'b000;
                     width10 = 3'b000;
                     width9 = 3'b000;
                     width8 = 3'b000;
                     width7 = 3'b000;
                     width6 = 3'b000;
                     width5 = 3'b000;
                     width4 = 3'b011;
                     width3 = 3'b011;
                     width2 = 3'b011;
                     width1 = 3'b011;
                     width0 = 3'b101;
                                    
                    writeAddr68 = {writeAddr[13:0]};
                    writeAddr67 = {writeAddr[13:0]};
                    writeAddr66 = {writeAddr[13:0]};
                    writeAddr65 = {writeAddr[13:0]};
                    writeAddr64 = {writeAddr[13:0]};
                    writeAddr63 = {writeAddr[13:0]};
                    writeAddr62 = {writeAddr[13:0]};
                    writeAddr61 = {writeAddr[13:0]};
                    writeAddr60 = {writeAddr[13:0]};
                    writeAddr59 = {writeAddr[13:0]};
                    writeAddr58 = {writeAddr[13:0]};
                    writeAddr57 = {writeAddr[13:0]};
                    writeAddr56 = {writeAddr[13:0]};
                    writeAddr55 = {writeAddr[13:0]};
                    writeAddr54 = {writeAddr[13:0]};
                    writeAddr53 = {writeAddr[13:0]};
                    writeAddr52 = {writeAddr[13:0]};
                    writeAddr51 = {writeAddr[13:0]};
                    writeAddr50 = {writeAddr[13:0]};
                    writeAddr49 = {writeAddr[13:0]};
                    writeAddr48 = {writeAddr[13:0]};
                    writeAddr47 = {writeAddr[13:0]};
                    writeAddr46 = {writeAddr[13:0]};
                    writeAddr45 = {writeAddr[13:0]};
                    writeAddr44 = {writeAddr[13:0]};
                    writeAddr43 = {writeAddr[13:0]};
                    writeAddr42 = {writeAddr[13:0]};
                    writeAddr41 = {writeAddr[13:0]};
                    writeAddr40 = {writeAddr[13:0]};
                    writeAddr39 = {writeAddr[13:0]};
                    writeAddr38 = {writeAddr[13:0]};
                    writeAddr37 = {writeAddr[13:0]};
                    writeAddr36 = {writeAddr[13:0]};
                    writeAddr35 = {writeAddr[13:0]};
                    writeAddr34 = {writeAddr[13:0]};
                    writeAddr33 = {writeAddr[13:0]};
                    writeAddr32 = {writeAddr[13:0]};
                    writeAddr31 = {writeAddr[13:0]};
                    writeAddr30 = {writeAddr[13:0]};
                    writeAddr29 = {writeAddr[13:0]};
                    writeAddr28 = {writeAddr[13:0]};
                    writeAddr27 = {writeAddr[13:0]};
                    writeAddr26 = {writeAddr[13:0]};
                    writeAddr25 = {writeAddr[13:0]};
                    writeAddr24 = {writeAddr[13:0]};
                    writeAddr23 = {writeAddr[13:0]};
                    writeAddr22 = {writeAddr[13:0]};
                    writeAddr21 = {writeAddr[13:0]};
                    writeAddr20 = {writeAddr[13:0]};
                    writeAddr19 = {writeAddr[13:0]};
                    writeAddr18 = {writeAddr[13:0]};
                    writeAddr17 = {writeAddr[13:0]};
                    writeAddr16 = {writeAddr[13:0]};
                    writeAddr15 = {writeAddr[13:0]};
                    writeAddr14 = {writeAddr[13:0]};
                    writeAddr13 = {writeAddr[13:0]};
                    writeAddr12 = {writeAddr[13:0]};
                    writeAddr11 = {writeAddr[13:0]};
                    writeAddr10 = {writeAddr[13:0]};
                    writeAddr9 = {writeAddr[13:0]};
                    writeAddr8 = {writeAddr[13:0]};
                    writeAddr7 = {writeAddr[13:0]};
                    writeAddr6 = {writeAddr[13:0]};
                    writeAddr5 = {writeAddr[13:0]};
                    writeAddr4 = {writeAddr[10:0], 3'b0};
                    writeAddr3 = {writeAddr[10:0], 3'b0};
                    writeAddr2 = {writeAddr[10:0], 3'b0};
                    writeAddr1 = {writeAddr[10:0], 3'b0};
                    writeAddr0 = {writeAddr[8:0], 5'b0};

                    readAddr68 = {readAddr[13:0]};
                    readAddr67 = {readAddr[13:0]};
                    readAddr66 = {readAddr[13:0]};
                    readAddr65 = {readAddr[13:0]};
                    readAddr64 = {readAddr[13:0]};
                    readAddr63 = {readAddr[13:0]};
                    readAddr62 = {readAddr[13:0]};
                    readAddr61 = {readAddr[13:0]};
                    readAddr60 = {readAddr[13:0]};
                    readAddr59 = {readAddr[13:0]};
                    readAddr58 = {readAddr[13:0]};
                    readAddr57 = {readAddr[13:0]};
                    readAddr56 = {readAddr[13:0]};
                    readAddr55 = {readAddr[13:0]};
                    readAddr54 = {readAddr[13:0]};
                    readAddr53 = {readAddr[13:0]};
                    readAddr52 = {readAddr[13:0]};
                    readAddr51 = {readAddr[13:0]};
                    readAddr50 = {readAddr[13:0]};
                    readAddr49 = {readAddr[13:0]};
                    readAddr48 = {readAddr[13:0]};
                    readAddr47 = {readAddr[13:0]};
                    readAddr46 = {readAddr[13:0]};
                    readAddr45 = {readAddr[13:0]};
                    readAddr44 = {readAddr[13:0]};
                    readAddr43 = {readAddr[13:0]};
                    readAddr42 = {readAddr[13:0]};
                    readAddr41 = {readAddr[13:0]};
                    readAddr40 = {readAddr[13:0]};
                    readAddr39 = {readAddr[13:0]};
                    readAddr38 = {readAddr[13:0]};
                    readAddr37 = {readAddr[13:0]};
                    readAddr36 = {readAddr[13:0]};
                    readAddr35 = {readAddr[13:0]};
                    readAddr34 = {readAddr[13:0]};
                    readAddr33 = {readAddr[13:0]};
                    readAddr32 = {readAddr[13:0]};
                    readAddr31 = {readAddr[13:0]};
                    readAddr30 = {readAddr[13:0]};
                    readAddr29 = {readAddr[13:0]};
                    readAddr28 = {readAddr[13:0]};
                    readAddr27 = {readAddr[13:0]};
                    readAddr26 = {readAddr[13:0]};
                    readAddr25 = {readAddr[13:0]};
                    readAddr24 = {readAddr[13:0]};
                    readAddr23 = {readAddr[13:0]};
                    readAddr22 = {readAddr[13:0]};
                    readAddr21 = {readAddr[13:0]};
                    readAddr20 = {readAddr[13:0]};
                    readAddr19 = {readAddr[13:0]};
                    readAddr18 = {readAddr[13:0]};
                    readAddr17 = {readAddr[13:0]};
                    readAddr16 = {readAddr[13:0]};
                    readAddr15 = {readAddr[13:0]};
                    readAddr14 = {readAddr[13:0]};
                    readAddr13 = {readAddr[13:0]};
                    readAddr12 = {readAddr[13:0]};
                    readAddr11 = {readAddr[13:0]};
                    readAddr10 = {readAddr[13:0]};
                    readAddr9 = {readAddr[13:0]};
                    readAddr8 = {readAddr[13:0]};
                    readAddr7 = {readAddr[13:0]};
                    readAddr6 = {readAddr[13:0]};
                    readAddr5 = {readAddr[13:0]};
                    readAddr4  = {readAddr[10:0],  3'b0};
                    readAddr3  = {readAddr[10:0],  3'b0};
                    readAddr2  = {readAddr[10:0],  3'b0};
                    readAddr1  = {readAddr[10:0],  3'b0};
                    readAddr0  = {readAddr[8:0],  5'b0};

                     writeData68 = {17'b0, writeData[31]};
                     writeData67 = {17'b0, writeData[30]};
                     writeData66 = {17'b0, writeData[29]};
                     writeData65 = {17'b0, writeData[28]};
                     writeData64 = {17'b0, writeData[27]};
                     writeData63 = {17'b0, writeData[26]};
                     writeData62 = {17'b0, writeData[25]};
                     writeData61 = {17'b0, writeData[24]};
                     writeData60 = {17'b0, writeData[23]};
                     writeData59 = {17'b0, writeData[22]};
                     writeData58 = {17'b0, writeData[21]};
                     writeData57 = {17'b0, writeData[20]};
                     writeData56 = {17'b0, writeData[19]};
                     writeData55 = {17'b0, writeData[18]};
                     writeData54 = {17'b0, writeData[17]};
                     writeData53 = {17'b0, writeData[16]};
                     writeData52 = {17'b0, writeData[15]};
                     writeData51 = {17'b0, writeData[14]};
                     writeData50 = {17'b0, writeData[13]};
                     writeData49 = {17'b0, writeData[12]};
                     writeData48 = {17'b0, writeData[11]};
                     writeData47 = {17'b0, writeData[10]};
                     writeData46 = {17'b0, writeData[9]};
                     writeData45 = {17'b0, writeData[8]};
                     writeData44 = {17'b0, writeData[7]};
                     writeData43 = {17'b0, writeData[6]};
                     writeData42 = {17'b0, writeData[5]};
                     writeData41 = {17'b0, writeData[4]};
                     writeData40 = {17'b0, writeData[3]};
                     writeData39 = {17'b0, writeData[2]};
                     writeData38 = {17'b0, writeData[1]};
                     writeData37 = {17'b0, writeData[0]};
                     writeData36 = {17'b0, writeData[31]};
                     writeData35 = {17'b0, writeData[30]};
                     writeData34 = {17'b0, writeData[29]};
                     writeData33 = {17'b0, writeData[28]};
                     writeData32 = {17'b0, writeData[27]};
                     writeData31 = {17'b0, writeData[26]};
                     writeData30 = {17'b0, writeData[25]};
                     writeData29 = {17'b0, writeData[24]};
                     writeData28 = {17'b0, writeData[23]};
                     writeData27 = {17'b0, writeData[22]};
                     writeData26 = {17'b0, writeData[21]};
                     writeData25 = {17'b0, writeData[20]};
                     writeData24 = {17'b0, writeData[19]};
                     writeData23 = {17'b0, writeData[18]};
                     writeData22 = {17'b0, writeData[17]};
                     writeData21 = {17'b0, writeData[16]};
                     writeData20 = {17'b0, writeData[15]};
                     writeData19 = {17'b0, writeData[14]};
                     writeData18 = {17'b0, writeData[13]};
                     writeData17 = {17'b0, writeData[12]};
                     writeData16 = {17'b0, writeData[11]};
                     writeData15 = {17'b0, writeData[10]};
                     writeData14 = {17'b0, writeData[9]};
                     writeData13 = {17'b0, writeData[8]};
                     writeData12 = {17'b0, writeData[7]};
                     writeData11 = {17'b0, writeData[6]};
                     writeData10 = {17'b0, writeData[5]};
                     writeData9 = {17'b0, writeData[4]};
                     writeData8 = {17'b0, writeData[3]};
                     writeData7 = {17'b0, writeData[2]};
                     writeData6 = {17'b0, writeData[1]};
                     writeData5 = {17'b0, writeData[0]};
                writeData4 = {10'b0, writeData[31:24]};
                writeData3 = {10'b0, writeData[23:16]};
                writeData2 = {10'b0, writeData[15:8]};
                writeData1 = {10'b0, writeData[7:0]};
                writeData0 = {1'b0, writeData[31:24], 1'b0, writeData[23:16], 1'b0, writeData[15:8], 1'b0, writeData[7:0]};

                case (writeAddr[15:9])
                  7'b0000000, 7'b0000001, 7'b0000010, 7'b0000011,
                         7'b0000100, 7'b0000101, 7'b0000110, 7'b0000111,
                         7'b0001000, 7'b0001001, 7'b0001010, 7'b0001011,
                         7'b0001100, 7'b0001101, 7'b0001110, 7'b0001111,
                         7'b0010000, 7'b0010001, 7'b0010010, 7'b0010011,
                         7'b0010100, 7'b0010101, 7'b0010110, 7'b0010111,
                         7'b0011000, 7'b0011001, 7'b0011010, 7'b0011011,
                         7'b0011100, 7'b0011101, 7'b0011110, 7'b0011111 : begin
                            wen_a68 = {1'b0, wen};
                            wen_a67 = {1'b0, wen};
                            wen_a66 = {1'b0, wen};
                            wen_a65 = {1'b0, wen};
                            wen_a64 = {1'b0, wen};
                            wen_a63 = {1'b0, wen};
                            wen_a62 = {1'b0, wen};
                            wen_a61 = {1'b0, wen};
                            wen_a60 = {1'b0, wen};
                            wen_a59 = {1'b0, wen};
                            wen_a58 = {1'b0, wen};
                            wen_a57 = {1'b0, wen};
                            wen_a56 = {1'b0, wen};
                            wen_a55 = {1'b0, wen};
                            wen_a54 = {1'b0, wen};
                            wen_a53 = {1'b0, wen};
                            wen_a52 = {1'b0, wen};
                            wen_a51 = {1'b0, wen};
                            wen_a50 = {1'b0, wen};
                            wen_a49 = {1'b0, wen};
                            wen_a48 = {1'b0, wen};
                            wen_a47 = {1'b0, wen};
                            wen_a46 = {1'b0, wen};
                            wen_a45 = {1'b0, wen};
                            wen_a44 = {1'b0, wen};
                            wen_a43 = {1'b0, wen};
                            wen_a42 = {1'b0, wen};
                            wen_a41 = {1'b0, wen};
                            wen_a40 = {1'b0, wen};
                            wen_a39 = {1'b0, wen};
                            wen_a38 = {1'b0, wen};
                            wen_a37 = {1'b0, wen};
                        wen_a36 = {1'b0, 1'b0};
                        wen_a35 = {1'b0, 1'b0};
                        wen_a34 = {1'b0, 1'b0};
                        wen_a33 = {1'b0, 1'b0};
                        wen_a32 = {1'b0, 1'b0};
                        wen_a31 = {1'b0, 1'b0};
                        wen_a30 = {1'b0, 1'b0};
                        wen_a29 = {1'b0, 1'b0};
                        wen_a28 = {1'b0, 1'b0};
                        wen_a27 = {1'b0, 1'b0};
                        wen_a26 = {1'b0, 1'b0};
                        wen_a25 = {1'b0, 1'b0};
                        wen_a24 = {1'b0, 1'b0};
                        wen_a23 = {1'b0, 1'b0};
                        wen_a22 = {1'b0, 1'b0};
                        wen_a21 = {1'b0, 1'b0};
                        wen_a20 = {1'b0, 1'b0};
                        wen_a19 = {1'b0, 1'b0};
                        wen_a18 = {1'b0, 1'b0};
                        wen_a17 = {1'b0, 1'b0};
                        wen_a16 = {1'b0, 1'b0};
                        wen_a15 = {1'b0, 1'b0};
                        wen_a14 = {1'b0, 1'b0};
                        wen_a13 = {1'b0, 1'b0};
                        wen_a12 = {1'b0, 1'b0};
                        wen_a11 = {1'b0, 1'b0};
                        wen_a10 = {1'b0, 1'b0};
                        wen_a9 = {1'b0, 1'b0};
                        wen_a8 = {1'b0, 1'b0};
                        wen_a7 = {1'b0, 1'b0};
                        wen_a6 = {1'b0, 1'b0};
                        wen_a5 = {1'b0, 1'b0};
                        wen_a4 = {1'b0, 1'b0};
                        wen_a3 = {1'b0, 1'b0};
                        wen_a2 = {1'b0, 1'b0};
                        wen_a1 = {1'b0, 1'b0};
                        wen_a0 = {1'b0, 1'b0};
                        wen_b0 = {1'b0, 1'b0};
                    end
                         7'b0100000, 7'b0100001, 7'b0100010, 7'b0100011,
                         7'b0100100, 7'b0100101, 7'b0100110, 7'b0100111,
                         7'b0101000, 7'b0101001, 7'b0101010, 7'b0101011,
                         7'b0101100, 7'b0101101, 7'b0101110, 7'b0101111,
                         7'b0110000, 7'b0110001, 7'b0110010, 7'b0110011,
                         7'b0110100, 7'b0110101, 7'b0110110, 7'b0110111,             
                         7'b0111000, 7'b0111001, 7'b0111010, 7'b0111011,
                         7'b0111100, 7'b0111101, 7'b0111110, 7'b0111111  : begin
                            wen_a68 = {1'b0, 1'b0};
                            wen_a67 = {1'b0, 1'b0};
                            wen_a66 = {1'b0, 1'b0};
                            wen_a65 = {1'b0, 1'b0};
                            wen_a64 = {1'b0, 1'b0};
                            wen_a63 = {1'b0, 1'b0};
                            wen_a62 = {1'b0, 1'b0};
                            wen_a61 = {1'b0, 1'b0};
                            wen_a60 = {1'b0, 1'b0};
                            wen_a59 = {1'b0, 1'b0};
                            wen_a58 = {1'b0, 1'b0};
                            wen_a57 = {1'b0, 1'b0};
                            wen_a56 = {1'b0, 1'b0};
                            wen_a55 = {1'b0, 1'b0};
                            wen_a54 = {1'b0, 1'b0};
                            wen_a53 = {1'b0, 1'b0};
                            wen_a52 = {1'b0, 1'b0};
                            wen_a51 = {1'b0, 1'b0};
                            wen_a50 = {1'b0, 1'b0};
                            wen_a49 = {1'b0, 1'b0};
                            wen_a48 = {1'b0, 1'b0};
                            wen_a47 = {1'b0, 1'b0};
                            wen_a46 = {1'b0, 1'b0};
                            wen_a45 = {1'b0, 1'b0};
                            wen_a44 = {1'b0, 1'b0};
                            wen_a43 = {1'b0, 1'b0};
                            wen_a42 = {1'b0, 1'b0};
                            wen_a41 = {1'b0, 1'b0};
                            wen_a40 = {1'b0, 1'b0};
                            wen_a39 = {1'b0, 1'b0};
                            wen_a38 = {1'b0, 1'b0};
                            wen_a37 = {1'b0, 1'b0};
                            wen_a36 = {1'b0, wen};
                            wen_a35 = {1'b0, wen};
                        wen_a34 = {1'b0, wen};
                        wen_a33 = {1'b0, wen};
                        wen_a32 = {1'b0, wen};
                        wen_a31 = {1'b0, wen};
                        wen_a30 = {1'b0, wen};
                        wen_a29 = {1'b0, wen};
                        wen_a28 = {1'b0, wen};
                        wen_a27 = {1'b0, wen};
                        wen_a26 = {1'b0, wen};
                        wen_a25 = {1'b0, wen};
                        wen_a24 = {1'b0, wen};
                        wen_a23 = {1'b0, wen};
                        wen_a22 = {1'b0, wen};
                        wen_a21 = {1'b0, wen};
                        wen_a20 = {1'b0, wen};
                        wen_a19 = {1'b0, wen};
                        wen_a18 = {1'b0, wen};
                        wen_a17 = {1'b0, wen};
                        wen_a16 = {1'b0, wen};
                        wen_a15 = {1'b0, wen};
                        wen_a14 = {1'b0, wen};
                        wen_a13 = {1'b0, wen};
                        wen_a12 = {1'b0, wen};
                        wen_a11 = {1'b0, wen};
                        wen_a10 = {1'b0, wen};
                        wen_a9 = {1'b0, wen};
                        wen_a8 = {1'b0, wen};
                        wen_a7 = {1'b0, wen};
                        wen_a6 = {1'b0, wen};
                        wen_a5 = {1'b0, wen};
                        wen_a4 = {1'b0, 1'b0};
                        wen_a3 = {1'b0, 1'b0};
                        wen_a2 = {1'b0, 1'b0};
                        wen_a1 = {1'b0, 1'b0};
                        wen_a0 = {1'b0, 1'b0};
                        wen_b0 = {1'b0, 1'b0};
                    end

                     7'b1000000, 7'b1000001, 7'b1000010, 7'b1000011 : begin
                        wen_a68 = {1'b0, 1'b0};
                        wen_a67 = {1'b0, 1'b0};
                        wen_a66 = {1'b0, 1'b0};
                        wen_a65 = {1'b0, 1'b0};
                        wen_a64 = {1'b0, 1'b0};
                        wen_a63 = {1'b0, 1'b0};
                        wen_a62 = {1'b0, 1'b0};
                        wen_a61 = {1'b0, 1'b0};
                        wen_a60 = {1'b0, 1'b0};
                        wen_a59 = {1'b0, 1'b0};
                        wen_a58 = {1'b0, 1'b0};
                        wen_a57 = {1'b0, 1'b0};
                        wen_a56 = {1'b0, 1'b0};
                        wen_a55 = {1'b0, 1'b0};
                        wen_a54 = {1'b0, 1'b0};
                        wen_a53 = {1'b0, 1'b0};
                        wen_a52 = {1'b0, 1'b0};
                        wen_a51 = {1'b0, 1'b0};
                        wen_a50 = {1'b0, 1'b0};
                        wen_a49 = {1'b0, 1'b0};
                        wen_a48 = {1'b0, 1'b0};
                        wen_a47 = {1'b0, 1'b0};
                        wen_a46 = {1'b0, 1'b0};
                        wen_a45 = {1'b0, 1'b0};
                        wen_a44 = {1'b0, 1'b0};
                        wen_a43 = {1'b0, 1'b0};
                        wen_a42 = {1'b0, 1'b0};
                        wen_a41 = {1'b0, 1'b0};
                        wen_a40 = {1'b0, 1'b0};
                        wen_a39 = {1'b0, 1'b0};
                        wen_a38 = {1'b0, 1'b0};
                        wen_a37 = {1'b0, 1'b0};
                        wen_a36 = {1'b0, 1'b0};
                        wen_a35 = {1'b0, 1'b0};
                        wen_a34 = {1'b0, 1'b0};
                        wen_a33 = {1'b0, 1'b0};
                        wen_a32 = {1'b0, 1'b0};
                        wen_a31 = {1'b0, 1'b0};
                        wen_a30 = {1'b0, 1'b0};
                        wen_a29 = {1'b0, 1'b0};
                        wen_a28 = {1'b0, 1'b0};
                        wen_a27 = {1'b0, 1'b0};
                        wen_a26 = {1'b0, 1'b0};
                        wen_a25 = {1'b0, 1'b0};
                        wen_a24 = {1'b0, 1'b0};
                        wen_a23 = {1'b0, 1'b0};
                        wen_a22 = {1'b0, 1'b0};
                        wen_a21 = {1'b0, 1'b0};
                        wen_a20 = {1'b0, 1'b0};
                        wen_a19 = {1'b0, 1'b0};
                        wen_a18 = {1'b0, 1'b0};
                        wen_a17 = {1'b0, 1'b0};
                        wen_a16 = {1'b0, 1'b0};
                        wen_a15 = {1'b0, 1'b0};
                        wen_a14 = {1'b0, 1'b0};
                        wen_a13 = {1'b0, 1'b0};
                        wen_a12 = {1'b0, 1'b0};
                        wen_a11 = {1'b0, 1'b0};
                        wen_a10 = {1'b0, 1'b0};
                        wen_a9 = {1'b0, 1'b0};
                        wen_a8 = {1'b0, 1'b0};
                        wen_a7 = {1'b0, 1'b0};
                        wen_a6 = {1'b0, 1'b0};
                        wen_a5 = {1'b0, 1'b0};
                        wen_a4 = {1'b0, wen};
                        wen_a3 = {1'b0, wen};
                        wen_a2 = {1'b0, wen};
                        wen_a1 = {1'b0, wen};
                        wen_a0 = {1'b0, 1'b0};
                        wen_b0 = {1'b0, 1'b0};
                    end
                    7'b1000100 : begin
                        wen_a68 = {1'b0, 1'b0};
                        wen_a67 = {1'b0, 1'b0};
                        wen_a66 = {1'b0, 1'b0};
                        wen_a65 = {1'b0, 1'b0};
                        wen_a64 = {1'b0, 1'b0};
                        wen_a63 = {1'b0, 1'b0};
                        wen_a62 = {1'b0, 1'b0};
                        wen_a61 = {1'b0, 1'b0};
                        wen_a60 = {1'b0, 1'b0};
                        wen_a59 = {1'b0, 1'b0};
                        wen_a58 = {1'b0, 1'b0};
                        wen_a57 = {1'b0, 1'b0};
                        wen_a56 = {1'b0, 1'b0};
                        wen_a55 = {1'b0, 1'b0};
                        wen_a54 = {1'b0, 1'b0};
                        wen_a53 = {1'b0, 1'b0};
                        wen_a52 = {1'b0, 1'b0};
                        wen_a51 = {1'b0, 1'b0};
                        wen_a50 = {1'b0, 1'b0};
                        wen_a49 = {1'b0, 1'b0};
                        wen_a48 = {1'b0, 1'b0};
                        wen_a47 = {1'b0, 1'b0};
                        wen_a46 = {1'b0, 1'b0};
                        wen_a45 = {1'b0, 1'b0};
                        wen_a44 = {1'b0, 1'b0};
                        wen_a43 = {1'b0, 1'b0};
                        wen_a42 = {1'b0, 1'b0};
                        wen_a41 = {1'b0, 1'b0};
                        wen_a40 = {1'b0, 1'b0};
                        wen_a39 = {1'b0, 1'b0};
                        wen_a38 = {1'b0, 1'b0};
                        wen_a37 = {1'b0, 1'b0};
                        wen_a36 = {1'b0, 1'b0};
                        wen_a35 = {1'b0, 1'b0};
                        wen_a34 = {1'b0, 1'b0};
                        wen_a33 = {1'b0, 1'b0};
                        wen_a32 = {1'b0, 1'b0};
                        wen_a31 = {1'b0, 1'b0};
                        wen_a30 = {1'b0, 1'b0};
                        wen_a29 = {1'b0, 1'b0};
                        wen_a28 = {1'b0, 1'b0};
                        wen_a27 = {1'b0, 1'b0};
                        wen_a26 = {1'b0, 1'b0};
                        wen_a25 = {1'b0, 1'b0};
                        wen_a24 = {1'b0, 1'b0};
                        wen_a23 = {1'b0, 1'b0};
                        wen_a22 = {1'b0, 1'b0};
                        wen_a21 = {1'b0, 1'b0};
                        wen_a20 = {1'b0, 1'b0};
                        wen_a19 = {1'b0, 1'b0};
                        wen_a18 = {1'b0, 1'b0};
                        wen_a17 = {1'b0, 1'b0};
                        wen_a16 = {1'b0, 1'b0};
                        wen_a15 = {1'b0, 1'b0};
                        wen_a14 = {1'b0, 1'b0};
                        wen_a13 = {1'b0, 1'b0};
                        wen_a12 = {1'b0, 1'b0};
                        wen_a11 = {1'b0, 1'b0};
                        wen_a10 = {1'b0, 1'b0};
                        wen_a9 = {1'b0, 1'b0};
                        wen_a8 = {1'b0, 1'b0};
                        wen_a7 = {1'b0, 1'b0};
                        wen_a6 = {1'b0, 1'b0};
                        wen_a5 = {1'b0, 1'b0};
                        wen_a4 = {1'b0, 1'b0};
                        wen_a3 = {1'b0, 1'b0};
                        wen_a2 = {1'b0, 1'b0};
                        wen_a1 = {1'b0, 1'b0};
                        wen_a0 = {wen,  wen};
                        wen_b0 = {wen,  wen};
                    end
                    default : begin
                        wen_a68 = {1'b0, 1'b0};
                        wen_a67 = {1'b0, 1'b0};
                        wen_a66 = {1'b0, 1'b0};
                        wen_a65 = {1'b0, 1'b0};
                        wen_a64 = {1'b0, 1'b0};
                        wen_a63 = {1'b0, 1'b0};
                        wen_a62 = {1'b0, 1'b0};
                        wen_a61 = {1'b0, 1'b0};
                        wen_a60 = {1'b0, 1'b0};
                        wen_a59 = {1'b0, 1'b0};
                        wen_a58 = {1'b0, 1'b0};
                        wen_a57 = {1'b0, 1'b0};
                        wen_a56 = {1'b0, 1'b0};
                        wen_a55 = {1'b0, 1'b0};
                        wen_a54 = {1'b0, 1'b0};
                        wen_a53 = {1'b0, 1'b0};
                        wen_a52 = {1'b0, 1'b0};
                        wen_a51 = {1'b0, 1'b0};
                        wen_a50 = {1'b0, 1'b0};
                        wen_a49 = {1'b0, 1'b0};
                        wen_a48 = {1'b0, 1'b0};
                        wen_a47 = {1'b0, 1'b0};
                        wen_a46 = {1'b0, 1'b0};
                        wen_a45 = {1'b0, 1'b0};
                        wen_a44 = {1'b0, 1'b0};
                        wen_a43 = {1'b0, 1'b0};
                        wen_a42 = {1'b0, 1'b0};
                        wen_a41 = {1'b0, 1'b0};
                        wen_a40 = {1'b0, 1'b0};
                        wen_a39 = {1'b0, 1'b0};
                        wen_a38 = {1'b0, 1'b0};
                        wen_a37 = {1'b0, 1'b0};
                        wen_a36 = {1'b0, 1'b0};
                        wen_a35 = {1'b0, 1'b0};
                        wen_a34 = {1'b0, 1'b0};
                        wen_a33 = {1'b0, 1'b0};
                        wen_a32 = {1'b0, 1'b0};
                        wen_a31 = {1'b0, 1'b0};
                        wen_a30 = {1'b0, 1'b0};
                        wen_a29 = {1'b0, 1'b0};
                        wen_a28 = {1'b0, 1'b0};
                        wen_a27 = {1'b0, 1'b0};
                        wen_a26 = {1'b0, 1'b0};
                        wen_a25 = {1'b0, 1'b0};
                        wen_a24 = {1'b0, 1'b0};
                        wen_a23 = {1'b0, 1'b0};
                        wen_a22 = {1'b0, 1'b0};
                        wen_a21 = {1'b0, 1'b0};
                        wen_a20 = {1'b0, 1'b0};
                        wen_a19 = {1'b0, 1'b0};
                        wen_a18 = {1'b0, 1'b0};
                        wen_a17 = {1'b0, 1'b0};
                        wen_a16 = {1'b0, 1'b0};
                        wen_a15 = {1'b0, 1'b0};
                        wen_a14 = {1'b0, 1'b0};
                        wen_a13 = {1'b0, 1'b0};
                        wen_a12 = {1'b0, 1'b0};
                        wen_a11 = {1'b0, 1'b0};
                        wen_a10 = {1'b0, 1'b0};
                        wen_a9 = {1'b0, 1'b0};
                        wen_a8 = {1'b0, 1'b0};
                        wen_a7 = {1'b0, 1'b0};
                        wen_a6 = {1'b0, 1'b0};
                        wen_a5 = {1'b0, 1'b0};
                        wen_a4 = {1'b0, 1'b0};
                        wen_a3 = {1'b0, 1'b0};
                        wen_a2 = {1'b0, 1'b0};
                        wen_a1 = {1'b0, 1'b0};
                        wen_a0 = {1'b0, 1'b0};
                        wen_b0 = {1'b0, 1'b0};
                    end
               endcase // case (writeAddr[15:9])

                case (ckRdAddr[15:9])

                       7'b0000000, 7'b0000001, 7'b0000010, 7'b0000011,
                         7'b0000100, 7'b0000101, 7'b0000110, 7'b0000111,
                         7'b0001000, 7'b0001001, 7'b0001010, 7'b0001011,
                         7'b0001100, 7'b0001101, 7'b0001110, 7'b0001111,
                         7'b0010000, 7'b0010001, 7'b0010010, 7'b0010011,
                         7'b0010100, 7'b0010101, 7'b0010110, 7'b0010111,
                         7'b0011000, 7'b0011001, 7'b0011010, 7'b0011011,
                         7'b0011100, 7'b0011101, 7'b0011110, 7'b0011111  : begin
                        readData = {
                                        readData68[0],
                                        readData67[0],
                                        readData66[0],
                                        readData65[0],
                                        readData64[0],
                                        readData63[0],
                                        readData62[0],
                                        readData61[0],
                                        readData60[0],
                                        readData59[0],
                                        readData58[0],
                                        readData57[0],
                                        readData56[0],
                                        readData55[0], 
                                        readData54[0],
                                        readData53[0],
                                        readData52[0],
                                        readData51[0],
                                        readData50[0],
                                        readData49[0],
                                        readData48[0],
                                        readData47[0],
                                        readData46[0],
                                        readData45[0],
                                        readData44[0],
                                        readData43[0],
                                        readData42[0],
                                        readData41[0],
                                        readData40[0],
                                        readData39[0],
                                        readData38[0],
                                        readData37[0]
                        };
                    end
                  7'b0100000, 7'b0100001, 7'b0100010, 7'b0100011,
                    7'b0100100, 7'b0100101, 7'b0100110, 7'b0100111,
                    7'b0101000, 7'b0101001, 7'b0101010, 7'b0101011,
                    7'b0101100, 7'b0101101, 7'b0101110, 7'b0101111,
                    7'b0110000, 7'b0110001, 7'b0110010, 7'b0110011,
                    7'b0110100, 7'b0110101, 7'b0110110, 7'b0110111,             
                    7'b0111000, 7'b0111001, 7'b0111010, 7'b0111011,
                    7'b0111100, 7'b0111101, 7'b0111110, 7'b0111111 : begin
                       readData  =  { readData36[0],
                                        readData35[0],
                                        readData34[0],
                                        readData33[0],
                                        readData32[0],
                                        readData31[0],
                                        readData30[0],
                                        readData29[0],
                                        readData28[0],
                                        readData27[0],
                                        readData26[0],
                                        readData25[0],
                                        readData24[0],
                                        readData23[0],
                                        readData22[0],
                                        readData21[0],
                                        readData20[0],
                                        readData19[0],
                                        readData18[0],
                                        readData17[0],
                                        readData16[0],
                                        readData15[0],
                                        readData14[0],
                                        readData13[0],
                                        readData12[0],
                                        readData11[0],
                                        readData10[0],
                                        readData9[0],
                                        readData8[0],
                                        readData7[0],
                                        readData6[0],
                                        readData5[0]
                                      };                       
                    end                  
                    7'b1000000, 7'b1000001, 7'b1000010, 7'b1000011 : begin
                        readData = {readData4[7:0],readData3[7:0],readData2[7:0],readData1[7:0]};
                    end
                    7'b1000100 : begin
                        readData = {readData0[34:27],readData0[25:18],readData0[16:9],readData0[7:0]};
                    end
                    default : begin
                       readData = 32'b0;
                    end
               endcase // case (ckRdAddr[15:9])                                    
           end // case: 35328

        endcase // case (DEPTH)       
    end // always @ (*)   


    //----------------------------------------------------------------------------------------
    // RAM1K18 blocks
    //----------------------------------------------------------------------------------------
    RAM1K18 block68 (
        .A_DOUT (readData68),           .B_DOUT (),
        .A_CLK (clk),                  .B_CLK (clk), 
        .A_ARST_N (resetn),            .B_ARST_N (resetn), 
        .A_BLK (3'b111),               .B_BLK (3'b111), 
        .A_DIN (writeData68),           .B_DIN (writeData68), 
        .A_ADDR (writeAddr68),          .B_ADDR (writeAddr68), 
        .A_WEN (wen_a68),               .B_WEN (wen_b68),
        .A_DOUT_CLK (1'b1),            .B_DOUT_CLK (1'b1), 
        .A_DOUT_EN (1'b1),             .B_DOUT_EN (1'b1), 
        .A_DOUT_ARST_N (1'b1),         .B_DOUT_ARST_N (1'b1), 
        .A_DOUT_SRST_N (1'b1),         .B_DOUT_SRST_N (1'b1), 
        .A_DOUT_LAT (1'b1),            .B_DOUT_LAT (1'b1),
        .A_WIDTH (width68),             .B_WIDTH (width68), 
        .A_WMODE (1'b0),               .B_WMODE (1'b0),
        .A_EN (1'b1),                  .B_EN (1'b1),
        .BUSY (lsram_512_BUSY_68),
        .SII_LOCK (1'b0)
    );

    RAM1K18 block67 (
        .A_DOUT (readData67),           .B_DOUT (),
        .A_CLK (clk),                  .B_CLK (clk), 
        .A_ARST_N (resetn),            .B_ARST_N (resetn), 
        .A_BLK (3'b111),               .B_BLK (3'b111), 
        .A_DIN (writeData67),           .B_DIN (writeData67), 
        .A_ADDR (writeAddr67),          .B_ADDR (writeAddr67), 
        .A_WEN (wen_a67),               .B_WEN (wen_b67),
        .A_DOUT_CLK (1'b1),            .B_DOUT_CLK (1'b1), 
        .A_DOUT_EN (1'b1),             .B_DOUT_EN (1'b1), 
        .A_DOUT_ARST_N (1'b1),         .B_DOUT_ARST_N (1'b1), 
        .A_DOUT_SRST_N (1'b1),         .B_DOUT_SRST_N (1'b1), 
        .A_DOUT_LAT (1'b1),            .B_DOUT_LAT (1'b1),
        .A_WIDTH (width67),             .B_WIDTH (width67), 
        .A_WMODE (1'b0),               .B_WMODE (1'b0),
        .A_EN (1'b1),                  .B_EN (1'b1),
        .BUSY (lsram_512_BUSY_67),
        .SII_LOCK (1'b0)
    );

    RAM1K18 block66 (
        .A_DOUT (readData66),           .B_DOUT (),
        .A_CLK (clk),                  .B_CLK (clk), 
        .A_ARST_N (resetn),            .B_ARST_N (resetn), 
        .A_BLK (3'b111),               .B_BLK (3'b111), 
        .A_DIN (writeData66),           .B_DIN (writeData66), 
        .A_ADDR (writeAddr66),          .B_ADDR (writeAddr66), 
        .A_WEN (wen_a66),               .B_WEN (wen_b66),
        .A_DOUT_CLK (1'b1),            .B_DOUT_CLK (1'b1), 
        .A_DOUT_EN (1'b1),             .B_DOUT_EN (1'b1), 
        .A_DOUT_ARST_N (1'b1),         .B_DOUT_ARST_N (1'b1), 
        .A_DOUT_SRST_N (1'b1),         .B_DOUT_SRST_N (1'b1), 
        .A_DOUT_LAT (1'b1),            .B_DOUT_LAT (1'b1),
        .A_WIDTH (width66),             .B_WIDTH (width66), 
        .A_WMODE (1'b0),               .B_WMODE (1'b0),
        .A_EN (1'b1),                  .B_EN (1'b1),
        .BUSY (lsram_512_BUSY_66),
        .SII_LOCK (1'b0)
    );

    RAM1K18 block65 (
        .A_DOUT (readData65),           .B_DOUT (),
        .A_CLK (clk),                  .B_CLK (clk), 
        .A_ARST_N (resetn),            .B_ARST_N (resetn), 
        .A_BLK (3'b111),               .B_BLK (3'b111), 
        .A_DIN (writeData65),           .B_DIN (writeData65), 
        .A_ADDR (writeAddr65),          .B_ADDR (writeAddr65), 
        .A_WEN (wen_a65),               .B_WEN (wen_b65),
        .A_DOUT_CLK (1'b1),            .B_DOUT_CLK (1'b1), 
        .A_DOUT_EN (1'b1),             .B_DOUT_EN (1'b1), 
        .A_DOUT_ARST_N (1'b1),         .B_DOUT_ARST_N (1'b1), 
        .A_DOUT_SRST_N (1'b1),         .B_DOUT_SRST_N (1'b1), 
        .A_DOUT_LAT (1'b1),            .B_DOUT_LAT (1'b1),
        .A_WIDTH (width65),             .B_WIDTH (width65), 
        .A_WMODE (1'b0),               .B_WMODE (1'b0),
        .A_EN (1'b1),                  .B_EN (1'b1),
        .BUSY (lsram_512_BUSY_65),
        .SII_LOCK (1'b0)
    );

    RAM1K18 block64 (
        .A_DOUT (readData64),           .B_DOUT (),
        .A_CLK (clk),                  .B_CLK (clk), 
        .A_ARST_N (resetn),            .B_ARST_N (resetn), 
        .A_BLK (3'b111),               .B_BLK (3'b111), 
        .A_DIN (writeData64),           .B_DIN (writeData64), 
        .A_ADDR (writeAddr64),          .B_ADDR (writeAddr64), 
        .A_WEN (wen_a64),               .B_WEN (wen_b64),
        .A_DOUT_CLK (1'b1),            .B_DOUT_CLK (1'b1), 
        .A_DOUT_EN (1'b1),             .B_DOUT_EN (1'b1), 
        .A_DOUT_ARST_N (1'b1),         .B_DOUT_ARST_N (1'b1), 
        .A_DOUT_SRST_N (1'b1),         .B_DOUT_SRST_N (1'b1), 
        .A_DOUT_LAT (1'b1),            .B_DOUT_LAT (1'b1),
        .A_WIDTH (width64),             .B_WIDTH (width64), 
        .A_WMODE (1'b0),               .B_WMODE (1'b0),
        .A_EN (1'b1),                  .B_EN (1'b1),
        .BUSY (lsram_512_BUSY_64),
        .SII_LOCK (1'b0)
    );

    RAM1K18 block63 (
        .A_DOUT (readData63),           .B_DOUT (),
        .A_CLK (clk),                  .B_CLK (clk), 
        .A_ARST_N (resetn),            .B_ARST_N (resetn), 
        .A_BLK (3'b111),               .B_BLK (3'b111), 
        .A_DIN (writeData63),           .B_DIN (writeData63), 
        .A_ADDR (writeAddr63),          .B_ADDR (writeAddr63), 
        .A_WEN (wen_a63),               .B_WEN (wen_b63),
        .A_DOUT_CLK (1'b1),            .B_DOUT_CLK (1'b1), 
        .A_DOUT_EN (1'b1),             .B_DOUT_EN (1'b1), 
        .A_DOUT_ARST_N (1'b1),         .B_DOUT_ARST_N (1'b1), 
        .A_DOUT_SRST_N (1'b1),         .B_DOUT_SRST_N (1'b1), 
        .A_DOUT_LAT (1'b1),            .B_DOUT_LAT (1'b1),
        .A_WIDTH (width63),             .B_WIDTH (width63), 
        .A_WMODE (1'b0),               .B_WMODE (1'b0),
        .A_EN (1'b1),                  .B_EN (1'b1),
        .BUSY (lsram_512_BUSY_63),
        .SII_LOCK (1'b0)
    );

    RAM1K18 block62 (
        .A_DOUT (readData62),           .B_DOUT (),
        .A_CLK (clk),                  .B_CLK (clk), 
        .A_ARST_N (resetn),            .B_ARST_N (resetn), 
        .A_BLK (3'b111),               .B_BLK (3'b111), 
        .A_DIN (writeData62),           .B_DIN (writeData62), 
        .A_ADDR (writeAddr62),          .B_ADDR (writeAddr62), 
        .A_WEN (wen_a62),               .B_WEN (wen_b62),
        .A_DOUT_CLK (1'b1),            .B_DOUT_CLK (1'b1), 
        .A_DOUT_EN (1'b1),             .B_DOUT_EN (1'b1), 
        .A_DOUT_ARST_N (1'b1),         .B_DOUT_ARST_N (1'b1), 
        .A_DOUT_SRST_N (1'b1),         .B_DOUT_SRST_N (1'b1), 
        .A_DOUT_LAT (1'b1),            .B_DOUT_LAT (1'b1),
        .A_WIDTH (width62),             .B_WIDTH (width62), 
        .A_WMODE (1'b0),               .B_WMODE (1'b0),
        .A_EN (1'b1),                  .B_EN (1'b1),
        .BUSY (lsram_512_BUSY_62),
        .SII_LOCK (1'b0)
    );

    RAM1K18 block61 (
        .A_DOUT (readData61),           .B_DOUT (),
        .A_CLK (clk),                  .B_CLK (clk), 
        .A_ARST_N (resetn),            .B_ARST_N (resetn), 
        .A_BLK (3'b111),               .B_BLK (3'b111), 
        .A_DIN (writeData61),           .B_DIN (writeData61), 
        .A_ADDR (writeAddr61),          .B_ADDR (writeAddr61), 
        .A_WEN (wen_a61),               .B_WEN (wen_b61),
        .A_DOUT_CLK (1'b1),            .B_DOUT_CLK (1'b1), 
        .A_DOUT_EN (1'b1),             .B_DOUT_EN (1'b1), 
        .A_DOUT_ARST_N (1'b1),         .B_DOUT_ARST_N (1'b1), 
        .A_DOUT_SRST_N (1'b1),         .B_DOUT_SRST_N (1'b1), 
        .A_DOUT_LAT (1'b1),            .B_DOUT_LAT (1'b1),
        .A_WIDTH (width61),             .B_WIDTH (width61), 
        .A_WMODE (1'b0),               .B_WMODE (1'b0),
        .A_EN (1'b1),                  .B_EN (1'b1),
        .BUSY (lsram_512_BUSY_61),
        .SII_LOCK (1'b0)
    );

    RAM1K18 block60 (
        .A_DOUT (readData60),           .B_DOUT (),
        .A_CLK (clk),                  .B_CLK (clk), 
        .A_ARST_N (resetn),            .B_ARST_N (resetn), 
        .A_BLK (3'b111),               .B_BLK (3'b111), 
        .A_DIN (writeData60),           .B_DIN (writeData60), 
        .A_ADDR (writeAddr60),          .B_ADDR (writeAddr60), 
        .A_WEN (wen_a60),               .B_WEN (wen_b60),
        .A_DOUT_CLK (1'b1),            .B_DOUT_CLK (1'b1), 
        .A_DOUT_EN (1'b1),             .B_DOUT_EN (1'b1), 
        .A_DOUT_ARST_N (1'b1),         .B_DOUT_ARST_N (1'b1), 
        .A_DOUT_SRST_N (1'b1),         .B_DOUT_SRST_N (1'b1), 
        .A_DOUT_LAT (1'b1),            .B_DOUT_LAT (1'b1),
        .A_WIDTH (width60),             .B_WIDTH (width60), 
        .A_WMODE (1'b0),               .B_WMODE (1'b0),
        .A_EN (1'b1),                  .B_EN (1'b1),
        .BUSY (lsram_512_BUSY_60),
        .SII_LOCK (1'b0)
    );

    RAM1K18 block59 (
        .A_DOUT (readData59),           .B_DOUT (),
        .A_CLK (clk),                  .B_CLK (clk), 
        .A_ARST_N (resetn),            .B_ARST_N (resetn), 
        .A_BLK (3'b111),               .B_BLK (3'b111), 
        .A_DIN (writeData59),           .B_DIN (writeData59), 
        .A_ADDR (writeAddr59),          .B_ADDR (writeAddr59), 
        .A_WEN (wen_a59),               .B_WEN (wen_b59),
        .A_DOUT_CLK (1'b1),            .B_DOUT_CLK (1'b1), 
        .A_DOUT_EN (1'b1),             .B_DOUT_EN (1'b1), 
        .A_DOUT_ARST_N (1'b1),         .B_DOUT_ARST_N (1'b1), 
        .A_DOUT_SRST_N (1'b1),         .B_DOUT_SRST_N (1'b1), 
        .A_DOUT_LAT (1'b1),            .B_DOUT_LAT (1'b1),
        .A_WIDTH (width59),             .B_WIDTH (width59), 
        .A_WMODE (1'b0),               .B_WMODE (1'b0),
        .A_EN (1'b1),                  .B_EN (1'b1),
        .BUSY (lsram_512_BUSY_59),
        .SII_LOCK (1'b0)
    );

    RAM1K18 block58 (
        .A_DOUT (readData58),           .B_DOUT (),
        .A_CLK (clk),                  .B_CLK (clk), 
        .A_ARST_N (resetn),            .B_ARST_N (resetn), 
        .A_BLK (3'b111),               .B_BLK (3'b111), 
        .A_DIN (writeData58),           .B_DIN (writeData58), 
        .A_ADDR (writeAddr58),          .B_ADDR (writeAddr58), 
        .A_WEN (wen_a58),               .B_WEN (wen_b58),
        .A_DOUT_CLK (1'b1),            .B_DOUT_CLK (1'b1), 
        .A_DOUT_EN (1'b1),             .B_DOUT_EN (1'b1), 
        .A_DOUT_ARST_N (1'b1),         .B_DOUT_ARST_N (1'b1), 
        .A_DOUT_SRST_N (1'b1),         .B_DOUT_SRST_N (1'b1), 
        .A_DOUT_LAT (1'b1),            .B_DOUT_LAT (1'b1),
        .A_WIDTH (width58),             .B_WIDTH (width58), 
        .A_WMODE (1'b0),               .B_WMODE (1'b0),
        .A_EN (1'b1),                  .B_EN (1'b1),
        .BUSY (lsram_512_BUSY_58),
        .SII_LOCK (1'b0)
    );

    RAM1K18 block57 (
        .A_DOUT (readData57),           .B_DOUT (),
        .A_CLK (clk),                  .B_CLK (clk), 
        .A_ARST_N (resetn),            .B_ARST_N (resetn), 
        .A_BLK (3'b111),               .B_BLK (3'b111), 
        .A_DIN (writeData57),           .B_DIN (writeData57), 
        .A_ADDR (writeAddr57),          .B_ADDR (writeAddr57), 
        .A_WEN (wen_a57),               .B_WEN (wen_b57),
        .A_DOUT_CLK (1'b1),            .B_DOUT_CLK (1'b1), 
        .A_DOUT_EN (1'b1),             .B_DOUT_EN (1'b1), 
        .A_DOUT_ARST_N (1'b1),         .B_DOUT_ARST_N (1'b1), 
        .A_DOUT_SRST_N (1'b1),         .B_DOUT_SRST_N (1'b1), 
        .A_DOUT_LAT (1'b1),            .B_DOUT_LAT (1'b1),
        .A_WIDTH (width57),             .B_WIDTH (width57), 
        .A_WMODE (1'b0),               .B_WMODE (1'b0),
        .A_EN (1'b1),                  .B_EN (1'b1),
        .BUSY (lsram_512_BUSY_57),
        .SII_LOCK (1'b0)
    );

    RAM1K18 block56 (
        .A_DOUT (readData56),           .B_DOUT (),
        .A_CLK (clk),                  .B_CLK (clk), 
        .A_ARST_N (resetn),            .B_ARST_N (resetn), 
        .A_BLK (3'b111),               .B_BLK (3'b111), 
        .A_DIN (writeData56),           .B_DIN (writeData56), 
        .A_ADDR (writeAddr56),          .B_ADDR (writeAddr56), 
        .A_WEN (wen_a56),               .B_WEN (wen_b56),
        .A_DOUT_CLK (1'b1),            .B_DOUT_CLK (1'b1), 
        .A_DOUT_EN (1'b1),             .B_DOUT_EN (1'b1), 
        .A_DOUT_ARST_N (1'b1),         .B_DOUT_ARST_N (1'b1), 
        .A_DOUT_SRST_N (1'b1),         .B_DOUT_SRST_N (1'b1), 
        .A_DOUT_LAT (1'b1),            .B_DOUT_LAT (1'b1),
        .A_WIDTH (width56),             .B_WIDTH (width56), 
        .A_WMODE (1'b0),               .B_WMODE (1'b0),
        .A_EN (1'b1),                  .B_EN (1'b1),
        .BUSY (lsram_512_BUSY_56),
        .SII_LOCK (1'b0)
    );

    RAM1K18 block55 (
        .A_DOUT (readData55),           .B_DOUT (),
        .A_CLK (clk),                  .B_CLK (clk), 
        .A_ARST_N (resetn),            .B_ARST_N (resetn), 
        .A_BLK (3'b111),               .B_BLK (3'b111), 
        .A_DIN (writeData55),           .B_DIN (writeData55), 
        .A_ADDR (writeAddr55),          .B_ADDR (writeAddr55), 
        .A_WEN (wen_a55),               .B_WEN (wen_b55),
        .A_DOUT_CLK (1'b1),            .B_DOUT_CLK (1'b1), 
        .A_DOUT_EN (1'b1),             .B_DOUT_EN (1'b1), 
        .A_DOUT_ARST_N (1'b1),         .B_DOUT_ARST_N (1'b1), 
        .A_DOUT_SRST_N (1'b1),         .B_DOUT_SRST_N (1'b1), 
        .A_DOUT_LAT (1'b1),            .B_DOUT_LAT (1'b1),
        .A_WIDTH (width55),             .B_WIDTH (width55), 
        .A_WMODE (1'b0),               .B_WMODE (1'b0),
        .A_EN (1'b1),                  .B_EN (1'b1),
        .BUSY (lsram_512_BUSY_55),
        .SII_LOCK (1'b0)
    );

    RAM1K18 block54 (
        .A_DOUT (readData54),           .B_DOUT (),
        .A_CLK (clk),                  .B_CLK (clk), 
        .A_ARST_N (resetn),            .B_ARST_N (resetn), 
        .A_BLK (3'b111),               .B_BLK (3'b111), 
        .A_DIN (writeData54),           .B_DIN (writeData54), 
        .A_ADDR (writeAddr54),          .B_ADDR (writeAddr54), 
        .A_WEN (wen_a54),               .B_WEN (wen_b54),
        .A_DOUT_CLK (1'b1),            .B_DOUT_CLK (1'b1), 
        .A_DOUT_EN (1'b1),             .B_DOUT_EN (1'b1), 
        .A_DOUT_ARST_N (1'b1),         .B_DOUT_ARST_N (1'b1), 
        .A_DOUT_SRST_N (1'b1),         .B_DOUT_SRST_N (1'b1), 
        .A_DOUT_LAT (1'b1),            .B_DOUT_LAT (1'b1),
        .A_WIDTH (width54),             .B_WIDTH (width54), 
        .A_WMODE (1'b0),               .B_WMODE (1'b0),
        .A_EN (1'b1),                  .B_EN (1'b1),
        .BUSY (lsram_512_BUSY_54),
        .SII_LOCK (1'b0)
    );

    RAM1K18 block53 (
        .A_DOUT (readData53),           .B_DOUT (),
        .A_CLK (clk),                  .B_CLK (clk), 
        .A_ARST_N (resetn),            .B_ARST_N (resetn), 
        .A_BLK (3'b111),               .B_BLK (3'b111), 
        .A_DIN (writeData53),           .B_DIN (writeData53), 
        .A_ADDR (writeAddr53),          .B_ADDR (writeAddr53), 
        .A_WEN (wen_a53),               .B_WEN (wen_b53),
        .A_DOUT_CLK (1'b1),            .B_DOUT_CLK (1'b1), 
        .A_DOUT_EN (1'b1),             .B_DOUT_EN (1'b1), 
        .A_DOUT_ARST_N (1'b1),         .B_DOUT_ARST_N (1'b1), 
        .A_DOUT_SRST_N (1'b1),         .B_DOUT_SRST_N (1'b1), 
        .A_DOUT_LAT (1'b1),            .B_DOUT_LAT (1'b1),
        .A_WIDTH (width53),             .B_WIDTH (width53), 
        .A_WMODE (1'b0),               .B_WMODE (1'b0),
        .A_EN (1'b1),                  .B_EN (1'b1),
        .BUSY (lsram_512_BUSY_53),
        .SII_LOCK (1'b0)
    );

    RAM1K18 block52 (
        .A_DOUT (readData52),           .B_DOUT (),
        .A_CLK (clk),                  .B_CLK (clk), 
        .A_ARST_N (resetn),            .B_ARST_N (resetn), 
        .A_BLK (3'b111),               .B_BLK (3'b111), 
        .A_DIN (writeData52),           .B_DIN (writeData52), 
        .A_ADDR (writeAddr52),          .B_ADDR (writeAddr52), 
        .A_WEN (wen_a52),               .B_WEN (wen_b52),
        .A_DOUT_CLK (1'b1),            .B_DOUT_CLK (1'b1), 
        .A_DOUT_EN (1'b1),             .B_DOUT_EN (1'b1), 
        .A_DOUT_ARST_N (1'b1),         .B_DOUT_ARST_N (1'b1), 
        .A_DOUT_SRST_N (1'b1),         .B_DOUT_SRST_N (1'b1), 
        .A_DOUT_LAT (1'b1),            .B_DOUT_LAT (1'b1),
        .A_WIDTH (width52),             .B_WIDTH (width52), 
        .A_WMODE (1'b0),               .B_WMODE (1'b0),
        .A_EN (1'b1),                  .B_EN (1'b1),
        .BUSY (lsram_512_BUSY_52),
        .SII_LOCK (1'b0)
    );

    RAM1K18 block51 (
        .A_DOUT (readData51),           .B_DOUT (),
        .A_CLK (clk),                  .B_CLK (clk), 
        .A_ARST_N (resetn),            .B_ARST_N (resetn), 
        .A_BLK (3'b111),               .B_BLK (3'b111), 
        .A_DIN (writeData51),           .B_DIN (writeData51), 
        .A_ADDR (writeAddr51),          .B_ADDR (writeAddr51), 
        .A_WEN (wen_a51),               .B_WEN (wen_b51),
        .A_DOUT_CLK (1'b1),            .B_DOUT_CLK (1'b1), 
        .A_DOUT_EN (1'b1),             .B_DOUT_EN (1'b1), 
        .A_DOUT_ARST_N (1'b1),         .B_DOUT_ARST_N (1'b1), 
        .A_DOUT_SRST_N (1'b1),         .B_DOUT_SRST_N (1'b1), 
        .A_DOUT_LAT (1'b1),            .B_DOUT_LAT (1'b1),
        .A_WIDTH (width51),             .B_WIDTH (width51), 
        .A_WMODE (1'b0),               .B_WMODE (1'b0),
        .A_EN (1'b1),                  .B_EN (1'b1),
        .BUSY (lsram_512_BUSY_51),
        .SII_LOCK (1'b0)
    );

    RAM1K18 block50 (
        .A_DOUT (readData50),           .B_DOUT (),
        .A_CLK (clk),                  .B_CLK (clk), 
        .A_ARST_N (resetn),            .B_ARST_N (resetn), 
        .A_BLK (3'b111),               .B_BLK (3'b111), 
        .A_DIN (writeData50),           .B_DIN (writeData50), 
        .A_ADDR (writeAddr50),          .B_ADDR (writeAddr50), 
        .A_WEN (wen_a50),               .B_WEN (wen_b50),
        .A_DOUT_CLK (1'b1),            .B_DOUT_CLK (1'b1), 
        .A_DOUT_EN (1'b1),             .B_DOUT_EN (1'b1), 
        .A_DOUT_ARST_N (1'b1),         .B_DOUT_ARST_N (1'b1), 
        .A_DOUT_SRST_N (1'b1),         .B_DOUT_SRST_N (1'b1), 
        .A_DOUT_LAT (1'b1),            .B_DOUT_LAT (1'b1),
        .A_WIDTH (width50),             .B_WIDTH (width50), 
        .A_WMODE (1'b0),               .B_WMODE (1'b0),
        .A_EN (1'b1),                  .B_EN (1'b1),
        .BUSY (lsram_512_BUSY_50),
        .SII_LOCK (1'b0)
    );

    RAM1K18 block49 (
        .A_DOUT (readData49),           .B_DOUT (),
        .A_CLK (clk),                  .B_CLK (clk), 
        .A_ARST_N (resetn),            .B_ARST_N (resetn), 
        .A_BLK (3'b111),               .B_BLK (3'b111), 
        .A_DIN (writeData49),           .B_DIN (writeData49), 
        .A_ADDR (writeAddr49),          .B_ADDR (writeAddr49), 
        .A_WEN (wen_a49),               .B_WEN (wen_b49),
        .A_DOUT_CLK (1'b1),            .B_DOUT_CLK (1'b1), 
        .A_DOUT_EN (1'b1),             .B_DOUT_EN (1'b1), 
        .A_DOUT_ARST_N (1'b1),         .B_DOUT_ARST_N (1'b1), 
        .A_DOUT_SRST_N (1'b1),         .B_DOUT_SRST_N (1'b1), 
        .A_DOUT_LAT (1'b1),            .B_DOUT_LAT (1'b1),
        .A_WIDTH (width49),             .B_WIDTH (width49), 
        .A_WMODE (1'b0),               .B_WMODE (1'b0),
        .A_EN (1'b1),                  .B_EN (1'b1),
        .BUSY (lsram_512_BUSY_49),
        .SII_LOCK (1'b0)
    );

    RAM1K18 block48 (
        .A_DOUT (readData48),           .B_DOUT (),
        .A_CLK (clk),                  .B_CLK (clk), 
        .A_ARST_N (resetn),            .B_ARST_N (resetn), 
        .A_BLK (3'b111),               .B_BLK (3'b111), 
        .A_DIN (writeData48),           .B_DIN (writeData48), 
        .A_ADDR (writeAddr48),          .B_ADDR (writeAddr48), 
        .A_WEN (wen_a48),               .B_WEN (wen_b48),
        .A_DOUT_CLK (1'b1),            .B_DOUT_CLK (1'b1), 
        .A_DOUT_EN (1'b1),             .B_DOUT_EN (1'b1), 
        .A_DOUT_ARST_N (1'b1),         .B_DOUT_ARST_N (1'b1), 
        .A_DOUT_SRST_N (1'b1),         .B_DOUT_SRST_N (1'b1), 
        .A_DOUT_LAT (1'b1),            .B_DOUT_LAT (1'b1),
        .A_WIDTH (width48),             .B_WIDTH (width48), 
        .A_WMODE (1'b0),               .B_WMODE (1'b0),
        .A_EN (1'b1),                  .B_EN (1'b1),
        .BUSY (lsram_512_BUSY_48),
        .SII_LOCK (1'b0)
    );

    RAM1K18 block47 (
        .A_DOUT (readData47),           .B_DOUT (),
        .A_CLK (clk),                  .B_CLK (clk), 
        .A_ARST_N (resetn),            .B_ARST_N (resetn), 
        .A_BLK (3'b111),               .B_BLK (3'b111), 
        .A_DIN (writeData47),           .B_DIN (writeData47), 
        .A_ADDR (writeAddr47),          .B_ADDR (writeAddr47), 
        .A_WEN (wen_a47),               .B_WEN (wen_b47),
        .A_DOUT_CLK (1'b1),            .B_DOUT_CLK (1'b1), 
        .A_DOUT_EN (1'b1),             .B_DOUT_EN (1'b1), 
        .A_DOUT_ARST_N (1'b1),         .B_DOUT_ARST_N (1'b1), 
        .A_DOUT_SRST_N (1'b1),         .B_DOUT_SRST_N (1'b1), 
        .A_DOUT_LAT (1'b1),            .B_DOUT_LAT (1'b1),
        .A_WIDTH (width47),             .B_WIDTH (width47), 
        .A_WMODE (1'b0),               .B_WMODE (1'b0),
        .A_EN (1'b1),                  .B_EN (1'b1),
        .BUSY (lsram_512_BUSY_47),
        .SII_LOCK (1'b0)
    );

    RAM1K18 block46 (
        .A_DOUT (readData46),           .B_DOUT (),
        .A_CLK (clk),                  .B_CLK (clk), 
        .A_ARST_N (resetn),            .B_ARST_N (resetn), 
        .A_BLK (3'b111),               .B_BLK (3'b111), 
        .A_DIN (writeData46),           .B_DIN (writeData46), 
        .A_ADDR (writeAddr46),          .B_ADDR (writeAddr46), 
        .A_WEN (wen_a46),               .B_WEN (wen_b46),
        .A_DOUT_CLK (1'b1),            .B_DOUT_CLK (1'b1), 
        .A_DOUT_EN (1'b1),             .B_DOUT_EN (1'b1), 
        .A_DOUT_ARST_N (1'b1),         .B_DOUT_ARST_N (1'b1), 
        .A_DOUT_SRST_N (1'b1),         .B_DOUT_SRST_N (1'b1), 
        .A_DOUT_LAT (1'b1),            .B_DOUT_LAT (1'b1),
        .A_WIDTH (width46),             .B_WIDTH (width46), 
        .A_WMODE (1'b0),               .B_WMODE (1'b0),
        .A_EN (1'b1),                  .B_EN (1'b1),
        .BUSY (lsram_512_BUSY_46),
        .SII_LOCK (1'b0)
    );

    RAM1K18 block45 (
        .A_DOUT (readData45),           .B_DOUT (),
        .A_CLK (clk),                  .B_CLK (clk), 
        .A_ARST_N (resetn),            .B_ARST_N (resetn), 
        .A_BLK (3'b111),               .B_BLK (3'b111), 
        .A_DIN (writeData45),           .B_DIN (writeData45), 
        .A_ADDR (writeAddr45),          .B_ADDR (writeAddr45), 
        .A_WEN (wen_a45),               .B_WEN (wen_b45),
        .A_DOUT_CLK (1'b1),            .B_DOUT_CLK (1'b1), 
        .A_DOUT_EN (1'b1),             .B_DOUT_EN (1'b1), 
        .A_DOUT_ARST_N (1'b1),         .B_DOUT_ARST_N (1'b1), 
        .A_DOUT_SRST_N (1'b1),         .B_DOUT_SRST_N (1'b1), 
        .A_DOUT_LAT (1'b1),            .B_DOUT_LAT (1'b1),
        .A_WIDTH (width45),             .B_WIDTH (width45), 
        .A_WMODE (1'b0),               .B_WMODE (1'b0),
        .A_EN (1'b1),                  .B_EN (1'b1),
        .BUSY (lsram_512_BUSY_45),
        .SII_LOCK (1'b0)
    );

    RAM1K18 block44 (
        .A_DOUT (readData44),           .B_DOUT (),
        .A_CLK (clk),                  .B_CLK (clk), 
        .A_ARST_N (resetn),            .B_ARST_N (resetn), 
        .A_BLK (3'b111),               .B_BLK (3'b111), 
        .A_DIN (writeData44),           .B_DIN (writeData44), 
        .A_ADDR (writeAddr44),          .B_ADDR (writeAddr44), 
        .A_WEN (wen_a44),               .B_WEN (wen_b44),
        .A_DOUT_CLK (1'b1),            .B_DOUT_CLK (1'b1), 
        .A_DOUT_EN (1'b1),             .B_DOUT_EN (1'b1), 
        .A_DOUT_ARST_N (1'b1),         .B_DOUT_ARST_N (1'b1), 
        .A_DOUT_SRST_N (1'b1),         .B_DOUT_SRST_N (1'b1), 
        .A_DOUT_LAT (1'b1),            .B_DOUT_LAT (1'b1),
        .A_WIDTH (width44),             .B_WIDTH (width44), 
        .A_WMODE (1'b0),               .B_WMODE (1'b0),
        .A_EN (1'b1),                  .B_EN (1'b1),
        .BUSY (lsram_512_BUSY_44),
        .SII_LOCK (1'b0)
    );

    RAM1K18 block43 (
        .A_DOUT (readData43),           .B_DOUT (),
        .A_CLK (clk),                  .B_CLK (clk), 
        .A_ARST_N (resetn),            .B_ARST_N (resetn), 
        .A_BLK (3'b111),               .B_BLK (3'b111), 
        .A_DIN (writeData43),           .B_DIN (writeData43), 
        .A_ADDR (writeAddr43),          .B_ADDR (writeAddr43), 
        .A_WEN (wen_a43),               .B_WEN (wen_b43),
        .A_DOUT_CLK (1'b1),            .B_DOUT_CLK (1'b1), 
        .A_DOUT_EN (1'b1),             .B_DOUT_EN (1'b1), 
        .A_DOUT_ARST_N (1'b1),         .B_DOUT_ARST_N (1'b1), 
        .A_DOUT_SRST_N (1'b1),         .B_DOUT_SRST_N (1'b1), 
        .A_DOUT_LAT (1'b1),            .B_DOUT_LAT (1'b1),
        .A_WIDTH (width43),             .B_WIDTH (width43), 
        .A_WMODE (1'b0),               .B_WMODE (1'b0),
        .A_EN (1'b1),                  .B_EN (1'b1),
        .BUSY (lsram_512_BUSY_43),
        .SII_LOCK (1'b0)
    );

    RAM1K18 block42 (
        .A_DOUT (readData42),           .B_DOUT (),
        .A_CLK (clk),                  .B_CLK (clk), 
        .A_ARST_N (resetn),            .B_ARST_N (resetn), 
        .A_BLK (3'b111),               .B_BLK (3'b111), 
        .A_DIN (writeData42),           .B_DIN (writeData42), 
        .A_ADDR (writeAddr42),          .B_ADDR (writeAddr42), 
        .A_WEN (wen_a42),               .B_WEN (wen_b42),
        .A_DOUT_CLK (1'b1),            .B_DOUT_CLK (1'b1), 
        .A_DOUT_EN (1'b1),             .B_DOUT_EN (1'b1), 
        .A_DOUT_ARST_N (1'b1),         .B_DOUT_ARST_N (1'b1), 
        .A_DOUT_SRST_N (1'b1),         .B_DOUT_SRST_N (1'b1), 
        .A_DOUT_LAT (1'b1),            .B_DOUT_LAT (1'b1),
        .A_WIDTH (width42),             .B_WIDTH (width42), 
        .A_WMODE (1'b0),               .B_WMODE (1'b0),
        .A_EN (1'b1),                  .B_EN (1'b1),
        .BUSY (lsram_512_BUSY_42),
        .SII_LOCK (1'b0)
    );

    RAM1K18 block41 (
        .A_DOUT (readData41),           .B_DOUT (),
        .A_CLK (clk),                  .B_CLK (clk), 
        .A_ARST_N (resetn),            .B_ARST_N (resetn), 
        .A_BLK (3'b111),               .B_BLK (3'b111), 
        .A_DIN (writeData41),           .B_DIN (writeData41), 
        .A_ADDR (writeAddr41),          .B_ADDR (writeAddr41), 
        .A_WEN (wen_a41),               .B_WEN (wen_b41),
        .A_DOUT_CLK (1'b1),            .B_DOUT_CLK (1'b1), 
        .A_DOUT_EN (1'b1),             .B_DOUT_EN (1'b1), 
        .A_DOUT_ARST_N (1'b1),         .B_DOUT_ARST_N (1'b1), 
        .A_DOUT_SRST_N (1'b1),         .B_DOUT_SRST_N (1'b1), 
        .A_DOUT_LAT (1'b1),            .B_DOUT_LAT (1'b1),
        .A_WIDTH (width41),             .B_WIDTH (width41), 
        .A_WMODE (1'b0),               .B_WMODE (1'b0),
        .A_EN (1'b1),                  .B_EN (1'b1),
        .BUSY (lsram_512_BUSY_41),
        .SII_LOCK (1'b0)
    );

    RAM1K18 block40 (
        .A_DOUT (readData40),           .B_DOUT (),
        .A_CLK (clk),                  .B_CLK (clk), 
        .A_ARST_N (resetn),            .B_ARST_N (resetn), 
        .A_BLK (3'b111),               .B_BLK (3'b111), 
        .A_DIN (writeData40),           .B_DIN (writeData40), 
        .A_ADDR (writeAddr40),          .B_ADDR (writeAddr40), 
        .A_WEN (wen_a40),               .B_WEN (wen_b40),
        .A_DOUT_CLK (1'b1),            .B_DOUT_CLK (1'b1), 
        .A_DOUT_EN (1'b1),             .B_DOUT_EN (1'b1), 
        .A_DOUT_ARST_N (1'b1),         .B_DOUT_ARST_N (1'b1), 
        .A_DOUT_SRST_N (1'b1),         .B_DOUT_SRST_N (1'b1), 
        .A_DOUT_LAT (1'b1),            .B_DOUT_LAT (1'b1),
        .A_WIDTH (width40),             .B_WIDTH (width40), 
        .A_WMODE (1'b0),               .B_WMODE (1'b0),
        .A_EN (1'b1),                  .B_EN (1'b1),
        .BUSY (lsram_512_BUSY_40),
        .SII_LOCK (1'b0)
    );

    RAM1K18 block39 (
        .A_DOUT (readData39),           .B_DOUT (),
        .A_CLK (clk),                  .B_CLK (clk), 
        .A_ARST_N (resetn),            .B_ARST_N (resetn), 
        .A_BLK (3'b111),               .B_BLK (3'b111), 
        .A_DIN (writeData39),           .B_DIN (writeData39), 
        .A_ADDR (writeAddr39),          .B_ADDR (writeAddr39), 
        .A_WEN (wen_a39),               .B_WEN (wen_b39),
        .A_DOUT_CLK (1'b1),            .B_DOUT_CLK (1'b1), 
        .A_DOUT_EN (1'b1),             .B_DOUT_EN (1'b1), 
        .A_DOUT_ARST_N (1'b1),         .B_DOUT_ARST_N (1'b1), 
        .A_DOUT_SRST_N (1'b1),         .B_DOUT_SRST_N (1'b1), 
        .A_DOUT_LAT (1'b1),            .B_DOUT_LAT (1'b1),
        .A_WIDTH (width39),             .B_WIDTH (width39), 
        .A_WMODE (1'b0),               .B_WMODE (1'b0),
        .A_EN (1'b1),                  .B_EN (1'b1),
        .BUSY (lsram_512_BUSY_39),
        .SII_LOCK (1'b0)
    );

    RAM1K18 block38 (
        .A_DOUT (readData38),           .B_DOUT (),
        .A_CLK (clk),                  .B_CLK (clk), 
        .A_ARST_N (resetn),            .B_ARST_N (resetn), 
        .A_BLK (3'b111),               .B_BLK (3'b111), 
        .A_DIN (writeData38),           .B_DIN (writeData38), 
        .A_ADDR (writeAddr38),          .B_ADDR (writeAddr38), 
        .A_WEN (wen_a38),               .B_WEN (wen_b38),
        .A_DOUT_CLK (1'b1),            .B_DOUT_CLK (1'b1), 
        .A_DOUT_EN (1'b1),             .B_DOUT_EN (1'b1), 
        .A_DOUT_ARST_N (1'b1),         .B_DOUT_ARST_N (1'b1), 
        .A_DOUT_SRST_N (1'b1),         .B_DOUT_SRST_N (1'b1), 
        .A_DOUT_LAT (1'b1),            .B_DOUT_LAT (1'b1),
        .A_WIDTH (width38),             .B_WIDTH (width38), 
        .A_WMODE (1'b0),               .B_WMODE (1'b0),
        .A_EN (1'b1),                  .B_EN (1'b1),
        .BUSY (lsram_512_BUSY_38),
        .SII_LOCK (1'b0)
    );

    RAM1K18 block37 (
        .A_DOUT (readData37),           .B_DOUT (),
        .A_CLK (clk),                  .B_CLK (clk), 
        .A_ARST_N (resetn),            .B_ARST_N (resetn), 
        .A_BLK (3'b111),               .B_BLK (3'b111), 
        .A_DIN (writeData37),           .B_DIN (writeData37), 
        .A_ADDR (writeAddr37),          .B_ADDR (writeAddr37), 
        .A_WEN (wen_a37),               .B_WEN (wen_b37),
        .A_DOUT_CLK (1'b1),            .B_DOUT_CLK (1'b1), 
        .A_DOUT_EN (1'b1),             .B_DOUT_EN (1'b1), 
        .A_DOUT_ARST_N (1'b1),         .B_DOUT_ARST_N (1'b1), 
        .A_DOUT_SRST_N (1'b1),         .B_DOUT_SRST_N (1'b1), 
        .A_DOUT_LAT (1'b1),            .B_DOUT_LAT (1'b1),
        .A_WIDTH (width37),             .B_WIDTH (width37), 
        .A_WMODE (1'b0),               .B_WMODE (1'b0),
        .A_EN (1'b1),                  .B_EN (1'b1),
        .BUSY (lsram_512_BUSY_37),
        .SII_LOCK (1'b0)
    );

    RAM1K18 block36 (
        .A_DOUT (readData36),           .B_DOUT (),
        .A_CLK (clk),                  .B_CLK (clk), 
        .A_ARST_N (resetn),            .B_ARST_N (resetn), 
        .A_BLK (3'b111),               .B_BLK (3'b111), 
        .A_DIN (writeData36),           .B_DIN (writeData36), 
        .A_ADDR (writeAddr36),          .B_ADDR (writeAddr36), 
        .A_WEN (wen_a36),               .B_WEN (wen_b36),
        .A_DOUT_CLK (1'b1),            .B_DOUT_CLK (1'b1), 
        .A_DOUT_EN (1'b1),             .B_DOUT_EN (1'b1), 
        .A_DOUT_ARST_N (1'b1),         .B_DOUT_ARST_N (1'b1), 
        .A_DOUT_SRST_N (1'b1),         .B_DOUT_SRST_N (1'b1), 
        .A_DOUT_LAT (1'b1),            .B_DOUT_LAT (1'b1),
        .A_WIDTH (width36),             .B_WIDTH (width36), 
        .A_WMODE (1'b0),               .B_WMODE (1'b0),
        .A_EN (1'b1),                  .B_EN (1'b1),
        .BUSY (lsram_512_BUSY_36),
        .SII_LOCK (1'b0)
    );

    RAM1K18 block35 (
        .A_DOUT (readData35),           .B_DOUT (),
        .A_CLK (clk),                  .B_CLK (clk), 
        .A_ARST_N (resetn),            .B_ARST_N (resetn), 
        .A_BLK (3'b111),               .B_BLK (3'b111), 
        .A_DIN (writeData35),           .B_DIN (writeData35), 
        .A_ADDR (writeAddr35),          .B_ADDR (writeAddr35), 
        .A_WEN (wen_a35),               .B_WEN (wen_b35),
        .A_DOUT_CLK (1'b1),            .B_DOUT_CLK (1'b1), 
        .A_DOUT_EN (1'b1),             .B_DOUT_EN (1'b1), 
        .A_DOUT_ARST_N (1'b1),         .B_DOUT_ARST_N (1'b1), 
        .A_DOUT_SRST_N (1'b1),         .B_DOUT_SRST_N (1'b1), 
        .A_DOUT_LAT (1'b1),            .B_DOUT_LAT (1'b1),
        .A_WIDTH (width35),             .B_WIDTH (width35), 
        .A_WMODE (1'b0),               .B_WMODE (1'b0),
        .A_EN (1'b1),                  .B_EN (1'b1),
        .BUSY (lsram_512_BUSY_35),
        .SII_LOCK (1'b0)
    );

    RAM1K18 block34 (
        .A_DOUT (readData34),           .B_DOUT (),
        .A_CLK (clk),                  .B_CLK (clk), 
        .A_ARST_N (resetn),            .B_ARST_N (resetn), 
        .A_BLK (3'b111),               .B_BLK (3'b111), 
        .A_DIN (writeData34),           .B_DIN (writeData34), 
        .A_ADDR (writeAddr34),          .B_ADDR (writeAddr34), 
        .A_WEN (wen_a34),               .B_WEN (wen_b34),
        .A_DOUT_CLK (1'b1),            .B_DOUT_CLK (1'b1), 
        .A_DOUT_EN (1'b1),             .B_DOUT_EN (1'b1), 
        .A_DOUT_ARST_N (1'b1),         .B_DOUT_ARST_N (1'b1), 
        .A_DOUT_SRST_N (1'b1),         .B_DOUT_SRST_N (1'b1), 
        .A_DOUT_LAT (1'b1),            .B_DOUT_LAT (1'b1),
        .A_WIDTH (width34),             .B_WIDTH (width34), 
        .A_WMODE (1'b0),               .B_WMODE (1'b0),
        .A_EN (1'b1),                  .B_EN (1'b1),
        .BUSY (lsram_512_BUSY_34),
        .SII_LOCK (1'b0)
    );

    RAM1K18 block33 (
        .A_DOUT (readData33),           .B_DOUT (),
        .A_CLK (clk),                  .B_CLK (clk), 
        .A_ARST_N (resetn),            .B_ARST_N (resetn), 
        .A_BLK (3'b111),               .B_BLK (3'b111), 
        .A_DIN (writeData33),           .B_DIN (writeData33), 
        .A_ADDR (writeAddr33),          .B_ADDR (writeAddr33), 
        .A_WEN (wen_a33),               .B_WEN (wen_b33),
        .A_DOUT_CLK (1'b1),            .B_DOUT_CLK (1'b1), 
        .A_DOUT_EN (1'b1),             .B_DOUT_EN (1'b1), 
        .A_DOUT_ARST_N (1'b1),         .B_DOUT_ARST_N (1'b1), 
        .A_DOUT_SRST_N (1'b1),         .B_DOUT_SRST_N (1'b1), 
        .A_DOUT_LAT (1'b1),            .B_DOUT_LAT (1'b1),
        .A_WIDTH (width33),             .B_WIDTH (width33), 
        .A_WMODE (1'b0),               .B_WMODE (1'b0),
        .A_EN (1'b1),                  .B_EN (1'b1),
        .BUSY (lsram_512_BUSY_33),
        .SII_LOCK (1'b0)
    );

    RAM1K18 block32 (
        .A_DOUT (readData32),           .B_DOUT (),
        .A_CLK (clk),                  .B_CLK (clk), 
        .A_ARST_N (resetn),            .B_ARST_N (resetn), 
        .A_BLK (3'b111),               .B_BLK (3'b111), 
        .A_DIN (writeData32),           .B_DIN (writeData32), 
        .A_ADDR (writeAddr32),          .B_ADDR (writeAddr32), 
        .A_WEN (wen_a32),               .B_WEN (wen_b32),
        .A_DOUT_CLK (1'b1),            .B_DOUT_CLK (1'b1), 
        .A_DOUT_EN (1'b1),             .B_DOUT_EN (1'b1), 
        .A_DOUT_ARST_N (1'b1),         .B_DOUT_ARST_N (1'b1), 
        .A_DOUT_SRST_N (1'b1),         .B_DOUT_SRST_N (1'b1), 
        .A_DOUT_LAT (1'b1),            .B_DOUT_LAT (1'b1),
        .A_WIDTH (width32),             .B_WIDTH (width32), 
        .A_WMODE (1'b0),               .B_WMODE (1'b0),
        .A_EN (1'b1),                  .B_EN (1'b1),
        .BUSY (lsram_512_BUSY_32),
        .SII_LOCK (1'b0)
    );

    RAM1K18 block31 (
        .A_DOUT (readData31),           .B_DOUT (),
        .A_CLK (clk),                  .B_CLK (clk), 
        .A_ARST_N (resetn),            .B_ARST_N (resetn), 
        .A_BLK (3'b111),               .B_BLK (3'b111), 
        .A_DIN (writeData31),           .B_DIN (writeData31), 
        .A_ADDR (writeAddr31),          .B_ADDR (writeAddr31), 
        .A_WEN (wen_a31),               .B_WEN (wen_b31),
        .A_DOUT_CLK (1'b1),            .B_DOUT_CLK (1'b1), 
        .A_DOUT_EN (1'b1),             .B_DOUT_EN (1'b1), 
        .A_DOUT_ARST_N (1'b1),         .B_DOUT_ARST_N (1'b1), 
        .A_DOUT_SRST_N (1'b1),         .B_DOUT_SRST_N (1'b1), 
        .A_DOUT_LAT (1'b1),            .B_DOUT_LAT (1'b1),
        .A_WIDTH (width31),             .B_WIDTH (width31), 
        .A_WMODE (1'b0),               .B_WMODE (1'b0),
        .A_EN (1'b1),                  .B_EN (1'b1),
        .BUSY (lsram_512_BUSY_31),
        .SII_LOCK (1'b0)
    );

    RAM1K18 block30 (
        .A_DOUT (readData30),           .B_DOUT (),
        .A_CLK (clk),                  .B_CLK (clk), 
        .A_ARST_N (resetn),            .B_ARST_N (resetn), 
        .A_BLK (3'b111),               .B_BLK (3'b111), 
        .A_DIN (writeData30),           .B_DIN (writeData30), 
        .A_ADDR (writeAddr30),          .B_ADDR (writeAddr30), 
        .A_WEN (wen_a30),               .B_WEN (wen_b30),
        .A_DOUT_CLK (1'b1),            .B_DOUT_CLK (1'b1), 
        .A_DOUT_EN (1'b1),             .B_DOUT_EN (1'b1), 
        .A_DOUT_ARST_N (1'b1),         .B_DOUT_ARST_N (1'b1), 
        .A_DOUT_SRST_N (1'b1),         .B_DOUT_SRST_N (1'b1), 
        .A_DOUT_LAT (1'b1),            .B_DOUT_LAT (1'b1),
        .A_WIDTH (width30),             .B_WIDTH (width30), 
        .A_WMODE (1'b0),               .B_WMODE (1'b0),
        .A_EN (1'b1),                  .B_EN (1'b1),
        .BUSY (lsram_512_BUSY_30),
        .SII_LOCK (1'b0)
    );

    RAM1K18 block29 (
        .A_DOUT (readData29),           .B_DOUT (),
        .A_CLK (clk),                  .B_CLK (clk), 
        .A_ARST_N (resetn),            .B_ARST_N (resetn), 
        .A_BLK (3'b111),               .B_BLK (3'b111), 
        .A_DIN (writeData29),           .B_DIN (writeData29), 
        .A_ADDR (writeAddr29),          .B_ADDR (writeAddr29), 
        .A_WEN (wen_a29),               .B_WEN (wen_b29),
        .A_DOUT_CLK (1'b1),            .B_DOUT_CLK (1'b1), 
        .A_DOUT_EN (1'b1),             .B_DOUT_EN (1'b1), 
        .A_DOUT_ARST_N (1'b1),         .B_DOUT_ARST_N (1'b1), 
        .A_DOUT_SRST_N (1'b1),         .B_DOUT_SRST_N (1'b1), 
        .A_DOUT_LAT (1'b1),            .B_DOUT_LAT (1'b1),
        .A_WIDTH (width29),             .B_WIDTH (width29), 
        .A_WMODE (1'b0),               .B_WMODE (1'b0),
        .A_EN (1'b1),                  .B_EN (1'b1),
        .BUSY (lsram_512_BUSY_29),
        .SII_LOCK (1'b0)
    );

    RAM1K18 block28 (
        .A_DOUT (readData28),           .B_DOUT (),
        .A_CLK (clk),                  .B_CLK (clk), 
        .A_ARST_N (resetn),            .B_ARST_N (resetn), 
        .A_BLK (3'b111),               .B_BLK (3'b111), 
        .A_DIN (writeData28),           .B_DIN (writeData28), 
        .A_ADDR (writeAddr28),          .B_ADDR (writeAddr28), 
        .A_WEN (wen_a28),               .B_WEN (wen_b28),
        .A_DOUT_CLK (1'b1),            .B_DOUT_CLK (1'b1), 
        .A_DOUT_EN (1'b1),             .B_DOUT_EN (1'b1), 
        .A_DOUT_ARST_N (1'b1),         .B_DOUT_ARST_N (1'b1), 
        .A_DOUT_SRST_N (1'b1),         .B_DOUT_SRST_N (1'b1), 
        .A_DOUT_LAT (1'b1),            .B_DOUT_LAT (1'b1),
        .A_WIDTH (width28),             .B_WIDTH (width28), 
        .A_WMODE (1'b0),               .B_WMODE (1'b0),
        .A_EN (1'b1),                  .B_EN (1'b1),
        .BUSY (lsram_512_BUSY_28),
        .SII_LOCK (1'b0)
    );

    RAM1K18 block27 (
        .A_DOUT (readData27),           .B_DOUT (),
        .A_CLK (clk),                  .B_CLK (clk), 
        .A_ARST_N (resetn),            .B_ARST_N (resetn), 
        .A_BLK (3'b111),               .B_BLK (3'b111), 
        .A_DIN (writeData27),           .B_DIN (writeData27), 
        .A_ADDR (writeAddr27),          .B_ADDR (writeAddr27), 
        .A_WEN (wen_a27),               .B_WEN (wen_b27),
        .A_DOUT_CLK (1'b1),            .B_DOUT_CLK (1'b1), 
        .A_DOUT_EN (1'b1),             .B_DOUT_EN (1'b1), 
        .A_DOUT_ARST_N (1'b1),         .B_DOUT_ARST_N (1'b1), 
        .A_DOUT_SRST_N (1'b1),         .B_DOUT_SRST_N (1'b1), 
        .A_DOUT_LAT (1'b1),            .B_DOUT_LAT (1'b1),
        .A_WIDTH (width27),             .B_WIDTH (width27), 
        .A_WMODE (1'b0),               .B_WMODE (1'b0),
        .A_EN (1'b1),                  .B_EN (1'b1),
        .BUSY (lsram_512_BUSY_27),
        .SII_LOCK (1'b0)
    );

    RAM1K18 block26 (
        .A_DOUT (readData26),           .B_DOUT (),
        .A_CLK (clk),                  .B_CLK (clk), 
        .A_ARST_N (resetn),            .B_ARST_N (resetn), 
        .A_BLK (3'b111),               .B_BLK (3'b111), 
        .A_DIN (writeData26),           .B_DIN (writeData26), 
        .A_ADDR (writeAddr26),          .B_ADDR (writeAddr26), 
        .A_WEN (wen_a26),               .B_WEN (wen_b26),
        .A_DOUT_CLK (1'b1),            .B_DOUT_CLK (1'b1), 
        .A_DOUT_EN (1'b1),             .B_DOUT_EN (1'b1), 
        .A_DOUT_ARST_N (1'b1),         .B_DOUT_ARST_N (1'b1), 
        .A_DOUT_SRST_N (1'b1),         .B_DOUT_SRST_N (1'b1), 
        .A_DOUT_LAT (1'b1),            .B_DOUT_LAT (1'b1),
        .A_WIDTH (width26),             .B_WIDTH (width26), 
        .A_WMODE (1'b0),               .B_WMODE (1'b0),
        .A_EN (1'b1),                  .B_EN (1'b1),
        .BUSY (lsram_512_BUSY_26),
        .SII_LOCK (1'b0)
    );

    RAM1K18 block25 (
        .A_DOUT (readData25),           .B_DOUT (),
        .A_CLK (clk),                  .B_CLK (clk), 
        .A_ARST_N (resetn),            .B_ARST_N (resetn), 
        .A_BLK (3'b111),               .B_BLK (3'b111), 
        .A_DIN (writeData25),           .B_DIN (writeData25), 
        .A_ADDR (writeAddr25),          .B_ADDR (writeAddr25), 
        .A_WEN (wen_a25),               .B_WEN (wen_b25),
        .A_DOUT_CLK (1'b1),            .B_DOUT_CLK (1'b1), 
        .A_DOUT_EN (1'b1),             .B_DOUT_EN (1'b1), 
        .A_DOUT_ARST_N (1'b1),         .B_DOUT_ARST_N (1'b1), 
        .A_DOUT_SRST_N (1'b1),         .B_DOUT_SRST_N (1'b1), 
        .A_DOUT_LAT (1'b1),            .B_DOUT_LAT (1'b1),
        .A_WIDTH (width25),             .B_WIDTH (width25), 
        .A_WMODE (1'b0),               .B_WMODE (1'b0),
        .A_EN (1'b1),                  .B_EN (1'b1),
        .BUSY (lsram_512_BUSY_25),
        .SII_LOCK (1'b0)
    );

    RAM1K18 block24 (
        .A_DOUT (readData24),           .B_DOUT (),
        .A_CLK (clk),                  .B_CLK (clk), 
        .A_ARST_N (resetn),            .B_ARST_N (resetn), 
        .A_BLK (3'b111),               .B_BLK (3'b111), 
        .A_DIN (writeData24),           .B_DIN (writeData24), 
        .A_ADDR (writeAddr24),          .B_ADDR (writeAddr24), 
        .A_WEN (wen_a24),               .B_WEN (wen_b24),
        .A_DOUT_CLK (1'b1),            .B_DOUT_CLK (1'b1), 
        .A_DOUT_EN (1'b1),             .B_DOUT_EN (1'b1), 
        .A_DOUT_ARST_N (1'b1),         .B_DOUT_ARST_N (1'b1), 
        .A_DOUT_SRST_N (1'b1),         .B_DOUT_SRST_N (1'b1), 
        .A_DOUT_LAT (1'b1),            .B_DOUT_LAT (1'b1),
        .A_WIDTH (width24),             .B_WIDTH (width24), 
        .A_WMODE (1'b0),               .B_WMODE (1'b0),
        .A_EN (1'b1),                  .B_EN (1'b1),
        .BUSY (lsram_512_BUSY_24),
        .SII_LOCK (1'b0)
    );

    RAM1K18 block23 (
        .A_DOUT (readData23),           .B_DOUT (),
        .A_CLK (clk),                  .B_CLK (clk), 
        .A_ARST_N (resetn),            .B_ARST_N (resetn), 
        .A_BLK (3'b111),               .B_BLK (3'b111), 
        .A_DIN (writeData23),           .B_DIN (writeData23), 
        .A_ADDR (writeAddr23),          .B_ADDR (writeAddr23), 
        .A_WEN (wen_a23),               .B_WEN (wen_b23),
        .A_DOUT_CLK (1'b1),            .B_DOUT_CLK (1'b1), 
        .A_DOUT_EN (1'b1),             .B_DOUT_EN (1'b1), 
        .A_DOUT_ARST_N (1'b1),         .B_DOUT_ARST_N (1'b1), 
        .A_DOUT_SRST_N (1'b1),         .B_DOUT_SRST_N (1'b1), 
        .A_DOUT_LAT (1'b1),            .B_DOUT_LAT (1'b1),
        .A_WIDTH (width23),             .B_WIDTH (width23), 
        .A_WMODE (1'b0),               .B_WMODE (1'b0),
        .A_EN (1'b1),                  .B_EN (1'b1),
        .BUSY (lsram_512_BUSY_23),
        .SII_LOCK (1'b0)
    );

    RAM1K18 block22 (
        .A_DOUT (readData22),           .B_DOUT (),
        .A_CLK (clk),                  .B_CLK (clk), 
        .A_ARST_N (resetn),            .B_ARST_N (resetn), 
        .A_BLK (3'b111),               .B_BLK (3'b111), 
        .A_DIN (writeData22),           .B_DIN (writeData22), 
        .A_ADDR (writeAddr22),          .B_ADDR (writeAddr22), 
        .A_WEN (wen_a22),               .B_WEN (wen_b22),
        .A_DOUT_CLK (1'b1),            .B_DOUT_CLK (1'b1), 
        .A_DOUT_EN (1'b1),             .B_DOUT_EN (1'b1), 
        .A_DOUT_ARST_N (1'b1),         .B_DOUT_ARST_N (1'b1), 
        .A_DOUT_SRST_N (1'b1),         .B_DOUT_SRST_N (1'b1), 
        .A_DOUT_LAT (1'b1),            .B_DOUT_LAT (1'b1),
        .A_WIDTH (width22),             .B_WIDTH (width22), 
        .A_WMODE (1'b0),               .B_WMODE (1'b0),
        .A_EN (1'b1),                  .B_EN (1'b1),
        .BUSY (lsram_512_BUSY_22),
        .SII_LOCK (1'b0)
    );

    RAM1K18 block21 (
        .A_DOUT (readData21),           .B_DOUT (),
        .A_CLK (clk),                  .B_CLK (clk), 
        .A_ARST_N (resetn),            .B_ARST_N (resetn), 
        .A_BLK (3'b111),               .B_BLK (3'b111), 
        .A_DIN (writeData21),           .B_DIN (writeData21), 
        .A_ADDR (writeAddr21),          .B_ADDR (writeAddr21), 
        .A_WEN (wen_a21),               .B_WEN (wen_b21),
        .A_DOUT_CLK (1'b1),            .B_DOUT_CLK (1'b1), 
        .A_DOUT_EN (1'b1),             .B_DOUT_EN (1'b1), 
        .A_DOUT_ARST_N (1'b1),         .B_DOUT_ARST_N (1'b1), 
        .A_DOUT_SRST_N (1'b1),         .B_DOUT_SRST_N (1'b1), 
        .A_DOUT_LAT (1'b1),            .B_DOUT_LAT (1'b1),
        .A_WIDTH (width21),             .B_WIDTH (width21), 
        .A_WMODE (1'b0),               .B_WMODE (1'b0),
        .A_EN (1'b1),                  .B_EN (1'b1),
        .BUSY (lsram_512_BUSY_21),
        .SII_LOCK (1'b0)
    );

    RAM1K18 block20 (
        .A_DOUT (readData20),           .B_DOUT (),
        .A_CLK (clk),                  .B_CLK (clk), 
        .A_ARST_N (resetn),            .B_ARST_N (resetn), 
        .A_BLK (3'b111),               .B_BLK (3'b111), 
        .A_DIN (writeData20),           .B_DIN (writeData20), 
        .A_ADDR (writeAddr20),          .B_ADDR (writeAddr20), 
        .A_WEN (wen_a20),               .B_WEN (wen_b20),
        .A_DOUT_CLK (1'b1),            .B_DOUT_CLK (1'b1), 
        .A_DOUT_EN (1'b1),             .B_DOUT_EN (1'b1), 
        .A_DOUT_ARST_N (1'b1),         .B_DOUT_ARST_N (1'b1), 
        .A_DOUT_SRST_N (1'b1),         .B_DOUT_SRST_N (1'b1), 
        .A_DOUT_LAT (1'b1),            .B_DOUT_LAT (1'b1),
        .A_WIDTH (width20),             .B_WIDTH (width20), 
        .A_WMODE (1'b0),               .B_WMODE (1'b0),
        .A_EN (1'b1),                  .B_EN (1'b1),
        .BUSY (lsram_512_BUSY_20),
        .SII_LOCK (1'b0)
    );

    RAM1K18 block19 (
        .A_DOUT (readData19),           .B_DOUT (),
        .A_CLK (clk),                  .B_CLK (clk), 
        .A_ARST_N (resetn),            .B_ARST_N (resetn), 
        .A_BLK (3'b111),               .B_BLK (3'b111), 
        .A_DIN (writeData19),           .B_DIN (writeData19), 
        .A_ADDR (writeAddr19),          .B_ADDR (writeAddr19), 
        .A_WEN (wen_a19),               .B_WEN (wen_b19),
        .A_DOUT_CLK (1'b1),            .B_DOUT_CLK (1'b1), 
        .A_DOUT_EN (1'b1),             .B_DOUT_EN (1'b1), 
        .A_DOUT_ARST_N (1'b1),         .B_DOUT_ARST_N (1'b1), 
        .A_DOUT_SRST_N (1'b1),         .B_DOUT_SRST_N (1'b1), 
        .A_DOUT_LAT (1'b1),            .B_DOUT_LAT (1'b1),
        .A_WIDTH (width19),             .B_WIDTH (width19), 
        .A_WMODE (1'b0),               .B_WMODE (1'b0),
        .A_EN (1'b1),                  .B_EN (1'b1),
        .BUSY (lsram_512_BUSY_19),
        .SII_LOCK (1'b0)
    );

    RAM1K18 block18 (
        .A_DOUT (readData18),           .B_DOUT (),
        .A_CLK (clk),                  .B_CLK (clk), 
        .A_ARST_N (resetn),            .B_ARST_N (resetn), 
        .A_BLK (3'b111),               .B_BLK (3'b111), 
        .A_DIN (writeData18),           .B_DIN (writeData18), 
        .A_ADDR (writeAddr18),          .B_ADDR (writeAddr18), 
        .A_WEN (wen_a18),               .B_WEN (wen_b18),
        .A_DOUT_CLK (1'b1),            .B_DOUT_CLK (1'b1), 
        .A_DOUT_EN (1'b1),             .B_DOUT_EN (1'b1), 
        .A_DOUT_ARST_N (1'b1),         .B_DOUT_ARST_N (1'b1), 
        .A_DOUT_SRST_N (1'b1),         .B_DOUT_SRST_N (1'b1), 
        .A_DOUT_LAT (1'b1),            .B_DOUT_LAT (1'b1),
        .A_WIDTH (width18),             .B_WIDTH (width18), 
        .A_WMODE (1'b0),               .B_WMODE (1'b0),
        .A_EN (1'b1),                  .B_EN (1'b1),
        .BUSY (lsram_512_BUSY_18),
        .SII_LOCK (1'b0)
    );

    RAM1K18 block17 (
        .A_DOUT (readData17),           .B_DOUT (),
        .A_CLK (clk),                  .B_CLK (clk), 
        .A_ARST_N (resetn),            .B_ARST_N (resetn), 
        .A_BLK (3'b111),               .B_BLK (3'b111), 
        .A_DIN (writeData17),           .B_DIN (writeData17), 
        .A_ADDR (writeAddr17),          .B_ADDR (writeAddr17), 
        .A_WEN (wen_a17),               .B_WEN (wen_b17),
        .A_DOUT_CLK (1'b1),            .B_DOUT_CLK (1'b1), 
        .A_DOUT_EN (1'b1),             .B_DOUT_EN (1'b1), 
        .A_DOUT_ARST_N (1'b1),         .B_DOUT_ARST_N (1'b1), 
        .A_DOUT_SRST_N (1'b1),         .B_DOUT_SRST_N (1'b1), 
        .A_DOUT_LAT (1'b1),            .B_DOUT_LAT (1'b1),
        .A_WIDTH (width17),             .B_WIDTH (width17), 
        .A_WMODE (1'b0),               .B_WMODE (1'b0),
        .A_EN (1'b1),                  .B_EN (1'b1),
        .BUSY (lsram_512_BUSY_17),
        .SII_LOCK (1'b0)
    );

    RAM1K18 block16 (
        .A_DOUT (readData16),           .B_DOUT (),
        .A_CLK (clk),                  .B_CLK (clk), 
        .A_ARST_N (resetn),            .B_ARST_N (resetn), 
        .A_BLK (3'b111),               .B_BLK (3'b111), 
        .A_DIN (writeData16),           .B_DIN (writeData16), 
        .A_ADDR (writeAddr16),          .B_ADDR (writeAddr16), 
        .A_WEN (wen_a16),               .B_WEN (wen_b16),
        .A_DOUT_CLK (1'b1),            .B_DOUT_CLK (1'b1), 
        .A_DOUT_EN (1'b1),             .B_DOUT_EN (1'b1), 
        .A_DOUT_ARST_N (1'b1),         .B_DOUT_ARST_N (1'b1), 
        .A_DOUT_SRST_N (1'b1),         .B_DOUT_SRST_N (1'b1), 
        .A_DOUT_LAT (1'b1),            .B_DOUT_LAT (1'b1),
        .A_WIDTH (width16),             .B_WIDTH (width16), 
        .A_WMODE (1'b0),               .B_WMODE (1'b0),
        .A_EN (1'b1),                  .B_EN (1'b1),
        .BUSY (lsram_512_BUSY_16),
        .SII_LOCK (1'b0)
    );

    RAM1K18 block15 (
        .A_DOUT (readData15),           .B_DOUT (),
        .A_CLK (clk),                  .B_CLK (clk), 
        .A_ARST_N (resetn),            .B_ARST_N (resetn), 
        .A_BLK (3'b111),               .B_BLK (3'b111), 
        .A_DIN (writeData15),           .B_DIN (writeData15), 
        .A_ADDR (writeAddr15),          .B_ADDR (writeAddr15), 
        .A_WEN (wen_a15),               .B_WEN (wen_b15),
        .A_DOUT_CLK (1'b1),            .B_DOUT_CLK (1'b1), 
        .A_DOUT_EN (1'b1),             .B_DOUT_EN (1'b1), 
        .A_DOUT_ARST_N (1'b1),         .B_DOUT_ARST_N (1'b1), 
        .A_DOUT_SRST_N (1'b1),         .B_DOUT_SRST_N (1'b1), 
        .A_DOUT_LAT (1'b1),            .B_DOUT_LAT (1'b1),
        .A_WIDTH (width15),             .B_WIDTH (width15), 
        .A_WMODE (1'b0),               .B_WMODE (1'b0),
        .A_EN (1'b1),                  .B_EN (1'b1),
        .BUSY (lsram_512_BUSY_15),
        .SII_LOCK (1'b0)
    );

    RAM1K18 block14 (
        .A_DOUT (readData14),           .B_DOUT (),
        .A_CLK (clk),                  .B_CLK (clk), 
        .A_ARST_N (resetn),            .B_ARST_N (resetn), 
        .A_BLK (3'b111),               .B_BLK (3'b111), 
        .A_DIN (writeData14),           .B_DIN (writeData14), 
        .A_ADDR (writeAddr14),          .B_ADDR (writeAddr14), 
        .A_WEN (wen_a14),               .B_WEN (wen_b14),
        .A_DOUT_CLK (1'b1),            .B_DOUT_CLK (1'b1), 
        .A_DOUT_EN (1'b1),             .B_DOUT_EN (1'b1), 
        .A_DOUT_ARST_N (1'b1),         .B_DOUT_ARST_N (1'b1), 
        .A_DOUT_SRST_N (1'b1),         .B_DOUT_SRST_N (1'b1), 
        .A_DOUT_LAT (1'b1),            .B_DOUT_LAT (1'b1),
        .A_WIDTH (width14),             .B_WIDTH (width14), 
        .A_WMODE (1'b0),               .B_WMODE (1'b0),
        .A_EN (1'b1),                  .B_EN (1'b1),
        .BUSY (lsram_512_BUSY_14),
        .SII_LOCK (1'b0)
    );

    RAM1K18 block13 (
        .A_DOUT (readData13),           .B_DOUT (),
        .A_CLK (clk),                  .B_CLK (clk), 
        .A_ARST_N (resetn),            .B_ARST_N (resetn), 
        .A_BLK (3'b111),               .B_BLK (3'b111), 
        .A_DIN (writeData13),           .B_DIN (writeData13), 
        .A_ADDR (writeAddr13),          .B_ADDR (writeAddr13), 
        .A_WEN (wen_a13),               .B_WEN (wen_b13),
        .A_DOUT_CLK (1'b1),            .B_DOUT_CLK (1'b1), 
        .A_DOUT_EN (1'b1),             .B_DOUT_EN (1'b1), 
        .A_DOUT_ARST_N (1'b1),         .B_DOUT_ARST_N (1'b1), 
        .A_DOUT_SRST_N (1'b1),         .B_DOUT_SRST_N (1'b1), 
        .A_DOUT_LAT (1'b1),            .B_DOUT_LAT (1'b1),
        .A_WIDTH (width13),             .B_WIDTH (width13), 
        .A_WMODE (1'b0),               .B_WMODE (1'b0),
        .A_EN (1'b1),                  .B_EN (1'b1),
        .BUSY (lsram_512_BUSY_13),
        .SII_LOCK (1'b0)
    );

    RAM1K18 block12 (
        .A_DOUT (readData12),           .B_DOUT (),
        .A_CLK (clk),                  .B_CLK (clk), 
        .A_ARST_N (resetn),            .B_ARST_N (resetn), 
        .A_BLK (3'b111),               .B_BLK (3'b111), 
        .A_DIN (writeData12),           .B_DIN (writeData12), 
        .A_ADDR (writeAddr12),          .B_ADDR (writeAddr12), 
        .A_WEN (wen_a12),               .B_WEN (wen_b12),
        .A_DOUT_CLK (1'b1),            .B_DOUT_CLK (1'b1), 
        .A_DOUT_EN (1'b1),             .B_DOUT_EN (1'b1), 
        .A_DOUT_ARST_N (1'b1),         .B_DOUT_ARST_N (1'b1), 
        .A_DOUT_SRST_N (1'b1),         .B_DOUT_SRST_N (1'b1), 
        .A_DOUT_LAT (1'b1),            .B_DOUT_LAT (1'b1),
        .A_WIDTH (width12),             .B_WIDTH (width12), 
        .A_WMODE (1'b0),               .B_WMODE (1'b0),
        .A_EN (1'b1),                  .B_EN (1'b1),
        .BUSY (lsram_512_BUSY_12),
        .SII_LOCK (1'b0)
    );

    RAM1K18 block11 (
        .A_DOUT (readData11),           .B_DOUT (),
        .A_CLK (clk),                  .B_CLK (clk), 
        .A_ARST_N (resetn),            .B_ARST_N (resetn), 
        .A_BLK (3'b111),               .B_BLK (3'b111), 
        .A_DIN (writeData11),           .B_DIN (writeData11), 
        .A_ADDR (writeAddr11),          .B_ADDR (writeAddr11), 
        .A_WEN (wen_a11),               .B_WEN (wen_b11),
        .A_DOUT_CLK (1'b1),            .B_DOUT_CLK (1'b1), 
        .A_DOUT_EN (1'b1),             .B_DOUT_EN (1'b1), 
        .A_DOUT_ARST_N (1'b1),         .B_DOUT_ARST_N (1'b1), 
        .A_DOUT_SRST_N (1'b1),         .B_DOUT_SRST_N (1'b1), 
        .A_DOUT_LAT (1'b1),            .B_DOUT_LAT (1'b1),
        .A_WIDTH (width11),             .B_WIDTH (width11), 
        .A_WMODE (1'b0),               .B_WMODE (1'b0),
        .A_EN (1'b1),                  .B_EN (1'b1),
        .BUSY (lsram_512_BUSY_11),
        .SII_LOCK (1'b0)
    );

    RAM1K18 block10 (
        .A_DOUT (readData10),           .B_DOUT (),
        .A_CLK (clk),                  .B_CLK (clk), 
        .A_ARST_N (resetn),            .B_ARST_N (resetn), 
        .A_BLK (3'b111),               .B_BLK (3'b111), 
        .A_DIN (writeData10),           .B_DIN (writeData10), 
        .A_ADDR (writeAddr10),          .B_ADDR (writeAddr10), 
        .A_WEN (wen_a10),               .B_WEN (wen_b10),
        .A_DOUT_CLK (1'b1),            .B_DOUT_CLK (1'b1), 
        .A_DOUT_EN (1'b1),             .B_DOUT_EN (1'b1), 
        .A_DOUT_ARST_N (1'b1),         .B_DOUT_ARST_N (1'b1), 
        .A_DOUT_SRST_N (1'b1),         .B_DOUT_SRST_N (1'b1), 
        .A_DOUT_LAT (1'b1),            .B_DOUT_LAT (1'b1),
        .A_WIDTH (width10),             .B_WIDTH (width10), 
        .A_WMODE (1'b0),               .B_WMODE (1'b0),
        .A_EN (1'b1),                  .B_EN (1'b1),
        .BUSY (lsram_512_BUSY_10),
        .SII_LOCK (1'b0)
    );

    RAM1K18 block9 (
        .A_DOUT (readData9),           .B_DOUT (),
        .A_CLK (clk),                  .B_CLK (clk), 
        .A_ARST_N (resetn),            .B_ARST_N (resetn), 
        .A_BLK (3'b111),               .B_BLK (3'b111), 
        .A_DIN (writeData9),           .B_DIN (writeData9), 
        .A_ADDR (writeAddr9),          .B_ADDR (writeAddr9), 
        .A_WEN (wen_a9),               .B_WEN (wen_b9),
        .A_DOUT_CLK (1'b1),            .B_DOUT_CLK (1'b1), 
        .A_DOUT_EN (1'b1),             .B_DOUT_EN (1'b1), 
        .A_DOUT_ARST_N (1'b1),         .B_DOUT_ARST_N (1'b1), 
        .A_DOUT_SRST_N (1'b1),         .B_DOUT_SRST_N (1'b1), 
        .A_DOUT_LAT (1'b1),            .B_DOUT_LAT (1'b1),
        .A_WIDTH (width9),             .B_WIDTH (width9), 
        .A_WMODE (1'b0),               .B_WMODE (1'b0),
        .A_EN (1'b1),                  .B_EN (1'b1),
        .BUSY (lsram_512_BUSY_9),
        .SII_LOCK (1'b0)
    );

    RAM1K18 block8 (
        .A_DOUT (readData8),           .B_DOUT (),
        .A_CLK (clk),                  .B_CLK (clk), 
        .A_ARST_N (resetn),            .B_ARST_N (resetn), 
        .A_BLK (3'b111),               .B_BLK (3'b111), 
        .A_DIN (writeData8),           .B_DIN (writeData8), 
        .A_ADDR (writeAddr8),          .B_ADDR (writeAddr8), 
        .A_WEN (wen_a8),               .B_WEN (wen_b8),
        .A_DOUT_CLK (1'b1),            .B_DOUT_CLK (1'b1), 
        .A_DOUT_EN (1'b1),             .B_DOUT_EN (1'b1), 
        .A_DOUT_ARST_N (1'b1),         .B_DOUT_ARST_N (1'b1), 
        .A_DOUT_SRST_N (1'b1),         .B_DOUT_SRST_N (1'b1), 
        .A_DOUT_LAT (1'b1),            .B_DOUT_LAT (1'b1),
        .A_WIDTH (width8),             .B_WIDTH (width8), 
        .A_WMODE (1'b0),               .B_WMODE (1'b0),
        .A_EN (1'b1),                  .B_EN (1'b1),
        .BUSY (lsram_512_BUSY_8),
        .SII_LOCK (1'b0)
    );

    RAM1K18 block7 (
        .A_DOUT (readData7),           .B_DOUT (),
        .A_CLK (clk),                  .B_CLK (clk), 
        .A_ARST_N (resetn),            .B_ARST_N (resetn), 
        .A_BLK (3'b111),               .B_BLK (3'b111), 
        .A_DIN (writeData7),           .B_DIN (writeData7), 
        .A_ADDR (writeAddr7),          .B_ADDR (writeAddr7), 
        .A_WEN (wen_a7),               .B_WEN (wen_b7),
        .A_DOUT_CLK (1'b1),            .B_DOUT_CLK (1'b1), 
        .A_DOUT_EN (1'b1),             .B_DOUT_EN (1'b1), 
        .A_DOUT_ARST_N (1'b1),         .B_DOUT_ARST_N (1'b1), 
        .A_DOUT_SRST_N (1'b1),         .B_DOUT_SRST_N (1'b1), 
        .A_DOUT_LAT (1'b1),            .B_DOUT_LAT (1'b1),
        .A_WIDTH (width7),             .B_WIDTH (width7), 
        .A_WMODE (1'b0),               .B_WMODE (1'b0),
        .A_EN (1'b1),                  .B_EN (1'b1),
        .BUSY (lsram_512_BUSY_7),
        .SII_LOCK (1'b0)
    );

  RAM1K18 block6 (
        .A_DOUT (readData6),           .B_DOUT (),
        .A_CLK (clk),                  .B_CLK (clk), 
        .A_ARST_N (resetn),            .B_ARST_N (resetn), 
        .A_BLK (3'b111),               .B_BLK (3'b111), 
        .A_DIN (writeData6),           .B_DIN (writeData6), 
        .A_ADDR (writeAddr6),          .B_ADDR (writeAddr6), 
        .A_WEN (wen_a6),               .B_WEN (wen_b6),
        .A_DOUT_CLK (1'b1),            .B_DOUT_CLK (1'b1), 
        .A_DOUT_EN (1'b1),             .B_DOUT_EN (1'b1), 
        .A_DOUT_ARST_N (1'b1),         .B_DOUT_ARST_N (1'b1), 
        .A_DOUT_SRST_N (1'b1),         .B_DOUT_SRST_N (1'b1), 
        .A_DOUT_LAT (1'b1),            .B_DOUT_LAT (1'b1),
        .A_WIDTH (width6),             .B_WIDTH (width6), 
        .A_WMODE (1'b0),               .B_WMODE (1'b0),
        .A_EN (1'b1),                  .B_EN (1'b1),
        .BUSY (lsram_512_BUSY_6),
        .SII_LOCK (1'b0)
    );

    RAM1K18 block5 (
        .A_DOUT (readData5),           .B_DOUT (),
        .A_CLK (clk),                  .B_CLK (clk), 
        .A_ARST_N (resetn),            .B_ARST_N (resetn), 
        .A_BLK (3'b111),               .B_BLK (3'b111), 
        .A_DIN (writeData5),           .B_DIN (writeData5), 
        .A_ADDR (writeAddr5),          .B_ADDR (writeAddr5), 
        .A_WEN (wen_a5),               .B_WEN (wen_b5),
        .A_DOUT_CLK (1'b1),            .B_DOUT_CLK (1'b1), 
        .A_DOUT_EN (1'b1),             .B_DOUT_EN (1'b1), 
        .A_DOUT_ARST_N (1'b1),         .B_DOUT_ARST_N (1'b1), 
        .A_DOUT_SRST_N (1'b1),         .B_DOUT_SRST_N (1'b1), 
        .A_DOUT_LAT (1'b1),            .B_DOUT_LAT (1'b1),
        .A_WIDTH (width5),             .B_WIDTH (width5), 
        .A_WMODE (1'b0),               .B_WMODE (1'b0),
        .A_EN (1'b1),                  .B_EN (1'b1),
        .BUSY (lsram_512_BUSY_5),
        .SII_LOCK (1'b0)
    );

    RAM1K18 block4 (
        .A_DOUT (readData4),           .B_DOUT (),
        .A_CLK (clk),                  .B_CLK (clk), 
        .A_ARST_N (resetn),            .B_ARST_N (resetn), 
        .A_BLK (3'b111),               .B_BLK (3'b111), 
        .A_DIN (writeData4),           .B_DIN (writeData4), 
        .A_ADDR (writeAddr4),          .B_ADDR (writeAddr4), 
        .A_WEN (wen_a4),               .B_WEN (wen_b4),
        .A_DOUT_CLK (1'b1),            .B_DOUT_CLK (1'b1), 
        .A_DOUT_EN (1'b1),             .B_DOUT_EN (1'b1), 
        .A_DOUT_ARST_N (1'b1),         .B_DOUT_ARST_N (1'b1), 
        .A_DOUT_SRST_N (1'b1),         .B_DOUT_SRST_N (1'b1), 
        .A_DOUT_LAT (1'b1),            .B_DOUT_LAT (1'b1),
        .A_WIDTH (width4),             .B_WIDTH (width4), 
        .A_WMODE (1'b0),               .B_WMODE (1'b0),
        .A_EN (1'b1),                  .B_EN (1'b1),
        .BUSY (lsram_512_BUSY_4),
        .SII_LOCK (1'b0)
    );

    RAM1K18 block3 (
        .A_DOUT (readData3),           .B_DOUT (),
        .A_CLK (clk),                  .B_CLK (clk), 
        .A_ARST_N (resetn),            .B_ARST_N (resetn), 
        .A_BLK (3'b111),               .B_BLK (3'b111), 
        .A_DIN (writeData3),           .B_DIN (writeData3), 
        .A_ADDR (writeAddr3),          .B_ADDR (writeAddr3), 
        .A_WEN (wen_a3),               .B_WEN (wen_b3),
        .A_DOUT_CLK (1'b1),            .B_DOUT_CLK (1'b1), 
        .A_DOUT_EN (1'b1),             .B_DOUT_EN (1'b1), 
        .A_DOUT_ARST_N (1'b1),         .B_DOUT_ARST_N (1'b1), 
        .A_DOUT_SRST_N (1'b1),         .B_DOUT_SRST_N (1'b1), 
        .A_DOUT_LAT (1'b1),            .B_DOUT_LAT (1'b1),
        .A_WIDTH (width3),             .B_WIDTH (width3), 
        .A_WMODE (1'b0),               .B_WMODE (1'b0),
        .A_EN (1'b1),                  .B_EN (1'b1),
        .BUSY (lsram_512_BUSY_3),
        .SII_LOCK (1'b0)
    );

    RAM1K18 block2 (
        .A_DOUT (readData2),           .B_DOUT (),
        .A_CLK (clk),                  .B_CLK (clk), 
        .A_ARST_N (resetn),            .B_ARST_N (resetn), 
        .A_BLK (3'b111),               .B_BLK (3'b111), 
        .A_DIN (writeData2),           .B_DIN (writeData2), 
        .A_ADDR (writeAddr2),          .B_ADDR (writeAddr2), 
        .A_WEN (wen_a2),               .B_WEN (wen_b2),
        .A_DOUT_CLK (1'b1),            .B_DOUT_CLK (1'b1), 
        .A_DOUT_EN (1'b1),             .B_DOUT_EN (1'b1), 
        .A_DOUT_ARST_N (1'b1),         .B_DOUT_ARST_N (1'b1), 
        .A_DOUT_SRST_N (1'b1),         .B_DOUT_SRST_N (1'b1), 
        .A_DOUT_LAT (1'b1),            .B_DOUT_LAT (1'b1),
        .A_WIDTH (width2),             .B_WIDTH (width2), 
        .A_WMODE (1'b0),               .B_WMODE (1'b0),
        .A_EN (1'b1),                  .B_EN (1'b1),
        .BUSY (lsram_512_BUSY_2),
        .SII_LOCK (1'b0)
    );

    RAM1K18 block1 (
        .A_DOUT (readData1),           .B_DOUT (),
        .A_CLK (clk),                  .B_CLK (clk), 
        .A_ARST_N (resetn),            .B_ARST_N (resetn), 
        .A_BLK (3'b111),               .B_BLK (3'b111), 
        .A_DIN (writeData1),           .B_DIN (writeData1), 
        .A_ADDR (writeAddr1),          .B_ADDR (writeAddr1), 
        .A_WEN (wen_a1),               .B_WEN (wen_b1),
        .A_DOUT_CLK (1'b1),            .B_DOUT_CLK (1'b1), 
        .A_DOUT_EN (1'b1),             .B_DOUT_EN (1'b1), 
        .A_DOUT_ARST_N (1'b1),         .B_DOUT_ARST_N (1'b1), 
        .A_DOUT_SRST_N (1'b1),         .B_DOUT_SRST_N (1'b1), 
        .A_DOUT_LAT (1'b1),            .B_DOUT_LAT (1'b1),
        .A_WIDTH (width1),             .B_WIDTH (width1), 
        .A_WMODE (1'b0),               .B_WMODE (1'b0),
        .A_EN (1'b1),                  .B_EN (1'b1),
        .BUSY (lsram_512_BUSY_1),
        .SII_LOCK (1'b0)
    );

    RAM1K18 block0 (
//        .A_DOUT (readData0[35:18]),    .B_DOUT (readData0[17:0]),
        .B_DOUT (readData0[35:18]),    .A_DOUT (readData0[17:0]),
        .A_CLK (clk),                  .B_CLK (clk), 
        .A_ARST_N (resetn),            .B_ARST_N (resetn), 
        .A_BLK (3'b111),               .B_BLK (3'b111), 
//        .A_DIN (writeData0[35:18]),    .B_DIN (writeData0[17:0]), 
        .B_DIN (writeData0[35:18]),    .A_DIN (writeData0[17:0]), 
        .A_ADDR (writeAddr0),          .B_ADDR (writeAddr0), 
        .A_WEN (wen_a0),               .B_WEN (wen_b0),
        .A_DOUT_CLK (1'b1),            .B_DOUT_CLK (1'b1), 
        .A_DOUT_EN (1'b1),             .B_DOUT_EN (1'b1), 
        .A_DOUT_ARST_N (1'b1),         .B_DOUT_ARST_N (1'b1), 
        .A_DOUT_SRST_N (1'b1),         .B_DOUT_SRST_N (1'b1), 
        .A_DOUT_LAT (1'b1),            .B_DOUT_LAT (1'b1),
        .A_WIDTH (width0),             .B_WIDTH (width0), 
        .A_WMODE (1'b0),               .B_WMODE (1'b0),
        .A_EN (1'b1),                  .B_EN (1'b1),
        .BUSY (lsram_512_BUSY_0),
        .SII_LOCK (1'b0)
    );


assign lsram_512_BUSY_all = lsram_512_BUSY_0 | lsram_512_BUSY_1 | lsram_512_BUSY_2 | lsram_512_BUSY_3 | lsram_512_BUSY_4 | lsram_512_BUSY_5 | 
                            lsram_512_BUSY_6 | lsram_512_BUSY_7 | lsram_512_BUSY_8 | lsram_512_BUSY_9 | lsram_512_BUSY_10 | lsram_512_BUSY_11 | 
                            lsram_512_BUSY_12 | lsram_512_BUSY_13 | lsram_512_BUSY_14 | lsram_512_BUSY_15 | lsram_512_BUSY_16 | lsram_512_BUSY_17 | 
                            lsram_512_BUSY_18 | lsram_512_BUSY_19 | lsram_512_BUSY_20 | lsram_512_BUSY_21 | lsram_512_BUSY_22 | lsram_512_BUSY_23 | 
                            lsram_512_BUSY_24 | lsram_512_BUSY_25 | lsram_512_BUSY_26 | lsram_512_BUSY_27 | lsram_512_BUSY_28 | lsram_512_BUSY_29 | 
                            lsram_512_BUSY_30 | lsram_512_BUSY_31 | lsram_512_BUSY_32 | lsram_512_BUSY_33 | lsram_512_BUSY_34 | lsram_512_BUSY_35 | 
                            lsram_512_BUSY_36 | lsram_512_BUSY_37 | lsram_512_BUSY_38 | lsram_512_BUSY_39 | lsram_512_BUSY_40 | lsram_512_BUSY_41 | 
                            lsram_512_BUSY_42 | lsram_512_BUSY_43 | lsram_512_BUSY_44 | lsram_512_BUSY_45 | lsram_512_BUSY_46 | lsram_512_BUSY_47 | 
                            lsram_512_BUSY_48 | lsram_512_BUSY_49 | lsram_512_BUSY_50 | lsram_512_BUSY_51 | lsram_512_BUSY_52 | lsram_512_BUSY_53 |                             
                            lsram_512_BUSY_54 | lsram_512_BUSY_55 | lsram_512_BUSY_56 | lsram_512_BUSY_57 | lsram_512_BUSY_58 | lsram_512_BUSY_59 | 
                            lsram_512_BUSY_60 | lsram_512_BUSY_61 | lsram_512_BUSY_62 | lsram_512_BUSY_63 | lsram_512_BUSY_64 | lsram_512_BUSY_65 | 
                            lsram_512_BUSY_66 | lsram_512_BUSY_67 | lsram_512_BUSY_68;


endmodule // lsram_512to35328x32

