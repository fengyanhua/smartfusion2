`timescale 1 ns/100 ps
// Version: v11.5 SP3 11.5.3.10


module RCOSC_25_50MHZ(
       CLKOUT
    );
output CLKOUT;

    parameter FREQUENCY = 50.0 ;
    
endmodule


module MSS_010(
       CAN_RXBUS_MGPIO3A_H2F_A,
       CAN_RXBUS_MGPIO3A_H2F_B,
       CAN_TX_EBL_MGPIO4A_H2F_A,
       CAN_TX_EBL_MGPIO4A_H2F_B,
       CAN_TXBUS_MGPIO2A_H2F_A,
       CAN_TXBUS_MGPIO2A_H2F_B,
       CLK_CONFIG_APB,
       COMMS_INT,
       CONFIG_PRESET_N,
       EDAC_ERROR,
       F_FM0_RDATA,
       F_FM0_READYOUT,
       F_FM0_RESP,
       F_HM0_ADDR,
       F_HM0_ENABLE,
       F_HM0_SEL,
       F_HM0_SIZE,
       F_HM0_TRANS1,
       F_HM0_WDATA,
       F_HM0_WRITE,
       FAB_CHRGVBUS,
       FAB_DISCHRGVBUS,
       FAB_DMPULLDOWN,
       FAB_DPPULLDOWN,
       FAB_DRVVBUS,
       FAB_IDPULLUP,
       FAB_OPMODE,
       FAB_SUSPENDM,
       FAB_TERMSEL,
       FAB_TXVALID,
       FAB_VCONTROL,
       FAB_VCONTROLLOADM,
       FAB_XCVRSEL,
       FAB_XDATAOUT,
       FACC_GLMUX_SEL,
       FIC32_0_MASTER,
       FIC32_1_MASTER,
       FPGA_RESET_N,
       GTX_CLK,
       H2F_INTERRUPT,
       H2F_NMI,
       H2FCALIB,
       I2C0_SCL_MGPIO31B_H2F_A,
       I2C0_SCL_MGPIO31B_H2F_B,
       I2C0_SDA_MGPIO30B_H2F_A,
       I2C0_SDA_MGPIO30B_H2F_B,
       I2C1_SCL_MGPIO1A_H2F_A,
       I2C1_SCL_MGPIO1A_H2F_B,
       I2C1_SDA_MGPIO0A_H2F_A,
       I2C1_SDA_MGPIO0A_H2F_B,
       MDCF,
       MDOENF,
       MDOF,
       MMUART0_CTS_MGPIO19B_H2F_A,
       MMUART0_CTS_MGPIO19B_H2F_B,
       MMUART0_DCD_MGPIO22B_H2F_A,
       MMUART0_DCD_MGPIO22B_H2F_B,
       MMUART0_DSR_MGPIO20B_H2F_A,
       MMUART0_DSR_MGPIO20B_H2F_B,
       MMUART0_DTR_MGPIO18B_H2F_A,
       MMUART0_DTR_MGPIO18B_H2F_B,
       MMUART0_RI_MGPIO21B_H2F_A,
       MMUART0_RI_MGPIO21B_H2F_B,
       MMUART0_RTS_MGPIO17B_H2F_A,
       MMUART0_RTS_MGPIO17B_H2F_B,
       MMUART0_RXD_MGPIO28B_H2F_A,
       MMUART0_RXD_MGPIO28B_H2F_B,
       MMUART0_SCK_MGPIO29B_H2F_A,
       MMUART0_SCK_MGPIO29B_H2F_B,
       MMUART0_TXD_MGPIO27B_H2F_A,
       MMUART0_TXD_MGPIO27B_H2F_B,
       MMUART1_DTR_MGPIO12B_H2F_A,
       MMUART1_RTS_MGPIO11B_H2F_A,
       MMUART1_RTS_MGPIO11B_H2F_B,
       MMUART1_RXD_MGPIO26B_H2F_A,
       MMUART1_RXD_MGPIO26B_H2F_B,
       MMUART1_SCK_MGPIO25B_H2F_A,
       MMUART1_SCK_MGPIO25B_H2F_B,
       MMUART1_TXD_MGPIO24B_H2F_A,
       MMUART1_TXD_MGPIO24B_H2F_B,
       MPLL_LOCK,
       PER2_FABRIC_PADDR,
       PER2_FABRIC_PENABLE,
       PER2_FABRIC_PSEL,
       PER2_FABRIC_PWDATA,
       PER2_FABRIC_PWRITE,
       RTC_MATCH,
       SLEEPDEEP,
       SLEEPHOLDACK,
       SLEEPING,
       SMBALERT_NO0,
       SMBALERT_NO1,
       SMBSUS_NO0,
       SMBSUS_NO1,
       SPI0_CLK_OUT,
       SPI0_SDI_MGPIO5A_H2F_A,
       SPI0_SDI_MGPIO5A_H2F_B,
       SPI0_SDO_MGPIO6A_H2F_A,
       SPI0_SDO_MGPIO6A_H2F_B,
       SPI0_SS0_MGPIO7A_H2F_A,
       SPI0_SS0_MGPIO7A_H2F_B,
       SPI0_SS1_MGPIO8A_H2F_A,
       SPI0_SS1_MGPIO8A_H2F_B,
       SPI0_SS2_MGPIO9A_H2F_A,
       SPI0_SS2_MGPIO9A_H2F_B,
       SPI0_SS3_MGPIO10A_H2F_A,
       SPI0_SS3_MGPIO10A_H2F_B,
       SPI0_SS4_MGPIO19A_H2F_A,
       SPI0_SS5_MGPIO20A_H2F_A,
       SPI0_SS6_MGPIO21A_H2F_A,
       SPI0_SS7_MGPIO22A_H2F_A,
       SPI1_CLK_OUT,
       SPI1_SDI_MGPIO11A_H2F_A,
       SPI1_SDI_MGPIO11A_H2F_B,
       SPI1_SDO_MGPIO12A_H2F_A,
       SPI1_SDO_MGPIO12A_H2F_B,
       SPI1_SS0_MGPIO13A_H2F_A,
       SPI1_SS0_MGPIO13A_H2F_B,
       SPI1_SS1_MGPIO14A_H2F_A,
       SPI1_SS1_MGPIO14A_H2F_B,
       SPI1_SS2_MGPIO15A_H2F_A,
       SPI1_SS2_MGPIO15A_H2F_B,
       SPI1_SS3_MGPIO16A_H2F_A,
       SPI1_SS3_MGPIO16A_H2F_B,
       SPI1_SS4_MGPIO17A_H2F_A,
       SPI1_SS5_MGPIO18A_H2F_A,
       SPI1_SS6_MGPIO23A_H2F_A,
       SPI1_SS7_MGPIO24A_H2F_A,
       TCGF,
       TRACECLK,
       TRACEDATA,
       TX_CLK,
       TX_ENF,
       TX_ERRF,
       TXCTL_EN_RIF,
       TXD_RIF,
       TXDF,
       TXEV,
       WDOGTIMEOUT,
       F_ARREADY_HREADYOUT1,
       F_AWREADY_HREADYOUT0,
       F_BID,
       F_BRESP_HRESP0,
       F_BVALID,
       F_RDATA_HRDATA01,
       F_RID,
       F_RLAST,
       F_RRESP_HRESP1,
       F_RVALID,
       F_WREADY,
       MDDR_FABRIC_PRDATA,
       MDDR_FABRIC_PREADY,
       MDDR_FABRIC_PSLVERR,
       CAN_RXBUS_F2H_SCP,
       CAN_TX_EBL_F2H_SCP,
       CAN_TXBUS_F2H_SCP,
       COLF,
       CRSF,
       F2_DMAREADY,
       F2H_INTERRUPT,
       F2HCALIB,
       F_DMAREADY,
       F_FM0_ADDR,
       F_FM0_ENABLE,
       F_FM0_MASTLOCK,
       F_FM0_READY,
       F_FM0_SEL,
       F_FM0_SIZE,
       F_FM0_TRANS1,
       F_FM0_WDATA,
       F_FM0_WRITE,
       F_HM0_RDATA,
       F_HM0_READY,
       F_HM0_RESP,
       FAB_AVALID,
       FAB_HOSTDISCON,
       FAB_IDDIG,
       FAB_LINESTATE,
       FAB_M3_RESET_N,
       FAB_PLL_LOCK,
       FAB_RXACTIVE,
       FAB_RXERROR,
       FAB_RXVALID,
       FAB_RXVALIDH,
       FAB_SESSEND,
       FAB_TXREADY,
       FAB_VBUSVALID,
       FAB_VSTATUS,
       FAB_XDATAIN,
       GTX_CLKPF,
       I2C0_BCLK,
       I2C0_SCL_F2H_SCP,
       I2C0_SDA_F2H_SCP,
       I2C1_BCLK,
       I2C1_SCL_F2H_SCP,
       I2C1_SDA_F2H_SCP,
       MDIF,
       MGPIO0A_F2H_GPIN,
       MGPIO10A_F2H_GPIN,
       MGPIO11A_F2H_GPIN,
       MGPIO11B_F2H_GPIN,
       MGPIO12A_F2H_GPIN,
       MGPIO13A_F2H_GPIN,
       MGPIO14A_F2H_GPIN,
       MGPIO15A_F2H_GPIN,
       MGPIO16A_F2H_GPIN,
       MGPIO17B_F2H_GPIN,
       MGPIO18B_F2H_GPIN,
       MGPIO19B_F2H_GPIN,
       MGPIO1A_F2H_GPIN,
       MGPIO20B_F2H_GPIN,
       MGPIO21B_F2H_GPIN,
       MGPIO22B_F2H_GPIN,
       MGPIO24B_F2H_GPIN,
       MGPIO25B_F2H_GPIN,
       MGPIO26B_F2H_GPIN,
       MGPIO27B_F2H_GPIN,
       MGPIO28B_F2H_GPIN,
       MGPIO29B_F2H_GPIN,
       MGPIO2A_F2H_GPIN,
       MGPIO30B_F2H_GPIN,
       MGPIO31B_F2H_GPIN,
       MGPIO3A_F2H_GPIN,
       MGPIO4A_F2H_GPIN,
       MGPIO5A_F2H_GPIN,
       MGPIO6A_F2H_GPIN,
       MGPIO7A_F2H_GPIN,
       MGPIO8A_F2H_GPIN,
       MGPIO9A_F2H_GPIN,
       MMUART0_CTS_F2H_SCP,
       MMUART0_DCD_F2H_SCP,
       MMUART0_DSR_F2H_SCP,
       MMUART0_DTR_F2H_SCP,
       MMUART0_RI_F2H_SCP,
       MMUART0_RTS_F2H_SCP,
       MMUART0_RXD_F2H_SCP,
       MMUART0_SCK_F2H_SCP,
       MMUART0_TXD_F2H_SCP,
       MMUART1_CTS_F2H_SCP,
       MMUART1_DCD_F2H_SCP,
       MMUART1_DSR_F2H_SCP,
       MMUART1_RI_F2H_SCP,
       MMUART1_RTS_F2H_SCP,
       MMUART1_RXD_F2H_SCP,
       MMUART1_SCK_F2H_SCP,
       MMUART1_TXD_F2H_SCP,
       PER2_FABRIC_PRDATA,
       PER2_FABRIC_PREADY,
       PER2_FABRIC_PSLVERR,
       RCGF,
       RX_CLKPF,
       RX_DVF,
       RX_ERRF,
       RX_EV,
       RXDF,
       SLEEPHOLDREQ,
       SMBALERT_NI0,
       SMBALERT_NI1,
       SMBSUS_NI0,
       SMBSUS_NI1,
       SPI0_CLK_IN,
       SPI0_SDI_F2H_SCP,
       SPI0_SDO_F2H_SCP,
       SPI0_SS0_F2H_SCP,
       SPI0_SS1_F2H_SCP,
       SPI0_SS2_F2H_SCP,
       SPI0_SS3_F2H_SCP,
       SPI1_CLK_IN,
       SPI1_SDI_F2H_SCP,
       SPI1_SDO_F2H_SCP,
       SPI1_SS0_F2H_SCP,
       SPI1_SS1_F2H_SCP,
       SPI1_SS2_F2H_SCP,
       SPI1_SS3_F2H_SCP,
       TX_CLKPF,
       USER_MSS_GPIO_RESET_N,
       USER_MSS_RESET_N,
       XCLK_FAB,
       CLK_BASE,
       CLK_MDDR_APB,
       F_ARADDR_HADDR1,
       F_ARBURST_HTRANS1,
       F_ARID_HSEL1,
       F_ARLEN_HBURST1,
       F_ARLOCK_HMASTLOCK1,
       F_ARSIZE_HSIZE1,
       F_ARVALID_HWRITE1,
       F_AWADDR_HADDR0,
       F_AWBURST_HTRANS0,
       F_AWID_HSEL0,
       F_AWLEN_HBURST0,
       F_AWLOCK_HMASTLOCK0,
       F_AWSIZE_HSIZE0,
       F_AWVALID_HWRITE0,
       F_BREADY,
       F_RMW_AXI,
       F_RREADY,
       F_WDATA_HWDATA01,
       F_WID_HREADY01,
       F_WLAST,
       F_WSTRB,
       F_WVALID,
       FPGA_MDDR_ARESET_N,
       MDDR_FABRIC_PADDR,
       MDDR_FABRIC_PENABLE,
       MDDR_FABRIC_PSEL,
       MDDR_FABRIC_PWDATA,
       MDDR_FABRIC_PWRITE,
       PRESET_N,
       CAN_RXBUS_USBA_DATA1_MGPIO3A_IN,
       CAN_TX_EBL_USBA_DATA2_MGPIO4A_IN,
       CAN_TXBUS_USBA_DATA0_MGPIO2A_IN,
       DM_IN,
       DRAM_DQ_IN,
       DRAM_DQS_IN,
       DRAM_FIFO_WE_IN,
       I2C0_SCL_USBC_DATA1_MGPIO31B_IN,
       I2C0_SDA_USBC_DATA0_MGPIO30B_IN,
       I2C1_SCL_USBA_DATA4_MGPIO1A_IN,
       I2C1_SDA_USBA_DATA3_MGPIO0A_IN,
       MMUART0_CTS_USBC_DATA7_MGPIO19B_IN,
       MMUART0_DCD_MGPIO22B_IN,
       MMUART0_DSR_MGPIO20B_IN,
       MMUART0_DTR_USBC_DATA6_MGPIO18B_IN,
       MMUART0_RI_MGPIO21B_IN,
       MMUART0_RTS_USBC_DATA5_MGPIO17B_IN,
       MMUART0_RXD_USBC_STP_MGPIO28B_IN,
       MMUART0_SCK_USBC_NXT_MGPIO29B_IN,
       MMUART0_TXD_USBC_DIR_MGPIO27B_IN,
       MMUART1_RXD_USBC_DATA3_MGPIO26B_IN,
       MMUART1_SCK_USBC_DATA4_MGPIO25B_IN,
       MMUART1_TXD_USBC_DATA2_MGPIO24B_IN,
       RGMII_GTX_CLK_RMII_CLK_USBB_XCLK_IN,
       RGMII_MDC_RMII_MDC_IN,
       RGMII_MDIO_RMII_MDIO_USBB_DATA7_IN,
       RGMII_RX_CLK_IN,
       RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_IN,
       RGMII_RXD0_RMII_RXD0_USBB_DATA0_IN,
       RGMII_RXD1_RMII_RXD1_USBB_DATA1_IN,
       RGMII_RXD2_RMII_RX_ER_USBB_DATA3_IN,
       RGMII_RXD3_USBB_DATA4_IN,
       RGMII_TX_CLK_IN,
       RGMII_TX_CTL_RMII_TX_EN_USBB_NXT_IN,
       RGMII_TXD0_RMII_TXD0_USBB_DIR_IN,
       RGMII_TXD1_RMII_TXD1_USBB_STP_IN,
       RGMII_TXD2_USBB_DATA5_IN,
       RGMII_TXD3_USBB_DATA6_IN,
       SPI0_SCK_USBA_XCLK_IN,
       SPI0_SDI_USBA_DIR_MGPIO5A_IN,
       SPI0_SDO_USBA_STP_MGPIO6A_IN,
       SPI0_SS0_USBA_NXT_MGPIO7A_IN,
       SPI0_SS1_USBA_DATA5_MGPIO8A_IN,
       SPI0_SS2_USBA_DATA6_MGPIO9A_IN,
       SPI0_SS3_USBA_DATA7_MGPIO10A_IN,
       SPI1_SCK_IN,
       SPI1_SDI_MGPIO11A_IN,
       SPI1_SDO_MGPIO12A_IN,
       SPI1_SS0_MGPIO13A_IN,
       SPI1_SS1_MGPIO14A_IN,
       SPI1_SS2_MGPIO15A_IN,
       SPI1_SS3_MGPIO16A_IN,
       SPI1_SS4_MGPIO17A_IN,
       SPI1_SS5_MGPIO18A_IN,
       SPI1_SS6_MGPIO23A_IN,
       SPI1_SS7_MGPIO24A_IN,
       USBC_XCLK_IN,
       CAN_RXBUS_USBA_DATA1_MGPIO3A_OUT,
       CAN_TX_EBL_USBA_DATA2_MGPIO4A_OUT,
       CAN_TXBUS_USBA_DATA0_MGPIO2A_OUT,
       DRAM_ADDR,
       DRAM_BA,
       DRAM_CASN,
       DRAM_CKE,
       DRAM_CLK,
       DRAM_CSN,
       DRAM_DM_RDQS_OUT,
       DRAM_DQ_OUT,
       DRAM_DQS_OUT,
       DRAM_FIFO_WE_OUT,
       DRAM_ODT,
       DRAM_RASN,
       DRAM_RSTN,
       DRAM_WEN,
       I2C0_SCL_USBC_DATA1_MGPIO31B_OUT,
       I2C0_SDA_USBC_DATA0_MGPIO30B_OUT,
       I2C1_SCL_USBA_DATA4_MGPIO1A_OUT,
       I2C1_SDA_USBA_DATA3_MGPIO0A_OUT,
       MMUART0_CTS_USBC_DATA7_MGPIO19B_OUT,
       MMUART0_DCD_MGPIO22B_OUT,
       MMUART0_DSR_MGPIO20B_OUT,
       MMUART0_DTR_USBC_DATA6_MGPIO18B_OUT,
       MMUART0_RI_MGPIO21B_OUT,
       MMUART0_RTS_USBC_DATA5_MGPIO17B_OUT,
       MMUART0_RXD_USBC_STP_MGPIO28B_OUT,
       MMUART0_SCK_USBC_NXT_MGPIO29B_OUT,
       MMUART0_TXD_USBC_DIR_MGPIO27B_OUT,
       MMUART1_RXD_USBC_DATA3_MGPIO26B_OUT,
       MMUART1_SCK_USBC_DATA4_MGPIO25B_OUT,
       MMUART1_TXD_USBC_DATA2_MGPIO24B_OUT,
       RGMII_GTX_CLK_RMII_CLK_USBB_XCLK_OUT,
       RGMII_MDC_RMII_MDC_OUT,
       RGMII_MDIO_RMII_MDIO_USBB_DATA7_OUT,
       RGMII_RX_CLK_OUT,
       RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_OUT,
       RGMII_RXD0_RMII_RXD0_USBB_DATA0_OUT,
       RGMII_RXD1_RMII_RXD1_USBB_DATA1_OUT,
       RGMII_RXD2_RMII_RX_ER_USBB_DATA3_OUT,
       RGMII_RXD3_USBB_DATA4_OUT,
       RGMII_TX_CLK_OUT,
       RGMII_TX_CTL_RMII_TX_EN_USBB_NXT_OUT,
       RGMII_TXD0_RMII_TXD0_USBB_DIR_OUT,
       RGMII_TXD1_RMII_TXD1_USBB_STP_OUT,
       RGMII_TXD2_USBB_DATA5_OUT,
       RGMII_TXD3_USBB_DATA6_OUT,
       SPI0_SCK_USBA_XCLK_OUT,
       SPI0_SDI_USBA_DIR_MGPIO5A_OUT,
       SPI0_SDO_USBA_STP_MGPIO6A_OUT,
       SPI0_SS0_USBA_NXT_MGPIO7A_OUT,
       SPI0_SS1_USBA_DATA5_MGPIO8A_OUT,
       SPI0_SS2_USBA_DATA6_MGPIO9A_OUT,
       SPI0_SS3_USBA_DATA7_MGPIO10A_OUT,
       SPI1_SCK_OUT,
       SPI1_SDI_MGPIO11A_OUT,
       SPI1_SDO_MGPIO12A_OUT,
       SPI1_SS0_MGPIO13A_OUT,
       SPI1_SS1_MGPIO14A_OUT,
       SPI1_SS2_MGPIO15A_OUT,
       SPI1_SS3_MGPIO16A_OUT,
       SPI1_SS4_MGPIO17A_OUT,
       SPI1_SS5_MGPIO18A_OUT,
       SPI1_SS6_MGPIO23A_OUT,
       SPI1_SS7_MGPIO24A_OUT,
       USBC_XCLK_OUT,
       CAN_RXBUS_USBA_DATA1_MGPIO3A_OE,
       CAN_TX_EBL_USBA_DATA2_MGPIO4A_OE,
       CAN_TXBUS_USBA_DATA0_MGPIO2A_OE,
       DM_OE,
       DRAM_DQ_OE,
       DRAM_DQS_OE,
       I2C0_SCL_USBC_DATA1_MGPIO31B_OE,
       I2C0_SDA_USBC_DATA0_MGPIO30B_OE,
       I2C1_SCL_USBA_DATA4_MGPIO1A_OE,
       I2C1_SDA_USBA_DATA3_MGPIO0A_OE,
       MMUART0_CTS_USBC_DATA7_MGPIO19B_OE,
       MMUART0_DCD_MGPIO22B_OE,
       MMUART0_DSR_MGPIO20B_OE,
       MMUART0_DTR_USBC_DATA6_MGPIO18B_OE,
       MMUART0_RI_MGPIO21B_OE,
       MMUART0_RTS_USBC_DATA5_MGPIO17B_OE,
       MMUART0_RXD_USBC_STP_MGPIO28B_OE,
       MMUART0_SCK_USBC_NXT_MGPIO29B_OE,
       MMUART0_TXD_USBC_DIR_MGPIO27B_OE,
       MMUART1_RXD_USBC_DATA3_MGPIO26B_OE,
       MMUART1_SCK_USBC_DATA4_MGPIO25B_OE,
       MMUART1_TXD_USBC_DATA2_MGPIO24B_OE,
       RGMII_GTX_CLK_RMII_CLK_USBB_XCLK_OE,
       RGMII_MDC_RMII_MDC_OE,
       RGMII_MDIO_RMII_MDIO_USBB_DATA7_OE,
       RGMII_RX_CLK_OE,
       RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_OE,
       RGMII_RXD0_RMII_RXD0_USBB_DATA0_OE,
       RGMII_RXD1_RMII_RXD1_USBB_DATA1_OE,
       RGMII_RXD2_RMII_RX_ER_USBB_DATA3_OE,
       RGMII_RXD3_USBB_DATA4_OE,
       RGMII_TX_CLK_OE,
       RGMII_TX_CTL_RMII_TX_EN_USBB_NXT_OE,
       RGMII_TXD0_RMII_TXD0_USBB_DIR_OE,
       RGMII_TXD1_RMII_TXD1_USBB_STP_OE,
       RGMII_TXD2_USBB_DATA5_OE,
       RGMII_TXD3_USBB_DATA6_OE,
       SPI0_SCK_USBA_XCLK_OE,
       SPI0_SDI_USBA_DIR_MGPIO5A_OE,
       SPI0_SDO_USBA_STP_MGPIO6A_OE,
       SPI0_SS0_USBA_NXT_MGPIO7A_OE,
       SPI0_SS1_USBA_DATA5_MGPIO8A_OE,
       SPI0_SS2_USBA_DATA6_MGPIO9A_OE,
       SPI0_SS3_USBA_DATA7_MGPIO10A_OE,
       SPI1_SCK_OE,
       SPI1_SDI_MGPIO11A_OE,
       SPI1_SDO_MGPIO12A_OE,
       SPI1_SS0_MGPIO13A_OE,
       SPI1_SS1_MGPIO14A_OE,
       SPI1_SS2_MGPIO15A_OE,
       SPI1_SS3_MGPIO16A_OE,
       SPI1_SS4_MGPIO17A_OE,
       SPI1_SS5_MGPIO18A_OE,
       SPI1_SS6_MGPIO23A_OE,
       SPI1_SS7_MGPIO24A_OE,
       USBC_XCLK_OE
    );
output CAN_RXBUS_MGPIO3A_H2F_A;
output CAN_RXBUS_MGPIO3A_H2F_B;
output CAN_TX_EBL_MGPIO4A_H2F_A;
output CAN_TX_EBL_MGPIO4A_H2F_B;
output CAN_TXBUS_MGPIO2A_H2F_A;
output CAN_TXBUS_MGPIO2A_H2F_B;
output CLK_CONFIG_APB;
output COMMS_INT;
output CONFIG_PRESET_N;
output [7:0] EDAC_ERROR;
output [31:0] F_FM0_RDATA;
output F_FM0_READYOUT;
output F_FM0_RESP;
output [31:0] F_HM0_ADDR;
output F_HM0_ENABLE;
output F_HM0_SEL;
output [1:0] F_HM0_SIZE;
output F_HM0_TRANS1;
output [31:0] F_HM0_WDATA;
output F_HM0_WRITE;
output FAB_CHRGVBUS;
output FAB_DISCHRGVBUS;
output FAB_DMPULLDOWN;
output FAB_DPPULLDOWN;
output FAB_DRVVBUS;
output FAB_IDPULLUP;
output [1:0] FAB_OPMODE;
output FAB_SUSPENDM;
output FAB_TERMSEL;
output FAB_TXVALID;
output [3:0] FAB_VCONTROL;
output FAB_VCONTROLLOADM;
output [1:0] FAB_XCVRSEL;
output [7:0] FAB_XDATAOUT;
output FACC_GLMUX_SEL;
output [1:0] FIC32_0_MASTER;
output [1:0] FIC32_1_MASTER;
output FPGA_RESET_N;
output GTX_CLK;
output [15:0] H2F_INTERRUPT;
output H2F_NMI;
output H2FCALIB;
output I2C0_SCL_MGPIO31B_H2F_A;
output I2C0_SCL_MGPIO31B_H2F_B;
output I2C0_SDA_MGPIO30B_H2F_A;
output I2C0_SDA_MGPIO30B_H2F_B;
output I2C1_SCL_MGPIO1A_H2F_A;
output I2C1_SCL_MGPIO1A_H2F_B;
output I2C1_SDA_MGPIO0A_H2F_A;
output I2C1_SDA_MGPIO0A_H2F_B;
output MDCF;
output MDOENF;
output MDOF;
output MMUART0_CTS_MGPIO19B_H2F_A;
output MMUART0_CTS_MGPIO19B_H2F_B;
output MMUART0_DCD_MGPIO22B_H2F_A;
output MMUART0_DCD_MGPIO22B_H2F_B;
output MMUART0_DSR_MGPIO20B_H2F_A;
output MMUART0_DSR_MGPIO20B_H2F_B;
output MMUART0_DTR_MGPIO18B_H2F_A;
output MMUART0_DTR_MGPIO18B_H2F_B;
output MMUART0_RI_MGPIO21B_H2F_A;
output MMUART0_RI_MGPIO21B_H2F_B;
output MMUART0_RTS_MGPIO17B_H2F_A;
output MMUART0_RTS_MGPIO17B_H2F_B;
output MMUART0_RXD_MGPIO28B_H2F_A;
output MMUART0_RXD_MGPIO28B_H2F_B;
output MMUART0_SCK_MGPIO29B_H2F_A;
output MMUART0_SCK_MGPIO29B_H2F_B;
output MMUART0_TXD_MGPIO27B_H2F_A;
output MMUART0_TXD_MGPIO27B_H2F_B;
output MMUART1_DTR_MGPIO12B_H2F_A;
output MMUART1_RTS_MGPIO11B_H2F_A;
output MMUART1_RTS_MGPIO11B_H2F_B;
output MMUART1_RXD_MGPIO26B_H2F_A;
output MMUART1_RXD_MGPIO26B_H2F_B;
output MMUART1_SCK_MGPIO25B_H2F_A;
output MMUART1_SCK_MGPIO25B_H2F_B;
output MMUART1_TXD_MGPIO24B_H2F_A;
output MMUART1_TXD_MGPIO24B_H2F_B;
output MPLL_LOCK;
output [15:2] PER2_FABRIC_PADDR;
output PER2_FABRIC_PENABLE;
output PER2_FABRIC_PSEL;
output [31:0] PER2_FABRIC_PWDATA;
output PER2_FABRIC_PWRITE;
output RTC_MATCH;
output SLEEPDEEP;
output SLEEPHOLDACK;
output SLEEPING;
output SMBALERT_NO0;
output SMBALERT_NO1;
output SMBSUS_NO0;
output SMBSUS_NO1;
output SPI0_CLK_OUT;
output SPI0_SDI_MGPIO5A_H2F_A;
output SPI0_SDI_MGPIO5A_H2F_B;
output SPI0_SDO_MGPIO6A_H2F_A;
output SPI0_SDO_MGPIO6A_H2F_B;
output SPI0_SS0_MGPIO7A_H2F_A;
output SPI0_SS0_MGPIO7A_H2F_B;
output SPI0_SS1_MGPIO8A_H2F_A;
output SPI0_SS1_MGPIO8A_H2F_B;
output SPI0_SS2_MGPIO9A_H2F_A;
output SPI0_SS2_MGPIO9A_H2F_B;
output SPI0_SS3_MGPIO10A_H2F_A;
output SPI0_SS3_MGPIO10A_H2F_B;
output SPI0_SS4_MGPIO19A_H2F_A;
output SPI0_SS5_MGPIO20A_H2F_A;
output SPI0_SS6_MGPIO21A_H2F_A;
output SPI0_SS7_MGPIO22A_H2F_A;
output SPI1_CLK_OUT;
output SPI1_SDI_MGPIO11A_H2F_A;
output SPI1_SDI_MGPIO11A_H2F_B;
output SPI1_SDO_MGPIO12A_H2F_A;
output SPI1_SDO_MGPIO12A_H2F_B;
output SPI1_SS0_MGPIO13A_H2F_A;
output SPI1_SS0_MGPIO13A_H2F_B;
output SPI1_SS1_MGPIO14A_H2F_A;
output SPI1_SS1_MGPIO14A_H2F_B;
output SPI1_SS2_MGPIO15A_H2F_A;
output SPI1_SS2_MGPIO15A_H2F_B;
output SPI1_SS3_MGPIO16A_H2F_A;
output SPI1_SS3_MGPIO16A_H2F_B;
output SPI1_SS4_MGPIO17A_H2F_A;
output SPI1_SS5_MGPIO18A_H2F_A;
output SPI1_SS6_MGPIO23A_H2F_A;
output SPI1_SS7_MGPIO24A_H2F_A;
output [9:0] TCGF;
output TRACECLK;
output [3:0] TRACEDATA;
output TX_CLK;
output TX_ENF;
output TX_ERRF;
output TXCTL_EN_RIF;
output [3:0] TXD_RIF;
output [7:0] TXDF;
output TXEV;
output WDOGTIMEOUT;
output F_ARREADY_HREADYOUT1;
output F_AWREADY_HREADYOUT0;
output [3:0] F_BID;
output [1:0] F_BRESP_HRESP0;
output F_BVALID;
output [63:0] F_RDATA_HRDATA01;
output [3:0] F_RID;
output F_RLAST;
output [1:0] F_RRESP_HRESP1;
output F_RVALID;
output F_WREADY;
output [15:0] MDDR_FABRIC_PRDATA;
output MDDR_FABRIC_PREADY;
output MDDR_FABRIC_PSLVERR;
input  CAN_RXBUS_F2H_SCP;
input  CAN_TX_EBL_F2H_SCP;
input  CAN_TXBUS_F2H_SCP;
input  COLF;
input  CRSF;
input  [1:0] F2_DMAREADY;
input  [15:0] F2H_INTERRUPT;
input  F2HCALIB;
input  [1:0] F_DMAREADY;
input  [31:0] F_FM0_ADDR;
input  F_FM0_ENABLE;
input  F_FM0_MASTLOCK;
input  F_FM0_READY;
input  F_FM0_SEL;
input  [1:0] F_FM0_SIZE;
input  F_FM0_TRANS1;
input  [31:0] F_FM0_WDATA;
input  F_FM0_WRITE;
input  [31:0] F_HM0_RDATA;
input  F_HM0_READY;
input  F_HM0_RESP;
input  FAB_AVALID;
input  FAB_HOSTDISCON;
input  FAB_IDDIG;
input  [1:0] FAB_LINESTATE;
input  FAB_M3_RESET_N;
input  FAB_PLL_LOCK;
input  FAB_RXACTIVE;
input  FAB_RXERROR;
input  FAB_RXVALID;
input  FAB_RXVALIDH;
input  FAB_SESSEND;
input  FAB_TXREADY;
input  FAB_VBUSVALID;
input  [7:0] FAB_VSTATUS;
input  [7:0] FAB_XDATAIN;
input  GTX_CLKPF;
input  I2C0_BCLK;
input  I2C0_SCL_F2H_SCP;
input  I2C0_SDA_F2H_SCP;
input  I2C1_BCLK;
input  I2C1_SCL_F2H_SCP;
input  I2C1_SDA_F2H_SCP;
input  MDIF;
input  MGPIO0A_F2H_GPIN;
input  MGPIO10A_F2H_GPIN;
input  MGPIO11A_F2H_GPIN;
input  MGPIO11B_F2H_GPIN;
input  MGPIO12A_F2H_GPIN;
input  MGPIO13A_F2H_GPIN;
input  MGPIO14A_F2H_GPIN;
input  MGPIO15A_F2H_GPIN;
input  MGPIO16A_F2H_GPIN;
input  MGPIO17B_F2H_GPIN;
input  MGPIO18B_F2H_GPIN;
input  MGPIO19B_F2H_GPIN;
input  MGPIO1A_F2H_GPIN;
input  MGPIO20B_F2H_GPIN;
input  MGPIO21B_F2H_GPIN;
input  MGPIO22B_F2H_GPIN;
input  MGPIO24B_F2H_GPIN;
input  MGPIO25B_F2H_GPIN;
input  MGPIO26B_F2H_GPIN;
input  MGPIO27B_F2H_GPIN;
input  MGPIO28B_F2H_GPIN;
input  MGPIO29B_F2H_GPIN;
input  MGPIO2A_F2H_GPIN;
input  MGPIO30B_F2H_GPIN;
input  MGPIO31B_F2H_GPIN;
input  MGPIO3A_F2H_GPIN;
input  MGPIO4A_F2H_GPIN;
input  MGPIO5A_F2H_GPIN;
input  MGPIO6A_F2H_GPIN;
input  MGPIO7A_F2H_GPIN;
input  MGPIO8A_F2H_GPIN;
input  MGPIO9A_F2H_GPIN;
input  MMUART0_CTS_F2H_SCP;
input  MMUART0_DCD_F2H_SCP;
input  MMUART0_DSR_F2H_SCP;
input  MMUART0_DTR_F2H_SCP;
input  MMUART0_RI_F2H_SCP;
input  MMUART0_RTS_F2H_SCP;
input  MMUART0_RXD_F2H_SCP;
input  MMUART0_SCK_F2H_SCP;
input  MMUART0_TXD_F2H_SCP;
input  MMUART1_CTS_F2H_SCP;
input  MMUART1_DCD_F2H_SCP;
input  MMUART1_DSR_F2H_SCP;
input  MMUART1_RI_F2H_SCP;
input  MMUART1_RTS_F2H_SCP;
input  MMUART1_RXD_F2H_SCP;
input  MMUART1_SCK_F2H_SCP;
input  MMUART1_TXD_F2H_SCP;
input  [31:0] PER2_FABRIC_PRDATA;
input  PER2_FABRIC_PREADY;
input  PER2_FABRIC_PSLVERR;
input  [9:0] RCGF;
input  RX_CLKPF;
input  RX_DVF;
input  RX_ERRF;
input  RX_EV;
input  [7:0] RXDF;
input  SLEEPHOLDREQ;
input  SMBALERT_NI0;
input  SMBALERT_NI1;
input  SMBSUS_NI0;
input  SMBSUS_NI1;
input  SPI0_CLK_IN;
input  SPI0_SDI_F2H_SCP;
input  SPI0_SDO_F2H_SCP;
input  SPI0_SS0_F2H_SCP;
input  SPI0_SS1_F2H_SCP;
input  SPI0_SS2_F2H_SCP;
input  SPI0_SS3_F2H_SCP;
input  SPI1_CLK_IN;
input  SPI1_SDI_F2H_SCP;
input  SPI1_SDO_F2H_SCP;
input  SPI1_SS0_F2H_SCP;
input  SPI1_SS1_F2H_SCP;
input  SPI1_SS2_F2H_SCP;
input  SPI1_SS3_F2H_SCP;
input  TX_CLKPF;
input  USER_MSS_GPIO_RESET_N;
input  USER_MSS_RESET_N;
input  XCLK_FAB;
input  CLK_BASE;
input  CLK_MDDR_APB;
input  [31:0] F_ARADDR_HADDR1;
input  [1:0] F_ARBURST_HTRANS1;
input  [3:0] F_ARID_HSEL1;
input  [3:0] F_ARLEN_HBURST1;
input  [1:0] F_ARLOCK_HMASTLOCK1;
input  [1:0] F_ARSIZE_HSIZE1;
input  F_ARVALID_HWRITE1;
input  [31:0] F_AWADDR_HADDR0;
input  [1:0] F_AWBURST_HTRANS0;
input  [3:0] F_AWID_HSEL0;
input  [3:0] F_AWLEN_HBURST0;
input  [1:0] F_AWLOCK_HMASTLOCK0;
input  [1:0] F_AWSIZE_HSIZE0;
input  F_AWVALID_HWRITE0;
input  F_BREADY;
input  F_RMW_AXI;
input  F_RREADY;
input  [63:0] F_WDATA_HWDATA01;
input  [3:0] F_WID_HREADY01;
input  F_WLAST;
input  [7:0] F_WSTRB;
input  F_WVALID;
input  FPGA_MDDR_ARESET_N;
input  [10:2] MDDR_FABRIC_PADDR;
input  MDDR_FABRIC_PENABLE;
input  MDDR_FABRIC_PSEL;
input  [15:0] MDDR_FABRIC_PWDATA;
input  MDDR_FABRIC_PWRITE;
input  PRESET_N;
input  CAN_RXBUS_USBA_DATA1_MGPIO3A_IN;
input  CAN_TX_EBL_USBA_DATA2_MGPIO4A_IN;
input  CAN_TXBUS_USBA_DATA0_MGPIO2A_IN;
input  [2:0] DM_IN;
input  [17:0] DRAM_DQ_IN;
input  [2:0] DRAM_DQS_IN;
input  [1:0] DRAM_FIFO_WE_IN;
input  I2C0_SCL_USBC_DATA1_MGPIO31B_IN;
input  I2C0_SDA_USBC_DATA0_MGPIO30B_IN;
input  I2C1_SCL_USBA_DATA4_MGPIO1A_IN;
input  I2C1_SDA_USBA_DATA3_MGPIO0A_IN;
input  MMUART0_CTS_USBC_DATA7_MGPIO19B_IN;
input  MMUART0_DCD_MGPIO22B_IN;
input  MMUART0_DSR_MGPIO20B_IN;
input  MMUART0_DTR_USBC_DATA6_MGPIO18B_IN;
input  MMUART0_RI_MGPIO21B_IN;
input  MMUART0_RTS_USBC_DATA5_MGPIO17B_IN;
input  MMUART0_RXD_USBC_STP_MGPIO28B_IN;
input  MMUART0_SCK_USBC_NXT_MGPIO29B_IN;
input  MMUART0_TXD_USBC_DIR_MGPIO27B_IN;
input  MMUART1_RXD_USBC_DATA3_MGPIO26B_IN;
input  MMUART1_SCK_USBC_DATA4_MGPIO25B_IN;
input  MMUART1_TXD_USBC_DATA2_MGPIO24B_IN;
input  RGMII_GTX_CLK_RMII_CLK_USBB_XCLK_IN;
input  RGMII_MDC_RMII_MDC_IN;
input  RGMII_MDIO_RMII_MDIO_USBB_DATA7_IN;
input  RGMII_RX_CLK_IN;
input  RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_IN;
input  RGMII_RXD0_RMII_RXD0_USBB_DATA0_IN;
input  RGMII_RXD1_RMII_RXD1_USBB_DATA1_IN;
input  RGMII_RXD2_RMII_RX_ER_USBB_DATA3_IN;
input  RGMII_RXD3_USBB_DATA4_IN;
input  RGMII_TX_CLK_IN;
input  RGMII_TX_CTL_RMII_TX_EN_USBB_NXT_IN;
input  RGMII_TXD0_RMII_TXD0_USBB_DIR_IN;
input  RGMII_TXD1_RMII_TXD1_USBB_STP_IN;
input  RGMII_TXD2_USBB_DATA5_IN;
input  RGMII_TXD3_USBB_DATA6_IN;
input  SPI0_SCK_USBA_XCLK_IN;
input  SPI0_SDI_USBA_DIR_MGPIO5A_IN;
input  SPI0_SDO_USBA_STP_MGPIO6A_IN;
input  SPI0_SS0_USBA_NXT_MGPIO7A_IN;
input  SPI0_SS1_USBA_DATA5_MGPIO8A_IN;
input  SPI0_SS2_USBA_DATA6_MGPIO9A_IN;
input  SPI0_SS3_USBA_DATA7_MGPIO10A_IN;
input  SPI1_SCK_IN;
input  SPI1_SDI_MGPIO11A_IN;
input  SPI1_SDO_MGPIO12A_IN;
input  SPI1_SS0_MGPIO13A_IN;
input  SPI1_SS1_MGPIO14A_IN;
input  SPI1_SS2_MGPIO15A_IN;
input  SPI1_SS3_MGPIO16A_IN;
input  SPI1_SS4_MGPIO17A_IN;
input  SPI1_SS5_MGPIO18A_IN;
input  SPI1_SS6_MGPIO23A_IN;
input  SPI1_SS7_MGPIO24A_IN;
input  USBC_XCLK_IN;
output CAN_RXBUS_USBA_DATA1_MGPIO3A_OUT;
output CAN_TX_EBL_USBA_DATA2_MGPIO4A_OUT;
output CAN_TXBUS_USBA_DATA0_MGPIO2A_OUT;
output [15:0] DRAM_ADDR;
output [2:0] DRAM_BA;
output DRAM_CASN;
output DRAM_CKE;
output DRAM_CLK;
output DRAM_CSN;
output [2:0] DRAM_DM_RDQS_OUT;
output [17:0] DRAM_DQ_OUT;
output [2:0] DRAM_DQS_OUT;
output [1:0] DRAM_FIFO_WE_OUT;
output DRAM_ODT;
output DRAM_RASN;
output DRAM_RSTN;
output DRAM_WEN;
output I2C0_SCL_USBC_DATA1_MGPIO31B_OUT;
output I2C0_SDA_USBC_DATA0_MGPIO30B_OUT;
output I2C1_SCL_USBA_DATA4_MGPIO1A_OUT;
output I2C1_SDA_USBA_DATA3_MGPIO0A_OUT;
output MMUART0_CTS_USBC_DATA7_MGPIO19B_OUT;
output MMUART0_DCD_MGPIO22B_OUT;
output MMUART0_DSR_MGPIO20B_OUT;
output MMUART0_DTR_USBC_DATA6_MGPIO18B_OUT;
output MMUART0_RI_MGPIO21B_OUT;
output MMUART0_RTS_USBC_DATA5_MGPIO17B_OUT;
output MMUART0_RXD_USBC_STP_MGPIO28B_OUT;
output MMUART0_SCK_USBC_NXT_MGPIO29B_OUT;
output MMUART0_TXD_USBC_DIR_MGPIO27B_OUT;
output MMUART1_RXD_USBC_DATA3_MGPIO26B_OUT;
output MMUART1_SCK_USBC_DATA4_MGPIO25B_OUT;
output MMUART1_TXD_USBC_DATA2_MGPIO24B_OUT;
output RGMII_GTX_CLK_RMII_CLK_USBB_XCLK_OUT;
output RGMII_MDC_RMII_MDC_OUT;
output RGMII_MDIO_RMII_MDIO_USBB_DATA7_OUT;
output RGMII_RX_CLK_OUT;
output RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_OUT;
output RGMII_RXD0_RMII_RXD0_USBB_DATA0_OUT;
output RGMII_RXD1_RMII_RXD1_USBB_DATA1_OUT;
output RGMII_RXD2_RMII_RX_ER_USBB_DATA3_OUT;
output RGMII_RXD3_USBB_DATA4_OUT;
output RGMII_TX_CLK_OUT;
output RGMII_TX_CTL_RMII_TX_EN_USBB_NXT_OUT;
output RGMII_TXD0_RMII_TXD0_USBB_DIR_OUT;
output RGMII_TXD1_RMII_TXD1_USBB_STP_OUT;
output RGMII_TXD2_USBB_DATA5_OUT;
output RGMII_TXD3_USBB_DATA6_OUT;
output SPI0_SCK_USBA_XCLK_OUT;
output SPI0_SDI_USBA_DIR_MGPIO5A_OUT;
output SPI0_SDO_USBA_STP_MGPIO6A_OUT;
output SPI0_SS0_USBA_NXT_MGPIO7A_OUT;
output SPI0_SS1_USBA_DATA5_MGPIO8A_OUT;
output SPI0_SS2_USBA_DATA6_MGPIO9A_OUT;
output SPI0_SS3_USBA_DATA7_MGPIO10A_OUT;
output SPI1_SCK_OUT;
output SPI1_SDI_MGPIO11A_OUT;
output SPI1_SDO_MGPIO12A_OUT;
output SPI1_SS0_MGPIO13A_OUT;
output SPI1_SS1_MGPIO14A_OUT;
output SPI1_SS2_MGPIO15A_OUT;
output SPI1_SS3_MGPIO16A_OUT;
output SPI1_SS4_MGPIO17A_OUT;
output SPI1_SS5_MGPIO18A_OUT;
output SPI1_SS6_MGPIO23A_OUT;
output SPI1_SS7_MGPIO24A_OUT;
output USBC_XCLK_OUT;
output CAN_RXBUS_USBA_DATA1_MGPIO3A_OE;
output CAN_TX_EBL_USBA_DATA2_MGPIO4A_OE;
output CAN_TXBUS_USBA_DATA0_MGPIO2A_OE;
output [2:0] DM_OE;
output [17:0] DRAM_DQ_OE;
output [2:0] DRAM_DQS_OE;
output I2C0_SCL_USBC_DATA1_MGPIO31B_OE;
output I2C0_SDA_USBC_DATA0_MGPIO30B_OE;
output I2C1_SCL_USBA_DATA4_MGPIO1A_OE;
output I2C1_SDA_USBA_DATA3_MGPIO0A_OE;
output MMUART0_CTS_USBC_DATA7_MGPIO19B_OE;
output MMUART0_DCD_MGPIO22B_OE;
output MMUART0_DSR_MGPIO20B_OE;
output MMUART0_DTR_USBC_DATA6_MGPIO18B_OE;
output MMUART0_RI_MGPIO21B_OE;
output MMUART0_RTS_USBC_DATA5_MGPIO17B_OE;
output MMUART0_RXD_USBC_STP_MGPIO28B_OE;
output MMUART0_SCK_USBC_NXT_MGPIO29B_OE;
output MMUART0_TXD_USBC_DIR_MGPIO27B_OE;
output MMUART1_RXD_USBC_DATA3_MGPIO26B_OE;
output MMUART1_SCK_USBC_DATA4_MGPIO25B_OE;
output MMUART1_TXD_USBC_DATA2_MGPIO24B_OE;
output RGMII_GTX_CLK_RMII_CLK_USBB_XCLK_OE;
output RGMII_MDC_RMII_MDC_OE;
output RGMII_MDIO_RMII_MDIO_USBB_DATA7_OE;
output RGMII_RX_CLK_OE;
output RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_OE;
output RGMII_RXD0_RMII_RXD0_USBB_DATA0_OE;
output RGMII_RXD1_RMII_RXD1_USBB_DATA1_OE;
output RGMII_RXD2_RMII_RX_ER_USBB_DATA3_OE;
output RGMII_RXD3_USBB_DATA4_OE;
output RGMII_TX_CLK_OE;
output RGMII_TX_CTL_RMII_TX_EN_USBB_NXT_OE;
output RGMII_TXD0_RMII_TXD0_USBB_DIR_OE;
output RGMII_TXD1_RMII_TXD1_USBB_STP_OE;
output RGMII_TXD2_USBB_DATA5_OE;
output RGMII_TXD3_USBB_DATA6_OE;
output SPI0_SCK_USBA_XCLK_OE;
output SPI0_SDI_USBA_DIR_MGPIO5A_OE;
output SPI0_SDO_USBA_STP_MGPIO6A_OE;
output SPI0_SS0_USBA_NXT_MGPIO7A_OE;
output SPI0_SS1_USBA_DATA5_MGPIO8A_OE;
output SPI0_SS2_USBA_DATA6_MGPIO9A_OE;
output SPI0_SS3_USBA_DATA7_MGPIO10A_OE;
output SPI1_SCK_OE;
output SPI1_SDI_MGPIO11A_OE;
output SPI1_SDO_MGPIO12A_OE;
output SPI1_SS0_MGPIO13A_OE;
output SPI1_SS1_MGPIO14A_OE;
output SPI1_SS2_MGPIO15A_OE;
output SPI1_SS3_MGPIO16A_OE;
output SPI1_SS4_MGPIO17A_OE;
output SPI1_SS5_MGPIO18A_OE;
output SPI1_SS6_MGPIO23A_OE;
output SPI1_SS7_MGPIO24A_OE;
output USBC_XCLK_OE;

    parameter INIT = 'h0 ;
    parameter ACT_UBITS = 'hFFFFFFFFFFFFFF ;
    parameter MEMORYFILE = "" ;
    parameter RTC_MAIN_XTL_FREQ = 0.0 ;
    parameter RTC_MAIN_XTL_MODE = "1" ;
    
endmodule


module coreapb3_iaddr_reg_0s_32_28(
       IADDR_REG,
       CoreAPB3_0_APBmslave4_PWDATA,
       PRDATA_0_iv_0_0_a2_0_18,
       PRDATA_0_iv_0_0_a2_0_17,
       MSS_RESET_N_M2F_c,
       FCCC_0_GL1,
       CoreAPB3_0_APBmslave4_PENABLE,
       CoreAPB3_0_APBmslave4_PWRITE
    );
output [31:0] IADDR_REG;
input  [31:0] CoreAPB3_0_APBmslave4_PWDATA;
input  [3:3] PRDATA_0_iv_0_0_a2_0_18;
input  [3:3] PRDATA_0_iv_0_0_a2_0_17;
input  MSS_RESET_N_M2F_c;
input  FCCC_0_GL1;
input  CoreAPB3_0_APBmslave4_PENABLE;
input  CoreAPB3_0_APBmslave4_PWRITE;

    wire VCC_net_1, IADDR_REG_0_sqmuxa, GND_net_1;
    
    SLE \IADDR_REG[26]  (.D(CoreAPB3_0_APBmslave4_PWDATA[26]), .CLK(
        FCCC_0_GL1), .EN(IADDR_REG_0_sqmuxa), .ALn(MSS_RESET_N_M2F_c), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(IADDR_REG[26]));
    SLE \IADDR_REG[30]  (.D(CoreAPB3_0_APBmslave4_PWDATA[30]), .CLK(
        FCCC_0_GL1), .EN(IADDR_REG_0_sqmuxa), .ALn(MSS_RESET_N_M2F_c), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(IADDR_REG[30]));
    SLE \IADDR_REG[25]  (.D(CoreAPB3_0_APBmslave4_PWDATA[25]), .CLK(
        FCCC_0_GL1), .EN(IADDR_REG_0_sqmuxa), .ALn(MSS_RESET_N_M2F_c), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(IADDR_REG[25]));
    SLE \IADDR_REG[27]  (.D(CoreAPB3_0_APBmslave4_PWDATA[27]), .CLK(
        FCCC_0_GL1), .EN(IADDR_REG_0_sqmuxa), .ALn(MSS_RESET_N_M2F_c), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(IADDR_REG[27]));
    SLE \IADDR_REG[14]  (.D(CoreAPB3_0_APBmslave4_PWDATA[14]), .CLK(
        FCCC_0_GL1), .EN(IADDR_REG_0_sqmuxa), .ALn(MSS_RESET_N_M2F_c), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(IADDR_REG[14]));
    SLE \IADDR_REG[18]  (.D(CoreAPB3_0_APBmslave4_PWDATA[18]), .CLK(
        FCCC_0_GL1), .EN(IADDR_REG_0_sqmuxa), .ALn(MSS_RESET_N_M2F_c), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(IADDR_REG[18]));
    SLE \IADDR_REG[8]  (.D(CoreAPB3_0_APBmslave4_PWDATA[8]), .CLK(
        FCCC_0_GL1), .EN(IADDR_REG_0_sqmuxa), .ALn(MSS_RESET_N_M2F_c), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(IADDR_REG[8]));
    VCC VCC (.Y(VCC_net_1));
    SLE \IADDR_REG[7]  (.D(CoreAPB3_0_APBmslave4_PWDATA[7]), .CLK(
        FCCC_0_GL1), .EN(IADDR_REG_0_sqmuxa), .ALn(MSS_RESET_N_M2F_c), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(IADDR_REG[7]));
    SLE \IADDR_REG[29]  (.D(CoreAPB3_0_APBmslave4_PWDATA[29]), .CLK(
        FCCC_0_GL1), .EN(IADDR_REG_0_sqmuxa), .ALn(MSS_RESET_N_M2F_c), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(IADDR_REG[29]));
    SLE \IADDR_REG[5]  (.D(CoreAPB3_0_APBmslave4_PWDATA[5]), .CLK(
        FCCC_0_GL1), .EN(IADDR_REG_0_sqmuxa), .ALn(MSS_RESET_N_M2F_c), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(IADDR_REG[5]));
    SLE \IADDR_REG[20]  (.D(CoreAPB3_0_APBmslave4_PWDATA[20]), .CLK(
        FCCC_0_GL1), .EN(IADDR_REG_0_sqmuxa), .ALn(MSS_RESET_N_M2F_c), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(IADDR_REG[20]));
    SLE \IADDR_REG[4]  (.D(CoreAPB3_0_APBmslave4_PWDATA[4]), .CLK(
        FCCC_0_GL1), .EN(IADDR_REG_0_sqmuxa), .ALn(MSS_RESET_N_M2F_c), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(IADDR_REG[4]));
    CFG4 #( .INIT(16'h8000) )  IADDR_REG_0_sqmuxa_0_a3_0_a3 (.A(
        CoreAPB3_0_APBmslave4_PENABLE), .B(
        CoreAPB3_0_APBmslave4_PWRITE), .C(PRDATA_0_iv_0_0_a2_0_18[3]), 
        .D(PRDATA_0_iv_0_0_a2_0_17[3]), .Y(IADDR_REG_0_sqmuxa));
    SLE \IADDR_REG[31]  (.D(CoreAPB3_0_APBmslave4_PWDATA[31]), .CLK(
        FCCC_0_GL1), .EN(IADDR_REG_0_sqmuxa), .ALn(MSS_RESET_N_M2F_c), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(IADDR_REG[31]));
    SLE \IADDR_REG[2]  (.D(CoreAPB3_0_APBmslave4_PWDATA[2]), .CLK(
        FCCC_0_GL1), .EN(IADDR_REG_0_sqmuxa), .ALn(MSS_RESET_N_M2F_c), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(IADDR_REG[2]));
    SLE \IADDR_REG[23]  (.D(CoreAPB3_0_APBmslave4_PWDATA[23]), .CLK(
        FCCC_0_GL1), .EN(IADDR_REG_0_sqmuxa), .ALn(MSS_RESET_N_M2F_c), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(IADDR_REG[23]));
    GND GND (.Y(GND_net_1));
    SLE \IADDR_REG[22]  (.D(CoreAPB3_0_APBmslave4_PWDATA[22]), .CLK(
        FCCC_0_GL1), .EN(IADDR_REG_0_sqmuxa), .ALn(MSS_RESET_N_M2F_c), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(IADDR_REG[22]));
    SLE \IADDR_REG[16]  (.D(CoreAPB3_0_APBmslave4_PWDATA[16]), .CLK(
        FCCC_0_GL1), .EN(IADDR_REG_0_sqmuxa), .ALn(MSS_RESET_N_M2F_c), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(IADDR_REG[16]));
    SLE \IADDR_REG[15]  (.D(CoreAPB3_0_APBmslave4_PWDATA[15]), .CLK(
        FCCC_0_GL1), .EN(IADDR_REG_0_sqmuxa), .ALn(MSS_RESET_N_M2F_c), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(IADDR_REG[15]));
    SLE \IADDR_REG[1]  (.D(CoreAPB3_0_APBmslave4_PWDATA[1]), .CLK(
        FCCC_0_GL1), .EN(IADDR_REG_0_sqmuxa), .ALn(MSS_RESET_N_M2F_c), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(IADDR_REG[1]));
    SLE \IADDR_REG[3]  (.D(CoreAPB3_0_APBmslave4_PWDATA[3]), .CLK(
        FCCC_0_GL1), .EN(IADDR_REG_0_sqmuxa), .ALn(MSS_RESET_N_M2F_c), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(IADDR_REG[3]));
    SLE \IADDR_REG[17]  (.D(CoreAPB3_0_APBmslave4_PWDATA[17]), .CLK(
        FCCC_0_GL1), .EN(IADDR_REG_0_sqmuxa), .ALn(MSS_RESET_N_M2F_c), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(IADDR_REG[17]));
    SLE \IADDR_REG[21]  (.D(CoreAPB3_0_APBmslave4_PWDATA[21]), .CLK(
        FCCC_0_GL1), .EN(IADDR_REG_0_sqmuxa), .ALn(MSS_RESET_N_M2F_c), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(IADDR_REG[21]));
    SLE \IADDR_REG[6]  (.D(CoreAPB3_0_APBmslave4_PWDATA[6]), .CLK(
        FCCC_0_GL1), .EN(IADDR_REG_0_sqmuxa), .ALn(MSS_RESET_N_M2F_c), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(IADDR_REG[6]));
    SLE \IADDR_REG[0]  (.D(CoreAPB3_0_APBmslave4_PWDATA[0]), .CLK(
        FCCC_0_GL1), .EN(IADDR_REG_0_sqmuxa), .ALn(MSS_RESET_N_M2F_c), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(IADDR_REG[0]));
    SLE \IADDR_REG[19]  (.D(CoreAPB3_0_APBmslave4_PWDATA[19]), .CLK(
        FCCC_0_GL1), .EN(IADDR_REG_0_sqmuxa), .ALn(MSS_RESET_N_M2F_c), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(IADDR_REG[19]));
    SLE \IADDR_REG[10]  (.D(CoreAPB3_0_APBmslave4_PWDATA[10]), .CLK(
        FCCC_0_GL1), .EN(IADDR_REG_0_sqmuxa), .ALn(MSS_RESET_N_M2F_c), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(IADDR_REG[10]));
    SLE \IADDR_REG[24]  (.D(CoreAPB3_0_APBmslave4_PWDATA[24]), .CLK(
        FCCC_0_GL1), .EN(IADDR_REG_0_sqmuxa), .ALn(MSS_RESET_N_M2F_c), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(IADDR_REG[24]));
    SLE \IADDR_REG[28]  (.D(CoreAPB3_0_APBmslave4_PWDATA[28]), .CLK(
        FCCC_0_GL1), .EN(IADDR_REG_0_sqmuxa), .ALn(MSS_RESET_N_M2F_c), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(IADDR_REG[28]));
    SLE \IADDR_REG[13]  (.D(CoreAPB3_0_APBmslave4_PWDATA[13]), .CLK(
        FCCC_0_GL1), .EN(IADDR_REG_0_sqmuxa), .ALn(MSS_RESET_N_M2F_c), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(IADDR_REG[13]));
    SLE \IADDR_REG[12]  (.D(CoreAPB3_0_APBmslave4_PWDATA[12]), .CLK(
        FCCC_0_GL1), .EN(IADDR_REG_0_sqmuxa), .ALn(MSS_RESET_N_M2F_c), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(IADDR_REG[12]));
    SLE \IADDR_REG[9]  (.D(CoreAPB3_0_APBmslave4_PWDATA[9]), .CLK(
        FCCC_0_GL1), .EN(IADDR_REG_0_sqmuxa), .ALn(MSS_RESET_N_M2F_c), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(IADDR_REG[9]));
    SLE \IADDR_REG[11]  (.D(CoreAPB3_0_APBmslave4_PWDATA[11]), .CLK(
        FCCC_0_GL1), .EN(IADDR_REG_0_sqmuxa), .ALn(MSS_RESET_N_M2F_c), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(IADDR_REG[11]));
    
endmodule


module COREAPB3_MUXPTOB3(
       PRDATA_0_iv_0_0_a2_1,
       PRDATA_0_iv_0_0_a2_0_17,
       PRDATA_0_iv_0_0_a2_0_18,
       hello_regs_MSS_0_FIC_0_APB_MASTER_PADDR,
       mem_8__2_i_0_0_a2,
       mem_0__2_i_0_0_a2,
       PRDATA_0_iv_0_0_a2_2_4,
       CoreAPB3_0_APBmslave5_PRDATA,
       PRDATA_reg,
       lsram_width32_PRDATA,
       GPIO_OUT_1_c,
       IADDR_REG,
       hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA,
       CoreAPB3_0_APBmslave4_PADDR_8,
       CoreAPB3_0_APBmslave4_PADDR_7,
       CoreAPB3_0_APBmslave4_PADDR_0,
       CoreAPB3_0_APBmslave4_PADDR_6,
       CoreAPB3_0_APBmslave4_PADDR_1,
       hello_regs_MSS_0_FIC_0_APB_MASTER_PSELx,
       N_928,
       CoreAPB3_0_APBmslave4_PWRITE,
       CoreAPB3_0_APBmslave4_PENABLE,
       PRDATA4,
       CoreAPB3_0_APBmslave4_PREADY,
       N_676_i_0
    );
output [3:3] PRDATA_0_iv_0_0_a2_1;
output [3:3] PRDATA_0_iv_0_0_a2_0_17;
output [3:3] PRDATA_0_iv_0_0_a2_0_18;
input  [27:9] hello_regs_MSS_0_FIC_0_APB_MASTER_PADDR;
input  [2:2] mem_8__2_i_0_0_a2;
input  [0:0] mem_0__2_i_0_0_a2;
output [3:3] PRDATA_0_iv_0_0_a2_2_4;
input  [7:0] CoreAPB3_0_APBmslave5_PRDATA;
input  [31:0] PRDATA_reg;
input  [31:0] lsram_width32_PRDATA;
input  [7:0] GPIO_OUT_1_c;
input  [31:0] IADDR_REG;
output [31:0] hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA;
input  CoreAPB3_0_APBmslave4_PADDR_8;
input  CoreAPB3_0_APBmslave4_PADDR_7;
input  CoreAPB3_0_APBmslave4_PADDR_0;
input  CoreAPB3_0_APBmslave4_PADDR_6;
input  CoreAPB3_0_APBmslave4_PADDR_1;
input  hello_regs_MSS_0_FIC_0_APB_MASTER_PSELx;
input  N_928;
input  CoreAPB3_0_APBmslave4_PWRITE;
input  CoreAPB3_0_APBmslave4_PENABLE;
input  PRDATA4;
input  CoreAPB3_0_APBmslave4_PREADY;
output N_676_i_0;

    wire \PRDATA_0_iv_0_0_a2_1_1[3]_net_1 , 
        \PRDATA_0_iv_0_0_0[3]_net_1 , \PRDATA_0_iv_0_0_1[3]_net_1 , 
        \PRDATA_0_iv_0_0_a3[3]_net_1 , 
        \PRDATA_0_iv_0_0_a2_0_18_1[3]_net_1 , 
        \PRDATA_0_iv_0_0_a2_0_18_8[3]_net_1 , 
        \PRDATA_0_iv_0_0_a2_0_18_9[3]_net_1 , 
        \PRDATA_0_iv_0_0_a2_0_18_7[3]_net_1 , 
        \PRDATA_0_iv_0_0_a2[3]_net_1 , \PRDATA_0_iv_0_0_a3_0[3] , 
        \PRDATA_0_iv_0_0_a2_0_17_2[3]_net_1 , 
        \PRDATA_0_iv_0_0_a2_2_4_2[3]_net_1 , N_688, 
        \PRDATA_0_iv_0_0_a3_2_0[3]_net_1 , 
        \PRDATA_0_iv_0_0_a3_0[2]_net_1 , 
        \PRDATA_0_iv_0_0_a3_0[1]_net_1 , 
        \PRDATA_0_iv_0_0_a3_0[0]_net_1 , 
        \PRDATA_0_iv_0_0_a3_0[7]_net_1 , 
        \PRDATA_0_iv_0_0_a3_0[6]_net_1 , 
        \PRDATA_0_iv_0_0_a3_0[5]_net_1 , 
        \PRDATA_0_iv_0_0_a3_0[4]_net_1 , \PRDATA_0_iv_0_0_1[1]_net_1 , 
        \PRDATA_0_iv_0_0_1[0]_net_1 , \PRDATA_0_iv_0_0_1[7]_net_1 , 
        \PRDATA_0_iv_0_0_1[2]_net_1 , \PRDATA_0_iv_0_0_1[5]_net_1 , 
        \PRDATA_0_iv_0_0_1[4]_net_1 , \PRDATA_0_iv_0_0_1[6]_net_1 , 
        \PRDATA_0_iv_0_0_0[10]_net_1 , \PRDATA_0_iv_0_0_0[18]_net_1 , 
        \PRDATA_0_iv_0_0_0[31]_net_1 , \PRDATA_0_iv_0_0_0[12]_net_1 , 
        \PRDATA_0_iv_0_0_0[26]_net_1 , \PRDATA_0_iv_0_0_0[25]_net_1 , 
        \PRDATA_0_iv_0_0_0[16]_net_1 , \PRDATA_0_iv_0_0_0[15]_net_1 , 
        \PRDATA_0_iv_0_0_0[17]_net_1 , \PRDATA_0_iv_0_0_0[19]_net_1 , 
        \PRDATA_0_iv_0_0_0[29]_net_1 , \PRDATA_0_iv_0_0_0[30]_net_1 , 
        \PRDATA_0_iv_0_0_0[8]_net_1 , \PRDATA_0_iv_0_0_0[11]_net_1 , 
        \PRDATA_0_iv_0_0_0[21]_net_1 , \PRDATA_0_iv_0_0_0[14]_net_1 , 
        \PRDATA_0_iv_0_0_0[27]_net_1 , \PRDATA_0_iv_0_0_0[28]_net_1 , 
        \PRDATA_0_iv_0_0_0[20]_net_1 , \PRDATA_0_iv_0_0_0[22]_net_1 , 
        \PRDATA_0_iv_0_0_0[13]_net_1 , \PRDATA_0_iv_0_0_0[9]_net_1 , 
        \PRDATA_0_iv_0_0_0[24]_net_1 , \PRDATA_0_iv_0_0_0[23]_net_1 , 
        \PRDATA_0_iv_0_0_a3_3_0[5]_net_1 , 
        \PRDATA_0_iv_0_0_a3_3_0[1]_net_1 , 
        \PRDATA_0_iv_0_0_a3_3_0[6]_net_1 , 
        \PRDATA_0_iv_0_0_a3_3_0[0]_net_1 , 
        \PRDATA_0_iv_0_0_a3_3_0[4]_net_1 , 
        \PRDATA_0_iv_0_0_a3_3_0[2]_net_1 , 
        \PRDATA_0_iv_0_0_a3_1_0[9]_net_1 , 
        \PRDATA_0_iv_0_0_a3_3_0[7]_net_1 , 
        \PRDATA_0_iv_0_0_a3_1_0[23]_net_1 , 
        \PRDATA_0_iv_0_0_0[1]_net_1 , \PRDATA_0_iv_0_0_0[0]_net_1 , 
        \PRDATA_0_iv_0_0_0[7]_net_1 , \PRDATA_0_iv_0_0_0[2]_net_1 , 
        \PRDATA_0_iv_0_0_0[5]_net_1 , \PRDATA_0_iv_0_0_0[4]_net_1 , 
        \PRDATA_0_iv_0_0_0[6]_net_1 , GND_net_1, VCC_net_1;
    
    CFG4 #( .INIT(16'hECA0) )  \PRDATA_0_iv_0_0_0[29]  (.A(
        \PRDATA_0_iv_0_0_a2[3]_net_1 ), .B(PRDATA4), .C(PRDATA_reg[29])
        , .D(lsram_width32_PRDATA[29]), .Y(
        \PRDATA_0_iv_0_0_0[29]_net_1 ));
    CFG4 #( .INIT(16'hECA0) )  \PRDATA_0_iv_0_0_0[10]  (.A(
        \PRDATA_0_iv_0_0_a2[3]_net_1 ), .B(PRDATA4), .C(PRDATA_reg[10])
        , .D(lsram_width32_PRDATA[10]), .Y(
        \PRDATA_0_iv_0_0_0[10]_net_1 ));
    CFG4 #( .INIT(16'hFF80) )  \PRDATA_0_iv_0_0_0[2]  (.A(
        mem_8__2_i_0_0_a2[2]), .B(GPIO_OUT_1_c[2]), .C(
        PRDATA_0_iv_0_0_a2_2_4[3]), .D(\PRDATA_0_iv_0_0_a3_0[2]_net_1 )
        , .Y(\PRDATA_0_iv_0_0_0[2]_net_1 ));
    CFG4 #( .INIT(16'hECA0) )  \PRDATA_0_iv_0_0_0[24]  (.A(
        \PRDATA_0_iv_0_0_a2[3]_net_1 ), .B(PRDATA4), .C(PRDATA_reg[24])
        , .D(lsram_width32_PRDATA[24]), .Y(
        \PRDATA_0_iv_0_0_0[24]_net_1 ));
    CFG4 #( .INIT(16'hECA0) )  \PRDATA_0_iv_0_0_0[22]  (.A(
        \PRDATA_0_iv_0_0_a2[3]_net_1 ), .B(PRDATA4), .C(PRDATA_reg[22])
        , .D(lsram_width32_PRDATA[22]), .Y(
        \PRDATA_0_iv_0_0_0[22]_net_1 ));
    CFG4 #( .INIT(16'h8000) )  \PRDATA_0_iv_0_0_a3_3_0[0]  (.A(N_688), 
        .B(IADDR_REG[0]), .C(\PRDATA_0_iv_0_0_a2_0_17_2[3]_net_1 ), .D(
        mem_0__2_i_0_0_a2[0]), .Y(\PRDATA_0_iv_0_0_a3_3_0[0]_net_1 ));
    CFG3 #( .INIT(8'hDF) )  N_676_i (.A(N_928), .B(
        CoreAPB3_0_APBmslave4_PREADY), .C(
        hello_regs_MSS_0_FIC_0_APB_MASTER_PADDR[26]), .Y(N_676_i_0));
    CFG4 #( .INIT(16'hECA0) )  \PRDATA_0_iv_0_0_0[31]  (.A(
        \PRDATA_0_iv_0_0_a2[3]_net_1 ), .B(PRDATA4), .C(PRDATA_reg[31])
        , .D(lsram_width32_PRDATA[31]), .Y(
        \PRDATA_0_iv_0_0_0[31]_net_1 ));
    CFG3 #( .INIT(8'hC4) )  \PRDATA_0_iv_0_0_a3_0_0[3]  (.A(
        CoreAPB3_0_APBmslave4_PENABLE), .B(PRDATA_reg[3]), .C(
        CoreAPB3_0_APBmslave4_PWRITE), .Y(\PRDATA_0_iv_0_0_a3_0[3] ));
    CFG4 #( .INIT(16'hECA0) )  \PRDATA_0_iv_0_0_0[18]  (.A(
        \PRDATA_0_iv_0_0_a2[3]_net_1 ), .B(PRDATA4), .C(PRDATA_reg[18])
        , .D(lsram_width32_PRDATA[18]), .Y(
        \PRDATA_0_iv_0_0_0[18]_net_1 ));
    CFG3 #( .INIT(8'hF8) )  \PRDATA_0_iv_0_0[9]  (.A(
        \PRDATA_0_iv_0_0_a3_1_0[9]_net_1 ), .B(
        PRDATA_0_iv_0_0_a2_0_18[3]), .C(\PRDATA_0_iv_0_0_0[9]_net_1 ), 
        .Y(hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[9]));
    CFG4 #( .INIT(16'hFFF8) )  \PRDATA_0_iv_0_0[4]  (.A(
        PRDATA_0_iv_0_0_a2_0_18[3]), .B(
        \PRDATA_0_iv_0_0_a3_3_0[4]_net_1 ), .C(
        \PRDATA_0_iv_0_0_1[4]_net_1 ), .D(\PRDATA_0_iv_0_0_0[4]_net_1 )
        , .Y(hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[4]));
    CFG4 #( .INIT(16'hF8F0) )  \PRDATA_0_iv_0_0[10]  (.A(
        PRDATA_0_iv_0_0_a2_0_17[3]), .B(IADDR_REG[10]), .C(
        \PRDATA_0_iv_0_0_0[10]_net_1 ), .D(PRDATA_0_iv_0_0_a2_0_18[3]), 
        .Y(hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[10]));
    CFG2 #( .INIT(4'h8) )  \PRDATA_0_iv_0_0_a3_2_0[3]  (.A(
        mem_8__2_i_0_0_a2[2]), .B(GPIO_OUT_1_c[3]), .Y(
        \PRDATA_0_iv_0_0_a3_2_0[3]_net_1 ));
    CFG4 #( .INIT(16'hECA0) )  \PRDATA_0_iv_0_0_0[9]  (.A(
        \PRDATA_0_iv_0_0_a2[3]_net_1 ), .B(PRDATA4), .C(PRDATA_reg[9]), 
        .D(lsram_width32_PRDATA[9]), .Y(\PRDATA_0_iv_0_0_0[9]_net_1 ));
    CFG4 #( .INIT(16'hF8F0) )  \PRDATA_0_iv_0_0[31]  (.A(
        PRDATA_0_iv_0_0_a2_0_17[3]), .B(IADDR_REG[31]), .C(
        \PRDATA_0_iv_0_0_0[31]_net_1 ), .D(PRDATA_0_iv_0_0_a2_0_18[3]), 
        .Y(hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[31]));
    CFG3 #( .INIT(8'h80) )  \PRDATA_0_iv_0_0_a3[3]  (.A(N_928), .B(
        hello_regs_MSS_0_FIC_0_APB_MASTER_PADDR[26]), .C(
        \PRDATA_0_iv_0_0_a3_0[3] ), .Y(\PRDATA_0_iv_0_0_a3[3]_net_1 ));
    VCC VCC (.Y(VCC_net_1));
    CFG4 #( .INIT(16'hECA0) )  \PRDATA_0_iv_0_0_0[21]  (.A(
        \PRDATA_0_iv_0_0_a2[3]_net_1 ), .B(PRDATA4), .C(PRDATA_reg[21])
        , .D(lsram_width32_PRDATA[21]), .Y(
        \PRDATA_0_iv_0_0_0[21]_net_1 ));
    CFG4 #( .INIT(16'hF8F0) )  \PRDATA_0_iv_0_0[8]  (.A(
        PRDATA_0_iv_0_0_a2_0_17[3]), .B(IADDR_REG[8]), .C(
        \PRDATA_0_iv_0_0_0[8]_net_1 ), .D(PRDATA_0_iv_0_0_a2_0_18[3]), 
        .Y(hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[8]));
    CFG4 #( .INIT(16'hECA0) )  \PRDATA_0_iv_0_0_0[8]  (.A(
        \PRDATA_0_iv_0_0_a2[3]_net_1 ), .B(PRDATA4), .C(PRDATA_reg[8]), 
        .D(lsram_width32_PRDATA[8]), .Y(\PRDATA_0_iv_0_0_0[8]_net_1 ));
    CFG4 #( .INIT(16'hFF80) )  \PRDATA_0_iv_0_0_0[7]  (.A(
        mem_8__2_i_0_0_a2[2]), .B(GPIO_OUT_1_c[7]), .C(
        PRDATA_0_iv_0_0_a2_2_4[3]), .D(\PRDATA_0_iv_0_0_a3_0[7]_net_1 )
        , .Y(\PRDATA_0_iv_0_0_0[7]_net_1 ));
    CFG4 #( .INIT(16'h4000) )  \PRDATA_0_iv_0_0_a2_1[3]  (.A(
        hello_regs_MSS_0_FIC_0_APB_MASTER_PADDR[27]), .B(
        hello_regs_MSS_0_FIC_0_APB_MASTER_PADDR[24]), .C(
        \PRDATA_0_iv_0_0_a2_1_1[3]_net_1 ), .D(
        hello_regs_MSS_0_FIC_0_APB_MASTER_PADDR[26]), .Y(
        PRDATA_0_iv_0_0_a2_1[3]));
    CFG4 #( .INIT(16'hECA0) )  \PRDATA_0_iv_0_0_0[30]  (.A(
        \PRDATA_0_iv_0_0_a2[3]_net_1 ), .B(PRDATA4), .C(PRDATA_reg[30])
        , .D(lsram_width32_PRDATA[30]), .Y(
        \PRDATA_0_iv_0_0_0[30]_net_1 ));
    CFG4 #( .INIT(16'hF8F0) )  \PRDATA_0_iv_0_0[20]  (.A(
        PRDATA_0_iv_0_0_a2_0_17[3]), .B(IADDR_REG[20]), .C(
        \PRDATA_0_iv_0_0_0[20]_net_1 ), .D(PRDATA_0_iv_0_0_a2_0_18[3]), 
        .Y(hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[20]));
    CFG4 #( .INIT(16'h8000) )  \PRDATA_0_iv_0_0_a3_3_0[4]  (.A(N_688), 
        .B(IADDR_REG[4]), .C(\PRDATA_0_iv_0_0_a2_0_17_2[3]_net_1 ), .D(
        mem_0__2_i_0_0_a2[0]), .Y(\PRDATA_0_iv_0_0_a3_3_0[4]_net_1 ));
    CFG4 #( .INIT(16'hECA0) )  \PRDATA_0_iv_0_0_1[5]  (.A(
        \PRDATA_0_iv_0_0_a2[3]_net_1 ), .B(PRDATA4), .C(PRDATA_reg[5]), 
        .D(lsram_width32_PRDATA[5]), .Y(\PRDATA_0_iv_0_0_1[5]_net_1 ));
    CFG4 #( .INIT(16'hECA0) )  \PRDATA_0_iv_0_0_0[27]  (.A(
        \PRDATA_0_iv_0_0_a2[3]_net_1 ), .B(PRDATA4), .C(PRDATA_reg[27])
        , .D(lsram_width32_PRDATA[27]), .Y(
        \PRDATA_0_iv_0_0_0[27]_net_1 ));
    CFG2 #( .INIT(4'h4) )  \PRDATA_0_iv_0_0_a2_1_1[3]  (.A(
        hello_regs_MSS_0_FIC_0_APB_MASTER_PADDR[25]), .B(
        hello_regs_MSS_0_FIC_0_APB_MASTER_PSELx), .Y(
        \PRDATA_0_iv_0_0_a2_1_1[3]_net_1 ));
    CFG4 #( .INIT(16'hFFF8) )  \PRDATA_0_iv_0_0[2]  (.A(
        PRDATA_0_iv_0_0_a2_0_18[3]), .B(
        \PRDATA_0_iv_0_0_a3_3_0[2]_net_1 ), .C(
        \PRDATA_0_iv_0_0_1[2]_net_1 ), .D(\PRDATA_0_iv_0_0_0[2]_net_1 )
        , .Y(hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[2]));
    CFG3 #( .INIT(8'h80) )  \PRDATA_0_iv_0_0_a2_0_17[3]  (.A(
        mem_0__2_i_0_0_a2[0]), .B(\PRDATA_0_iv_0_0_a2_0_17_2[3]_net_1 )
        , .C(N_688), .Y(PRDATA_0_iv_0_0_a2_0_17[3]));
    CFG4 #( .INIT(16'hF8F0) )  \PRDATA_0_iv_0_0[13]  (.A(
        PRDATA_0_iv_0_0_a2_0_17[3]), .B(IADDR_REG[13]), .C(
        \PRDATA_0_iv_0_0_0[13]_net_1 ), .D(PRDATA_0_iv_0_0_a2_0_18[3]), 
        .Y(hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[13]));
    CFG4 #( .INIT(16'hF8F0) )  \PRDATA_0_iv_0_0[19]  (.A(
        PRDATA_0_iv_0_0_a2_0_17[3]), .B(IADDR_REG[19]), .C(
        \PRDATA_0_iv_0_0_0[19]_net_1 ), .D(PRDATA_0_iv_0_0_a2_0_18[3]), 
        .Y(hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[19]));
    CFG2 #( .INIT(4'h8) )  \PRDATA_0_iv_0_0_a3_0[4]  (.A(
        PRDATA_0_iv_0_0_a2_1[3]), .B(CoreAPB3_0_APBmslave5_PRDATA[4]), 
        .Y(\PRDATA_0_iv_0_0_a3_0[4]_net_1 ));
    CFG4 #( .INIT(16'hEAC0) )  \PRDATA_0_iv_0_0_1[3]  (.A(
        \PRDATA_0_iv_0_0_a3_2_0[3]_net_1 ), .B(lsram_width32_PRDATA[3])
        , .C(PRDATA4), .D(PRDATA_0_iv_0_0_a2_2_4[3]), .Y(
        \PRDATA_0_iv_0_0_1[3]_net_1 ));
    CFG4 #( .INIT(16'hECA0) )  \PRDATA_0_iv_0_0_0[26]  (.A(
        \PRDATA_0_iv_0_0_a2[3]_net_1 ), .B(PRDATA4), .C(PRDATA_reg[26])
        , .D(lsram_width32_PRDATA[26]), .Y(
        \PRDATA_0_iv_0_0_0[26]_net_1 ));
    CFG2 #( .INIT(4'h8) )  \PRDATA_0_iv_0_0_a3_0[1]  (.A(
        PRDATA_0_iv_0_0_a2_1[3]), .B(CoreAPB3_0_APBmslave5_PRDATA[1]), 
        .Y(\PRDATA_0_iv_0_0_a3_0[1]_net_1 ));
    CFG3 #( .INIT(8'h01) )  \PRDATA_0_iv_0_a2_2[3]  (.A(
        CoreAPB3_0_APBmslave4_PADDR_0), .B(
        CoreAPB3_0_APBmslave4_PADDR_6), .C(
        CoreAPB3_0_APBmslave4_PADDR_1), .Y(N_688));
    CFG4 #( .INIT(16'h8000) )  \PRDATA_0_iv_0_0_a3_3_0[5]  (.A(N_688), 
        .B(IADDR_REG[5]), .C(\PRDATA_0_iv_0_0_a2_0_17_2[3]_net_1 ), .D(
        mem_0__2_i_0_0_a2[0]), .Y(\PRDATA_0_iv_0_0_a3_3_0[5]_net_1 ));
    CFG4 #( .INIT(16'hECA0) )  \PRDATA_0_iv_0_0_1[1]  (.A(
        \PRDATA_0_iv_0_0_a2[3]_net_1 ), .B(PRDATA4), .C(PRDATA_reg[1]), 
        .D(lsram_width32_PRDATA[1]), .Y(\PRDATA_0_iv_0_0_1[1]_net_1 ));
    CFG4 #( .INIT(16'hB000) )  \PRDATA_0_iv_0_0_a2[3]  (.A(
        CoreAPB3_0_APBmslave4_PWRITE), .B(
        CoreAPB3_0_APBmslave4_PENABLE), .C(
        hello_regs_MSS_0_FIC_0_APB_MASTER_PADDR[26]), .D(N_928), .Y(
        \PRDATA_0_iv_0_0_a2[3]_net_1 ));
    CFG4 #( .INIT(16'hF8F0) )  \PRDATA_0_iv_0_0[15]  (.A(
        PRDATA_0_iv_0_0_a2_0_17[3]), .B(IADDR_REG[15]), .C(
        \PRDATA_0_iv_0_0_0[15]_net_1 ), .D(PRDATA_0_iv_0_0_a2_0_18[3]), 
        .Y(hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[15]));
    CFG4 #( .INIT(16'hFF80) )  \PRDATA_0_iv_0_0_0[1]  (.A(
        mem_8__2_i_0_0_a2[2]), .B(GPIO_OUT_1_c[1]), .C(
        PRDATA_0_iv_0_0_a2_2_4[3]), .D(\PRDATA_0_iv_0_0_a3_0[1]_net_1 )
        , .Y(\PRDATA_0_iv_0_0_0[1]_net_1 ));
    CFG4 #( .INIT(16'hFFF8) )  \PRDATA_0_iv_0_0[6]  (.A(
        PRDATA_0_iv_0_0_a2_0_18[3]), .B(
        \PRDATA_0_iv_0_0_a3_3_0[6]_net_1 ), .C(
        \PRDATA_0_iv_0_0_1[6]_net_1 ), .D(\PRDATA_0_iv_0_0_0[6]_net_1 )
        , .Y(hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[6]));
    CFG2 #( .INIT(4'h8) )  \PRDATA_0_iv_0_0_a3_0[0]  (.A(
        PRDATA_0_iv_0_0_a2_1[3]), .B(CoreAPB3_0_APBmslave5_PRDATA[0]), 
        .Y(\PRDATA_0_iv_0_0_a3_0[0]_net_1 ));
    CFG4 #( .INIT(16'hECA0) )  \PRDATA_0_iv_0_0_0[25]  (.A(
        \PRDATA_0_iv_0_0_a2[3]_net_1 ), .B(PRDATA4), .C(PRDATA_reg[25])
        , .D(lsram_width32_PRDATA[25]), .Y(
        \PRDATA_0_iv_0_0_0[25]_net_1 ));
    CFG4 #( .INIT(16'hECA0) )  \PRDATA_0_iv_0_0_0[13]  (.A(
        \PRDATA_0_iv_0_0_a2[3]_net_1 ), .B(PRDATA4), .C(PRDATA_reg[13])
        , .D(lsram_width32_PRDATA[13]), .Y(
        \PRDATA_0_iv_0_0_0[13]_net_1 ));
    CFG4 #( .INIT(16'hECA0) )  \PRDATA_0_iv_0_0_0[20]  (.A(
        \PRDATA_0_iv_0_0_a2[3]_net_1 ), .B(PRDATA4), .C(PRDATA_reg[20])
        , .D(lsram_width32_PRDATA[20]), .Y(
        \PRDATA_0_iv_0_0_0[20]_net_1 ));
    CFG3 #( .INIT(8'hF8) )  \PRDATA_0_iv_0_0[23]  (.A(
        \PRDATA_0_iv_0_0_a3_1_0[23]_net_1 ), .B(
        PRDATA_0_iv_0_0_a2_0_18[3]), .C(\PRDATA_0_iv_0_0_0[23]_net_1 ), 
        .Y(hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[23]));
    CFG4 #( .INIT(16'hF8F0) )  \PRDATA_0_iv_0_0[14]  (.A(
        PRDATA_0_iv_0_0_a2_0_17[3]), .B(IADDR_REG[14]), .C(
        \PRDATA_0_iv_0_0_0[14]_net_1 ), .D(PRDATA_0_iv_0_0_a2_0_18[3]), 
        .Y(hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[14]));
    CFG4 #( .INIT(16'hF8F0) )  \PRDATA_0_iv_0_0[29]  (.A(
        PRDATA_0_iv_0_0_a2_0_17[3]), .B(IADDR_REG[29]), .C(
        \PRDATA_0_iv_0_0_0[29]_net_1 ), .D(PRDATA_0_iv_0_0_a2_0_18[3]), 
        .Y(hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[29]));
    GND GND (.Y(GND_net_1));
    CFG4 #( .INIT(16'h0001) )  \PRDATA_0_iv_0_0_a2_0_18_8[3]  (.A(
        hello_regs_MSS_0_FIC_0_APB_MASTER_PADDR[20]), .B(
        hello_regs_MSS_0_FIC_0_APB_MASTER_PADDR[13]), .C(
        hello_regs_MSS_0_FIC_0_APB_MASTER_PADDR[14]), .D(
        hello_regs_MSS_0_FIC_0_APB_MASTER_PADDR[12]), .Y(
        \PRDATA_0_iv_0_0_a2_0_18_8[3]_net_1 ));
    CFG4 #( .INIT(16'hF8F0) )  \PRDATA_0_iv_0_0[25]  (.A(
        PRDATA_0_iv_0_0_a2_0_17[3]), .B(IADDR_REG[25]), .C(
        \PRDATA_0_iv_0_0_0[25]_net_1 ), .D(PRDATA_0_iv_0_0_a2_0_18[3]), 
        .Y(hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[25]));
    CFG4 #( .INIT(16'hECA0) )  \PRDATA_0_iv_0_0_0[28]  (.A(
        \PRDATA_0_iv_0_0_a2[3]_net_1 ), .B(PRDATA4), .C(PRDATA_reg[28])
        , .D(lsram_width32_PRDATA[28]), .Y(
        \PRDATA_0_iv_0_0_0[28]_net_1 ));
    CFG4 #( .INIT(16'hECA0) )  \PRDATA_0_iv_0_0_1[6]  (.A(
        \PRDATA_0_iv_0_0_a2[3]_net_1 ), .B(PRDATA4), .C(PRDATA_reg[6]), 
        .D(lsram_width32_PRDATA[6]), .Y(\PRDATA_0_iv_0_0_1[6]_net_1 ));
    CFG4 #( .INIT(16'h4000) )  \PRDATA_0_iv_0_0_a2_2_4[3]  (.A(
        hello_regs_MSS_0_FIC_0_APB_MASTER_PADDR[27]), .B(
        hello_regs_MSS_0_FIC_0_APB_MASTER_PSELx), .C(N_688), .D(
        \PRDATA_0_iv_0_0_a2_2_4_2[3]_net_1 ), .Y(
        PRDATA_0_iv_0_0_a2_2_4[3]));
    CFG4 #( .INIT(16'hF8F0) )  \PRDATA_0_iv_0_0[18]  (.A(
        PRDATA_0_iv_0_0_a2_0_17[3]), .B(IADDR_REG[18]), .C(
        \PRDATA_0_iv_0_0_0[18]_net_1 ), .D(PRDATA_0_iv_0_0_a2_0_18[3]), 
        .Y(hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[18]));
    CFG4 #( .INIT(16'hFFF8) )  \PRDATA_0_iv_0_0[0]  (.A(
        PRDATA_0_iv_0_0_a2_0_18[3]), .B(
        \PRDATA_0_iv_0_0_a3_3_0[0]_net_1 ), .C(
        \PRDATA_0_iv_0_0_1[0]_net_1 ), .D(\PRDATA_0_iv_0_0_0[0]_net_1 )
        , .Y(hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[0]));
    CFG4 #( .INIT(16'hECA0) )  \PRDATA_0_iv_0_0_0[19]  (.A(
        \PRDATA_0_iv_0_0_a2[3]_net_1 ), .B(PRDATA4), .C(PRDATA_reg[19])
        , .D(lsram_width32_PRDATA[19]), .Y(
        \PRDATA_0_iv_0_0_0[19]_net_1 ));
    CFG4 #( .INIT(16'hF8F0) )  \PRDATA_0_iv_0_0[24]  (.A(
        PRDATA_0_iv_0_0_a2_0_17[3]), .B(IADDR_REG[24]), .C(
        \PRDATA_0_iv_0_0_0[24]_net_1 ), .D(PRDATA_0_iv_0_0_a2_0_18[3]), 
        .Y(hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[24]));
    CFG4 #( .INIT(16'hFFF8) )  \PRDATA_0_iv_0_0[1]  (.A(
        PRDATA_0_iv_0_0_a2_0_18[3]), .B(
        \PRDATA_0_iv_0_0_a3_3_0[1]_net_1 ), .C(
        \PRDATA_0_iv_0_0_1[1]_net_1 ), .D(\PRDATA_0_iv_0_0_0[1]_net_1 )
        , .Y(hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[1]));
    CFG4 #( .INIT(16'hECA0) )  \PRDATA_0_iv_0_0_0[14]  (.A(
        \PRDATA_0_iv_0_0_a2[3]_net_1 ), .B(PRDATA4), .C(PRDATA_reg[14])
        , .D(lsram_width32_PRDATA[14]), .Y(
        \PRDATA_0_iv_0_0_0[14]_net_1 ));
    CFG4 #( .INIT(16'hECA0) )  \PRDATA_0_iv_0_0_0[12]  (.A(
        \PRDATA_0_iv_0_0_a2[3]_net_1 ), .B(PRDATA4), .C(PRDATA_reg[12])
        , .D(lsram_width32_PRDATA[12]), .Y(
        \PRDATA_0_iv_0_0_0[12]_net_1 ));
    CFG4 #( .INIT(16'hECA0) )  \PRDATA_0_iv_0_0_1[0]  (.A(
        \PRDATA_0_iv_0_0_a2[3]_net_1 ), .B(PRDATA4), .C(PRDATA_reg[0]), 
        .D(lsram_width32_PRDATA[0]), .Y(\PRDATA_0_iv_0_0_1[0]_net_1 ));
    CFG4 #( .INIT(16'h0001) )  \PRDATA_0_iv_0_0_a2_0_18_9[3]  (.A(
        hello_regs_MSS_0_FIC_0_APB_MASTER_PADDR[17]), .B(
        hello_regs_MSS_0_FIC_0_APB_MASTER_PADDR[23]), .C(
        hello_regs_MSS_0_FIC_0_APB_MASTER_PADDR[22]), .D(
        hello_regs_MSS_0_FIC_0_APB_MASTER_PADDR[18]), .Y(
        \PRDATA_0_iv_0_0_a2_0_18_9[3]_net_1 ));
    CFG4 #( .INIT(16'hFF80) )  \PRDATA_0_iv_0_0_0[6]  (.A(
        mem_8__2_i_0_0_a2[2]), .B(GPIO_OUT_1_c[6]), .C(
        PRDATA_0_iv_0_0_a2_2_4[3]), .D(\PRDATA_0_iv_0_0_a3_0[6]_net_1 )
        , .Y(\PRDATA_0_iv_0_0_0[6]_net_1 ));
    CFG4 #( .INIT(16'hF8F0) )  \PRDATA_0_iv_0_0[11]  (.A(
        PRDATA_0_iv_0_0_a2_0_17[3]), .B(IADDR_REG[11]), .C(
        \PRDATA_0_iv_0_0_0[11]_net_1 ), .D(PRDATA_0_iv_0_0_a2_0_18[3]), 
        .Y(hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[11]));
    CFG2 #( .INIT(4'h8) )  \PRDATA_0_iv_0_0_a3_0[7]  (.A(
        PRDATA_0_iv_0_0_a2_1[3]), .B(CoreAPB3_0_APBmslave5_PRDATA[7]), 
        .Y(\PRDATA_0_iv_0_0_a3_0[7]_net_1 ));
    CFG4 #( .INIT(16'hFF80) )  \PRDATA_0_iv_0_0_0[0]  (.A(
        mem_8__2_i_0_0_a2[2]), .B(GPIO_OUT_1_c[0]), .C(
        PRDATA_0_iv_0_0_a2_2_4[3]), .D(\PRDATA_0_iv_0_0_a3_0[0]_net_1 )
        , .Y(\PRDATA_0_iv_0_0_0[0]_net_1 ));
    CFG2 #( .INIT(4'h8) )  \PRDATA_0_iv_0_0_a3_0[5]  (.A(
        PRDATA_0_iv_0_0_a2_1[3]), .B(CoreAPB3_0_APBmslave5_PRDATA[5]), 
        .Y(\PRDATA_0_iv_0_0_a3_0[5]_net_1 ));
    CFG4 #( .INIT(16'hFF8F) )  \PRDATA_0_iv_0_0[3]  (.A(
        CoreAPB3_0_APBmslave5_PRDATA[3]), .B(PRDATA_0_iv_0_0_a2_1[3]), 
        .C(\PRDATA_0_iv_0_0_0[3]_net_1 ), .D(
        \PRDATA_0_iv_0_0_1[3]_net_1 ), .Y(
        hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[3]));
    CFG4 #( .INIT(16'hFFF8) )  \PRDATA_0_iv_0_0[7]  (.A(
        PRDATA_0_iv_0_0_a2_0_18[3]), .B(
        \PRDATA_0_iv_0_0_a3_3_0[7]_net_1 ), .C(
        \PRDATA_0_iv_0_0_1[7]_net_1 ), .D(\PRDATA_0_iv_0_0_0[7]_net_1 )
        , .Y(hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[7]));
    CFG4 #( .INIT(16'hF8F0) )  \PRDATA_0_iv_0_0[30]  (.A(
        PRDATA_0_iv_0_0_a2_0_17[3]), .B(IADDR_REG[30]), .C(
        \PRDATA_0_iv_0_0_0[30]_net_1 ), .D(PRDATA_0_iv_0_0_a2_0_18[3]), 
        .Y(hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[30]));
    CFG4 #( .INIT(16'hF8F0) )  \PRDATA_0_iv_0_0[28]  (.A(
        PRDATA_0_iv_0_0_a2_0_17[3]), .B(IADDR_REG[28]), .C(
        \PRDATA_0_iv_0_0_0[28]_net_1 ), .D(PRDATA_0_iv_0_0_a2_0_18[3]), 
        .Y(hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[28]));
    CFG4 #( .INIT(16'hECA0) )  \PRDATA_0_iv_0_0_1[4]  (.A(
        \PRDATA_0_iv_0_0_a2[3]_net_1 ), .B(PRDATA4), .C(PRDATA_reg[4]), 
        .D(lsram_width32_PRDATA[4]), .Y(\PRDATA_0_iv_0_0_1[4]_net_1 ));
    CFG4 #( .INIT(16'hFFF8) )  \PRDATA_0_iv_0_0[5]  (.A(
        PRDATA_0_iv_0_0_a2_0_18[3]), .B(
        \PRDATA_0_iv_0_0_a3_3_0[5]_net_1 ), .C(
        \PRDATA_0_iv_0_0_1[5]_net_1 ), .D(\PRDATA_0_iv_0_0_0[5]_net_1 )
        , .Y(hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[5]));
    CFG4 #( .INIT(16'hF8F0) )  \PRDATA_0_iv_0_0[17]  (.A(
        PRDATA_0_iv_0_0_a2_0_17[3]), .B(IADDR_REG[17]), .C(
        \PRDATA_0_iv_0_0_0[17]_net_1 ), .D(PRDATA_0_iv_0_0_a2_0_18[3]), 
        .Y(hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[17]));
    CFG4 #( .INIT(16'h8000) )  \PRDATA_0_iv_0_0_a3_3_0[2]  (.A(N_688), 
        .B(IADDR_REG[2]), .C(\PRDATA_0_iv_0_0_a2_0_17_2[3]_net_1 ), .D(
        mem_0__2_i_0_0_a2[0]), .Y(\PRDATA_0_iv_0_0_a3_3_0[2]_net_1 ));
    CFG4 #( .INIT(16'hF8F0) )  \PRDATA_0_iv_0_0[12]  (.A(
        PRDATA_0_iv_0_0_a2_0_17[3]), .B(IADDR_REG[12]), .C(
        \PRDATA_0_iv_0_0_0[12]_net_1 ), .D(PRDATA_0_iv_0_0_a2_0_18[3]), 
        .Y(hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[12]));
    CFG4 #( .INIT(16'h0080) )  \PRDATA_0_iv_0_0_a2_2_4_2[3]  (.A(
        CoreAPB3_0_APBmslave4_PADDR_7), .B(
        hello_regs_MSS_0_FIC_0_APB_MASTER_PADDR[25]), .C(
        hello_regs_MSS_0_FIC_0_APB_MASTER_PADDR[26]), .D(
        hello_regs_MSS_0_FIC_0_APB_MASTER_PADDR[24]), .Y(
        \PRDATA_0_iv_0_0_a2_2_4_2[3]_net_1 ));
    CFG4 #( .INIT(16'hECA0) )  \PRDATA_0_iv_0_0_1[2]  (.A(
        \PRDATA_0_iv_0_0_a2[3]_net_1 ), .B(PRDATA4), .C(PRDATA_reg[2]), 
        .D(lsram_width32_PRDATA[2]), .Y(\PRDATA_0_iv_0_0_1[2]_net_1 ));
    CFG4 #( .INIT(16'hF8F0) )  \PRDATA_0_iv_0_0[21]  (.A(
        PRDATA_0_iv_0_0_a2_0_17[3]), .B(IADDR_REG[21]), .C(
        \PRDATA_0_iv_0_0_0[21]_net_1 ), .D(PRDATA_0_iv_0_0_a2_0_18[3]), 
        .Y(hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[21]));
    CFG4 #( .INIT(16'h8000) )  \PRDATA_0_iv_0_0_a3_1_0[9]  (.A(N_688), 
        .B(IADDR_REG[9]), .C(\PRDATA_0_iv_0_0_a2_0_17_2[3]_net_1 ), .D(
        mem_0__2_i_0_0_a2[0]), .Y(\PRDATA_0_iv_0_0_a3_1_0[9]_net_1 ));
    CFG4 #( .INIT(16'h007F) )  \PRDATA_0_iv_0_0_0[3]  (.A(
        PRDATA_0_iv_0_0_a2_0_17[3]), .B(PRDATA_0_iv_0_0_a2_0_18[3]), 
        .C(IADDR_REG[3]), .D(\PRDATA_0_iv_0_0_a3[3]_net_1 ), .Y(
        \PRDATA_0_iv_0_0_0[3]_net_1 ));
    CFG4 #( .INIT(16'hECA0) )  \PRDATA_0_iv_0_0_0[11]  (.A(
        \PRDATA_0_iv_0_0_a2[3]_net_1 ), .B(PRDATA4), .C(PRDATA_reg[11])
        , .D(lsram_width32_PRDATA[11]), .Y(
        \PRDATA_0_iv_0_0_0[11]_net_1 ));
    CFG4 #( .INIT(16'hF8F0) )  \PRDATA_0_iv_0_0[16]  (.A(
        PRDATA_0_iv_0_0_a2_0_17[3]), .B(IADDR_REG[16]), .C(
        \PRDATA_0_iv_0_0_0[16]_net_1 ), .D(PRDATA_0_iv_0_0_a2_0_18[3]), 
        .Y(hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[16]));
    CFG4 #( .INIT(16'h8000) )  \PRDATA_0_iv_0_0_a2_0_18[3]  (.A(N_928), 
        .B(\PRDATA_0_iv_0_0_a2_0_18_1[3]_net_1 ), .C(
        \PRDATA_0_iv_0_0_a2_0_18_8[3]_net_1 ), .D(
        \PRDATA_0_iv_0_0_a2_0_18_9[3]_net_1 ), .Y(
        PRDATA_0_iv_0_0_a2_0_18[3]));
    CFG4 #( .INIT(16'hECA0) )  \PRDATA_0_iv_0_0_0[23]  (.A(
        \PRDATA_0_iv_0_0_a2[3]_net_1 ), .B(PRDATA4), .C(PRDATA_reg[23])
        , .D(lsram_width32_PRDATA[23]), .Y(
        \PRDATA_0_iv_0_0_0[23]_net_1 ));
    CFG4 #( .INIT(16'hECA0) )  \PRDATA_0_iv_0_0_0[17]  (.A(
        \PRDATA_0_iv_0_0_a2[3]_net_1 ), .B(PRDATA4), .C(PRDATA_reg[17])
        , .D(lsram_width32_PRDATA[17]), .Y(
        \PRDATA_0_iv_0_0_0[17]_net_1 ));
    CFG4 #( .INIT(16'hF8F0) )  \PRDATA_0_iv_0_0[27]  (.A(
        PRDATA_0_iv_0_0_a2_0_17[3]), .B(IADDR_REG[27]), .C(
        \PRDATA_0_iv_0_0_0[27]_net_1 ), .D(PRDATA_0_iv_0_0_a2_0_18[3]), 
        .Y(hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[27]));
    CFG4 #( .INIT(16'hF8F0) )  \PRDATA_0_iv_0_0[22]  (.A(
        PRDATA_0_iv_0_0_a2_0_17[3]), .B(IADDR_REG[22]), .C(
        \PRDATA_0_iv_0_0_0[22]_net_1 ), .D(PRDATA_0_iv_0_0_a2_0_18[3]), 
        .Y(hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[22]));
    CFG4 #( .INIT(16'h8000) )  \PRDATA_0_iv_0_0_a3_3_0[6]  (.A(N_688), 
        .B(IADDR_REG[6]), .C(\PRDATA_0_iv_0_0_a2_0_17_2[3]_net_1 ), .D(
        mem_0__2_i_0_0_a2[0]), .Y(\PRDATA_0_iv_0_0_a3_3_0[6]_net_1 ));
    CFG4 #( .INIT(16'h8000) )  \PRDATA_0_iv_0_0_a3_3_0[7]  (.A(N_688), 
        .B(IADDR_REG[7]), .C(\PRDATA_0_iv_0_0_a2_0_17_2[3]_net_1 ), .D(
        mem_0__2_i_0_0_a2[0]), .Y(\PRDATA_0_iv_0_0_a3_3_0[7]_net_1 ));
    CFG4 #( .INIT(16'h8000) )  \PRDATA_0_iv_0_0_a3_1_0[23]  (.A(N_688), 
        .B(IADDR_REG[23]), .C(\PRDATA_0_iv_0_0_a2_0_17_2[3]_net_1 ), 
        .D(mem_0__2_i_0_0_a2[0]), .Y(
        \PRDATA_0_iv_0_0_a3_1_0[23]_net_1 ));
    CFG3 #( .INIT(8'h10) )  \PRDATA_0_iv_0_0_a2_0_18_1[3]  (.A(
        hello_regs_MSS_0_FIC_0_APB_MASTER_PADDR[10]), .B(
        CoreAPB3_0_APBmslave4_PADDR_8), .C(
        \PRDATA_0_iv_0_0_a2_0_18_7[3]_net_1 ), .Y(
        \PRDATA_0_iv_0_0_a2_0_18_1[3]_net_1 ));
    CFG4 #( .INIT(16'hFF80) )  \PRDATA_0_iv_0_0_0[5]  (.A(
        mem_8__2_i_0_0_a2[2]), .B(GPIO_OUT_1_c[5]), .C(
        PRDATA_0_iv_0_0_a2_2_4[3]), .D(\PRDATA_0_iv_0_0_a3_0[5]_net_1 )
        , .Y(\PRDATA_0_iv_0_0_0[5]_net_1 ));
    CFG4 #( .INIT(16'hECA0) )  \PRDATA_0_iv_0_0_0[16]  (.A(
        \PRDATA_0_iv_0_0_a2[3]_net_1 ), .B(PRDATA4), .C(PRDATA_reg[16])
        , .D(lsram_width32_PRDATA[16]), .Y(
        \PRDATA_0_iv_0_0_0[16]_net_1 ));
    CFG4 #( .INIT(16'h0001) )  \PRDATA_0_iv_0_0_a2_0_18_7[3]  (.A(
        CoreAPB3_0_APBmslave4_PADDR_7), .B(
        hello_regs_MSS_0_FIC_0_APB_MASTER_PADDR[16]), .C(
        hello_regs_MSS_0_FIC_0_APB_MASTER_PADDR[15]), .D(
        hello_regs_MSS_0_FIC_0_APB_MASTER_PADDR[11]), .Y(
        \PRDATA_0_iv_0_0_a2_0_18_7[3]_net_1 ));
    CFG4 #( .INIT(16'h0001) )  \PRDATA_0_iv_0_0_a2_0_17_2[3]  (.A(
        hello_regs_MSS_0_FIC_0_APB_MASTER_PADDR[21]), .B(
        hello_regs_MSS_0_FIC_0_APB_MASTER_PADDR[9]), .C(
        hello_regs_MSS_0_FIC_0_APB_MASTER_PADDR[19]), .D(
        hello_regs_MSS_0_FIC_0_APB_MASTER_PADDR[26]), .Y(
        \PRDATA_0_iv_0_0_a2_0_17_2[3]_net_1 ));
    CFG4 #( .INIT(16'hFF80) )  \PRDATA_0_iv_0_0_0[4]  (.A(
        mem_8__2_i_0_0_a2[2]), .B(GPIO_OUT_1_c[4]), .C(
        PRDATA_0_iv_0_0_a2_2_4[3]), .D(\PRDATA_0_iv_0_0_a3_0[4]_net_1 )
        , .Y(\PRDATA_0_iv_0_0_0[4]_net_1 ));
    CFG4 #( .INIT(16'hF8F0) )  \PRDATA_0_iv_0_0[26]  (.A(
        PRDATA_0_iv_0_0_a2_0_17[3]), .B(IADDR_REG[26]), .C(
        \PRDATA_0_iv_0_0_0[26]_net_1 ), .D(PRDATA_0_iv_0_0_a2_0_18[3]), 
        .Y(hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[26]));
    CFG4 #( .INIT(16'h8000) )  \PRDATA_0_iv_0_0_a3_3_0[1]  (.A(N_688), 
        .B(IADDR_REG[1]), .C(\PRDATA_0_iv_0_0_a2_0_17_2[3]_net_1 ), .D(
        mem_0__2_i_0_0_a2[0]), .Y(\PRDATA_0_iv_0_0_a3_3_0[1]_net_1 ));
    CFG4 #( .INIT(16'hECA0) )  \PRDATA_0_iv_0_0_1[7]  (.A(
        \PRDATA_0_iv_0_0_a2[3]_net_1 ), .B(PRDATA4), .C(PRDATA_reg[7]), 
        .D(lsram_width32_PRDATA[7]), .Y(\PRDATA_0_iv_0_0_1[7]_net_1 ));
    CFG2 #( .INIT(4'h8) )  \PRDATA_0_iv_0_0_a3_0[6]  (.A(
        PRDATA_0_iv_0_0_a2_1[3]), .B(CoreAPB3_0_APBmslave5_PRDATA[6]), 
        .Y(\PRDATA_0_iv_0_0_a3_0[6]_net_1 ));
    CFG2 #( .INIT(4'h8) )  \PRDATA_0_iv_0_0_a3_0[2]  (.A(
        PRDATA_0_iv_0_0_a2_1[3]), .B(CoreAPB3_0_APBmslave5_PRDATA[2]), 
        .Y(\PRDATA_0_iv_0_0_a3_0[2]_net_1 ));
    CFG4 #( .INIT(16'hECA0) )  \PRDATA_0_iv_0_0_0[15]  (.A(
        \PRDATA_0_iv_0_0_a2[3]_net_1 ), .B(PRDATA4), .C(PRDATA_reg[15])
        , .D(lsram_width32_PRDATA[15]), .Y(
        \PRDATA_0_iv_0_0_0[15]_net_1 ));
    
endmodule


module CoreAPB3_Z1(
       PRDATA_0_iv_0_0_a2_1,
       hello_regs_MSS_0_FIC_0_APB_MASTER_PADDR,
       mem_8__2_i_0_0_a2,
       mem_0__2_i_0_0_a2,
       PRDATA_0_iv_0_0_a2_2_4,
       CoreAPB3_0_APBmslave5_PRDATA,
       PRDATA_reg,
       lsram_width32_PRDATA,
       GPIO_OUT_1_c,
       hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA,
       CoreAPB3_0_APBmslave4_PWDATA,
       CoreAPB3_0_APBmslave4_PADDR_8,
       CoreAPB3_0_APBmslave4_PADDR_7,
       CoreAPB3_0_APBmslave4_PADDR_0,
       CoreAPB3_0_APBmslave4_PADDR_6,
       CoreAPB3_0_APBmslave4_PADDR_1,
       hello_regs_MSS_0_FIC_0_APB_MASTER_PSELx,
       N_928,
       CoreAPB3_0_APBmslave4_PWRITE,
       CoreAPB3_0_APBmslave4_PENABLE,
       PRDATA4,
       CoreAPB3_0_APBmslave4_PREADY,
       N_676_i_0,
       MSS_RESET_N_M2F_c,
       FCCC_0_GL1
    );
output [3:3] PRDATA_0_iv_0_0_a2_1;
input  [27:9] hello_regs_MSS_0_FIC_0_APB_MASTER_PADDR;
input  [2:2] mem_8__2_i_0_0_a2;
input  [0:0] mem_0__2_i_0_0_a2;
output [3:3] PRDATA_0_iv_0_0_a2_2_4;
input  [7:0] CoreAPB3_0_APBmslave5_PRDATA;
input  [31:0] PRDATA_reg;
input  [31:0] lsram_width32_PRDATA;
input  [7:0] GPIO_OUT_1_c;
output [31:0] hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA;
input  [31:0] CoreAPB3_0_APBmslave4_PWDATA;
input  CoreAPB3_0_APBmslave4_PADDR_8;
input  CoreAPB3_0_APBmslave4_PADDR_7;
input  CoreAPB3_0_APBmslave4_PADDR_0;
input  CoreAPB3_0_APBmslave4_PADDR_6;
input  CoreAPB3_0_APBmslave4_PADDR_1;
input  hello_regs_MSS_0_FIC_0_APB_MASTER_PSELx;
input  N_928;
input  CoreAPB3_0_APBmslave4_PWRITE;
input  CoreAPB3_0_APBmslave4_PENABLE;
input  PRDATA4;
input  CoreAPB3_0_APBmslave4_PREADY;
output N_676_i_0;
input  MSS_RESET_N_M2F_c;
input  FCCC_0_GL1;

    wire \PRDATA_0_iv_0_0_a2_0_17[3] , \PRDATA_0_iv_0_0_a2_0_18[3] , 
        \IADDR_REG[0] , \IADDR_REG[1] , \IADDR_REG[2] , \IADDR_REG[3] , 
        \IADDR_REG[4] , \IADDR_REG[5] , \IADDR_REG[6] , \IADDR_REG[7] , 
        \IADDR_REG[8] , \IADDR_REG[9] , \IADDR_REG[10] , 
        \IADDR_REG[11] , \IADDR_REG[12] , \IADDR_REG[13] , 
        \IADDR_REG[14] , \IADDR_REG[15] , \IADDR_REG[16] , 
        \IADDR_REG[17] , \IADDR_REG[18] , \IADDR_REG[19] , 
        \IADDR_REG[20] , \IADDR_REG[21] , \IADDR_REG[22] , 
        \IADDR_REG[23] , \IADDR_REG[24] , \IADDR_REG[25] , 
        \IADDR_REG[26] , \IADDR_REG[27] , \IADDR_REG[28] , 
        \IADDR_REG[29] , \IADDR_REG[30] , \IADDR_REG[31] , GND_net_1, 
        VCC_net_1;
    
    coreapb3_iaddr_reg_0s_32_28 \g_iaddr_reg.genblk3.iaddr_reg  (
        .IADDR_REG({\IADDR_REG[31] , \IADDR_REG[30] , \IADDR_REG[29] , 
        \IADDR_REG[28] , \IADDR_REG[27] , \IADDR_REG[26] , 
        \IADDR_REG[25] , \IADDR_REG[24] , \IADDR_REG[23] , 
        \IADDR_REG[22] , \IADDR_REG[21] , \IADDR_REG[20] , 
        \IADDR_REG[19] , \IADDR_REG[18] , \IADDR_REG[17] , 
        \IADDR_REG[16] , \IADDR_REG[15] , \IADDR_REG[14] , 
        \IADDR_REG[13] , \IADDR_REG[12] , \IADDR_REG[11] , 
        \IADDR_REG[10] , \IADDR_REG[9] , \IADDR_REG[8] , 
        \IADDR_REG[7] , \IADDR_REG[6] , \IADDR_REG[5] , \IADDR_REG[4] , 
        \IADDR_REG[3] , \IADDR_REG[2] , \IADDR_REG[1] , \IADDR_REG[0] })
        , .CoreAPB3_0_APBmslave4_PWDATA({
        CoreAPB3_0_APBmslave4_PWDATA[31], 
        CoreAPB3_0_APBmslave4_PWDATA[30], 
        CoreAPB3_0_APBmslave4_PWDATA[29], 
        CoreAPB3_0_APBmslave4_PWDATA[28], 
        CoreAPB3_0_APBmslave4_PWDATA[27], 
        CoreAPB3_0_APBmslave4_PWDATA[26], 
        CoreAPB3_0_APBmslave4_PWDATA[25], 
        CoreAPB3_0_APBmslave4_PWDATA[24], 
        CoreAPB3_0_APBmslave4_PWDATA[23], 
        CoreAPB3_0_APBmslave4_PWDATA[22], 
        CoreAPB3_0_APBmslave4_PWDATA[21], 
        CoreAPB3_0_APBmslave4_PWDATA[20], 
        CoreAPB3_0_APBmslave4_PWDATA[19], 
        CoreAPB3_0_APBmslave4_PWDATA[18], 
        CoreAPB3_0_APBmslave4_PWDATA[17], 
        CoreAPB3_0_APBmslave4_PWDATA[16], 
        CoreAPB3_0_APBmslave4_PWDATA[15], 
        CoreAPB3_0_APBmslave4_PWDATA[14], 
        CoreAPB3_0_APBmslave4_PWDATA[13], 
        CoreAPB3_0_APBmslave4_PWDATA[12], 
        CoreAPB3_0_APBmslave4_PWDATA[11], 
        CoreAPB3_0_APBmslave4_PWDATA[10], 
        CoreAPB3_0_APBmslave4_PWDATA[9], 
        CoreAPB3_0_APBmslave4_PWDATA[8], 
        CoreAPB3_0_APBmslave4_PWDATA[7], 
        CoreAPB3_0_APBmslave4_PWDATA[6], 
        CoreAPB3_0_APBmslave4_PWDATA[5], 
        CoreAPB3_0_APBmslave4_PWDATA[4], 
        CoreAPB3_0_APBmslave4_PWDATA[3], 
        CoreAPB3_0_APBmslave4_PWDATA[2], 
        CoreAPB3_0_APBmslave4_PWDATA[1], 
        CoreAPB3_0_APBmslave4_PWDATA[0]}), .PRDATA_0_iv_0_0_a2_0_18({
        \PRDATA_0_iv_0_0_a2_0_18[3] }), .PRDATA_0_iv_0_0_a2_0_17({
        \PRDATA_0_iv_0_0_a2_0_17[3] }), .MSS_RESET_N_M2F_c(
        MSS_RESET_N_M2F_c), .FCCC_0_GL1(FCCC_0_GL1), 
        .CoreAPB3_0_APBmslave4_PENABLE(CoreAPB3_0_APBmslave4_PENABLE), 
        .CoreAPB3_0_APBmslave4_PWRITE(CoreAPB3_0_APBmslave4_PWRITE));
    VCC VCC (.Y(VCC_net_1));
    COREAPB3_MUXPTOB3 u_mux_p_to_b3 (.PRDATA_0_iv_0_0_a2_1({
        PRDATA_0_iv_0_0_a2_1[3]}), .PRDATA_0_iv_0_0_a2_0_17({
        \PRDATA_0_iv_0_0_a2_0_17[3] }), .PRDATA_0_iv_0_0_a2_0_18({
        \PRDATA_0_iv_0_0_a2_0_18[3] }), 
        .hello_regs_MSS_0_FIC_0_APB_MASTER_PADDR({
        hello_regs_MSS_0_FIC_0_APB_MASTER_PADDR[27], 
        hello_regs_MSS_0_FIC_0_APB_MASTER_PADDR[26], 
        hello_regs_MSS_0_FIC_0_APB_MASTER_PADDR[25], 
        hello_regs_MSS_0_FIC_0_APB_MASTER_PADDR[24], 
        hello_regs_MSS_0_FIC_0_APB_MASTER_PADDR[23], 
        hello_regs_MSS_0_FIC_0_APB_MASTER_PADDR[22], 
        hello_regs_MSS_0_FIC_0_APB_MASTER_PADDR[21], 
        hello_regs_MSS_0_FIC_0_APB_MASTER_PADDR[20], 
        hello_regs_MSS_0_FIC_0_APB_MASTER_PADDR[19], 
        hello_regs_MSS_0_FIC_0_APB_MASTER_PADDR[18], 
        hello_regs_MSS_0_FIC_0_APB_MASTER_PADDR[17], 
        hello_regs_MSS_0_FIC_0_APB_MASTER_PADDR[16], 
        hello_regs_MSS_0_FIC_0_APB_MASTER_PADDR[15], 
        hello_regs_MSS_0_FIC_0_APB_MASTER_PADDR[14], 
        hello_regs_MSS_0_FIC_0_APB_MASTER_PADDR[13], 
        hello_regs_MSS_0_FIC_0_APB_MASTER_PADDR[12], 
        hello_regs_MSS_0_FIC_0_APB_MASTER_PADDR[11], 
        hello_regs_MSS_0_FIC_0_APB_MASTER_PADDR[10], 
        hello_regs_MSS_0_FIC_0_APB_MASTER_PADDR[9]}), 
        .mem_8__2_i_0_0_a2({mem_8__2_i_0_0_a2[2]}), .mem_0__2_i_0_0_a2({
        mem_0__2_i_0_0_a2[0]}), .PRDATA_0_iv_0_0_a2_2_4({
        PRDATA_0_iv_0_0_a2_2_4[3]}), .CoreAPB3_0_APBmslave5_PRDATA({
        CoreAPB3_0_APBmslave5_PRDATA[7], 
        CoreAPB3_0_APBmslave5_PRDATA[6], 
        CoreAPB3_0_APBmslave5_PRDATA[5], 
        CoreAPB3_0_APBmslave5_PRDATA[4], 
        CoreAPB3_0_APBmslave5_PRDATA[3], 
        CoreAPB3_0_APBmslave5_PRDATA[2], 
        CoreAPB3_0_APBmslave5_PRDATA[1], 
        CoreAPB3_0_APBmslave5_PRDATA[0]}), .PRDATA_reg({PRDATA_reg[31], 
        PRDATA_reg[30], PRDATA_reg[29], PRDATA_reg[28], PRDATA_reg[27], 
        PRDATA_reg[26], PRDATA_reg[25], PRDATA_reg[24], PRDATA_reg[23], 
        PRDATA_reg[22], PRDATA_reg[21], PRDATA_reg[20], PRDATA_reg[19], 
        PRDATA_reg[18], PRDATA_reg[17], PRDATA_reg[16], PRDATA_reg[15], 
        PRDATA_reg[14], PRDATA_reg[13], PRDATA_reg[12], PRDATA_reg[11], 
        PRDATA_reg[10], PRDATA_reg[9], PRDATA_reg[8], PRDATA_reg[7], 
        PRDATA_reg[6], PRDATA_reg[5], PRDATA_reg[4], PRDATA_reg[3], 
        PRDATA_reg[2], PRDATA_reg[1], PRDATA_reg[0]}), 
        .lsram_width32_PRDATA({lsram_width32_PRDATA[31], 
        lsram_width32_PRDATA[30], lsram_width32_PRDATA[29], 
        lsram_width32_PRDATA[28], lsram_width32_PRDATA[27], 
        lsram_width32_PRDATA[26], lsram_width32_PRDATA[25], 
        lsram_width32_PRDATA[24], lsram_width32_PRDATA[23], 
        lsram_width32_PRDATA[22], lsram_width32_PRDATA[21], 
        lsram_width32_PRDATA[20], lsram_width32_PRDATA[19], 
        lsram_width32_PRDATA[18], lsram_width32_PRDATA[17], 
        lsram_width32_PRDATA[16], lsram_width32_PRDATA[15], 
        lsram_width32_PRDATA[14], lsram_width32_PRDATA[13], 
        lsram_width32_PRDATA[12], lsram_width32_PRDATA[11], 
        lsram_width32_PRDATA[10], lsram_width32_PRDATA[9], 
        lsram_width32_PRDATA[8], lsram_width32_PRDATA[7], 
        lsram_width32_PRDATA[6], lsram_width32_PRDATA[5], 
        lsram_width32_PRDATA[4], lsram_width32_PRDATA[3], 
        lsram_width32_PRDATA[2], lsram_width32_PRDATA[1], 
        lsram_width32_PRDATA[0]}), .GPIO_OUT_1_c({GPIO_OUT_1_c[7], 
        GPIO_OUT_1_c[6], GPIO_OUT_1_c[5], GPIO_OUT_1_c[4], 
        GPIO_OUT_1_c[3], GPIO_OUT_1_c[2], GPIO_OUT_1_c[1], 
        GPIO_OUT_1_c[0]}), .IADDR_REG({\IADDR_REG[31] , 
        \IADDR_REG[30] , \IADDR_REG[29] , \IADDR_REG[28] , 
        \IADDR_REG[27] , \IADDR_REG[26] , \IADDR_REG[25] , 
        \IADDR_REG[24] , \IADDR_REG[23] , \IADDR_REG[22] , 
        \IADDR_REG[21] , \IADDR_REG[20] , \IADDR_REG[19] , 
        \IADDR_REG[18] , \IADDR_REG[17] , \IADDR_REG[16] , 
        \IADDR_REG[15] , \IADDR_REG[14] , \IADDR_REG[13] , 
        \IADDR_REG[12] , \IADDR_REG[11] , \IADDR_REG[10] , 
        \IADDR_REG[9] , \IADDR_REG[8] , \IADDR_REG[7] , \IADDR_REG[6] , 
        \IADDR_REG[5] , \IADDR_REG[4] , \IADDR_REG[3] , \IADDR_REG[2] , 
        \IADDR_REG[1] , \IADDR_REG[0] }), 
        .hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA({
        hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[31], 
        hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[30], 
        hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[29], 
        hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[28], 
        hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[27], 
        hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[26], 
        hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[25], 
        hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[24], 
        hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[23], 
        hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[22], 
        hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[21], 
        hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[20], 
        hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[19], 
        hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[18], 
        hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[17], 
        hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[16], 
        hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[15], 
        hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[14], 
        hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[13], 
        hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[12], 
        hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[11], 
        hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[10], 
        hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[9], 
        hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[8], 
        hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[7], 
        hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[6], 
        hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[5], 
        hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[4], 
        hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[3], 
        hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[2], 
        hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[1], 
        hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[0]}), 
        .CoreAPB3_0_APBmslave4_PADDR_8(CoreAPB3_0_APBmslave4_PADDR_8), 
        .CoreAPB3_0_APBmslave4_PADDR_7(CoreAPB3_0_APBmslave4_PADDR_7), 
        .CoreAPB3_0_APBmslave4_PADDR_0(CoreAPB3_0_APBmslave4_PADDR_0), 
        .CoreAPB3_0_APBmslave4_PADDR_6(CoreAPB3_0_APBmslave4_PADDR_6), 
        .CoreAPB3_0_APBmslave4_PADDR_1(CoreAPB3_0_APBmslave4_PADDR_1), 
        .hello_regs_MSS_0_FIC_0_APB_MASTER_PSELx(
        hello_regs_MSS_0_FIC_0_APB_MASTER_PSELx), .N_928(N_928), 
        .CoreAPB3_0_APBmslave4_PWRITE(CoreAPB3_0_APBmslave4_PWRITE), 
        .CoreAPB3_0_APBmslave4_PENABLE(CoreAPB3_0_APBmslave4_PENABLE), 
        .PRDATA4(PRDATA4), .CoreAPB3_0_APBmslave4_PREADY(
        CoreAPB3_0_APBmslave4_PREADY), .N_676_i_0(N_676_i_0));
    GND GND (.Y(GND_net_1));
    
endmodule


module hello_regs_OSC_0_OSC(
       OSC_0_RCOSC_25_50MHZ_CCC_OUT_RCOSC_25_50MHZ_CCC
    );
output OSC_0_RCOSC_25_50MHZ_CCC_OUT_RCOSC_25_50MHZ_CCC;

    wire GND_net_1, VCC_net_1;
    
    RCOSC_25_50MHZ #( .FREQUENCY(50.0) )  I_RCOSC_25_50MHZ (.CLKOUT(
        OSC_0_RCOSC_25_50MHZ_CCC_OUT_RCOSC_25_50MHZ_CCC));
    VCC VCC (.Y(VCC_net_1));
    GND GND (.Y(GND_net_1));
    
endmodule


module hello_regs_MSS(
       CoreAPB3_0_APBmslave4_PADDR,
       hello_regs_MSS_0_FIC_0_APB_MASTER_PADDR,
       CoreAPB3_0_APBmslave4_PWDATA,
       hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA,
       MSS_RESET_N_M2F_c,
       MMUART_0_TXD,
       MMUART_0_RXD,
       CoreAPB3_0_APBmslave4_PENABLE,
       hello_regs_MSS_0_FIC_0_APB_MASTER_PSELx,
       CoreAPB3_0_APBmslave4_PWRITE,
       N_676_i_0,
       FCCC_0_LOCK,
       FCCC_0_GL1
    );
output [8:0] CoreAPB3_0_APBmslave4_PADDR;
output [27:9] hello_regs_MSS_0_FIC_0_APB_MASTER_PADDR;
output [31:0] CoreAPB3_0_APBmslave4_PWDATA;
input  [31:0] hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA;
output MSS_RESET_N_M2F_c;
output MMUART_0_TXD;
input  MMUART_0_RXD;
output CoreAPB3_0_APBmslave4_PENABLE;
output hello_regs_MSS_0_FIC_0_APB_MASTER_PSELx;
output CoreAPB3_0_APBmslave4_PWRITE;
input  N_676_i_0;
input  FCCC_0_LOCK;
input  FCCC_0_GL1;

    wire FPGA_RESET_N, 
        MSS_ADLIB_INST_MMUART0_TXD_USBC_DIR_MGPIO27B_OUT, 
        MSS_ADLIB_INST_MMUART0_TXD_USBC_DIR_MGPIO27B_OE, 
        MMUART_0_RXD_PAD_Y, VCC_net_1, GND_net_1;
    
    INBUF MMUART_0_RXD_PAD (.PAD(MMUART_0_RXD), .Y(MMUART_0_RXD_PAD_Y));
    VCC VCC (.Y(VCC_net_1));
    CLKINT MSS_ADLIB_INST_RNIUO3B (.A(FPGA_RESET_N), .Y(
        MSS_RESET_N_M2F_c));
    MSS_010 #( .INIT(1438'h00000000003612000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000F00000000F000000000000000000000000000000007FFFFFFFB000001007C33C000000006092C0104003FFFFE400000000000010000000000F41C000001FEDFDC010842108421000001FE34001FF8000000400000000020091007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF)
        , .ACT_UBITS(56'hFFFFFFFFFFFFFF), .MEMORYFILE("ENVM_init.mem")
        , .RTC_MAIN_XTL_FREQ(0.0), .RTC_MAIN_XTL_MODE("") )  
        MSS_ADLIB_INST (.CAN_RXBUS_MGPIO3A_H2F_A(), 
        .CAN_RXBUS_MGPIO3A_H2F_B(), .CAN_TX_EBL_MGPIO4A_H2F_A(), 
        .CAN_TX_EBL_MGPIO4A_H2F_B(), .CAN_TXBUS_MGPIO2A_H2F_A(), 
        .CAN_TXBUS_MGPIO2A_H2F_B(), .CLK_CONFIG_APB(), .COMMS_INT(), 
        .CONFIG_PRESET_N(), .EDAC_ERROR({nc0, nc1, nc2, nc3, nc4, nc5, 
        nc6, nc7}), .F_FM0_RDATA({nc8, nc9, nc10, nc11, nc12, nc13, 
        nc14, nc15, nc16, nc17, nc18, nc19, nc20, nc21, nc22, nc23, 
        nc24, nc25, nc26, nc27, nc28, nc29, nc30, nc31, nc32, nc33, 
        nc34, nc35, nc36, nc37, nc38, nc39}), .F_FM0_READYOUT(), 
        .F_FM0_RESP(), .F_HM0_ADDR({nc40, nc41, nc42, nc43, 
        hello_regs_MSS_0_FIC_0_APB_MASTER_PADDR[27], 
        hello_regs_MSS_0_FIC_0_APB_MASTER_PADDR[26], 
        hello_regs_MSS_0_FIC_0_APB_MASTER_PADDR[25], 
        hello_regs_MSS_0_FIC_0_APB_MASTER_PADDR[24], 
        hello_regs_MSS_0_FIC_0_APB_MASTER_PADDR[23], 
        hello_regs_MSS_0_FIC_0_APB_MASTER_PADDR[22], 
        hello_regs_MSS_0_FIC_0_APB_MASTER_PADDR[21], 
        hello_regs_MSS_0_FIC_0_APB_MASTER_PADDR[20], 
        hello_regs_MSS_0_FIC_0_APB_MASTER_PADDR[19], 
        hello_regs_MSS_0_FIC_0_APB_MASTER_PADDR[18], 
        hello_regs_MSS_0_FIC_0_APB_MASTER_PADDR[17], 
        hello_regs_MSS_0_FIC_0_APB_MASTER_PADDR[16], 
        hello_regs_MSS_0_FIC_0_APB_MASTER_PADDR[15], 
        hello_regs_MSS_0_FIC_0_APB_MASTER_PADDR[14], 
        hello_regs_MSS_0_FIC_0_APB_MASTER_PADDR[13], 
        hello_regs_MSS_0_FIC_0_APB_MASTER_PADDR[12], 
        hello_regs_MSS_0_FIC_0_APB_MASTER_PADDR[11], 
        hello_regs_MSS_0_FIC_0_APB_MASTER_PADDR[10], 
        hello_regs_MSS_0_FIC_0_APB_MASTER_PADDR[9], 
        CoreAPB3_0_APBmslave4_PADDR[8], CoreAPB3_0_APBmslave4_PADDR[7], 
        CoreAPB3_0_APBmslave4_PADDR[6], CoreAPB3_0_APBmslave4_PADDR[5], 
        CoreAPB3_0_APBmslave4_PADDR[4], CoreAPB3_0_APBmslave4_PADDR[3], 
        CoreAPB3_0_APBmslave4_PADDR[2], CoreAPB3_0_APBmslave4_PADDR[1], 
        CoreAPB3_0_APBmslave4_PADDR[0]}), .F_HM0_ENABLE(
        CoreAPB3_0_APBmslave4_PENABLE), .F_HM0_SEL(
        hello_regs_MSS_0_FIC_0_APB_MASTER_PSELx), .F_HM0_SIZE({nc44, 
        nc45}), .F_HM0_TRANS1(), .F_HM0_WDATA({
        CoreAPB3_0_APBmslave4_PWDATA[31], 
        CoreAPB3_0_APBmslave4_PWDATA[30], 
        CoreAPB3_0_APBmslave4_PWDATA[29], 
        CoreAPB3_0_APBmslave4_PWDATA[28], 
        CoreAPB3_0_APBmslave4_PWDATA[27], 
        CoreAPB3_0_APBmslave4_PWDATA[26], 
        CoreAPB3_0_APBmslave4_PWDATA[25], 
        CoreAPB3_0_APBmslave4_PWDATA[24], 
        CoreAPB3_0_APBmslave4_PWDATA[23], 
        CoreAPB3_0_APBmslave4_PWDATA[22], 
        CoreAPB3_0_APBmslave4_PWDATA[21], 
        CoreAPB3_0_APBmslave4_PWDATA[20], 
        CoreAPB3_0_APBmslave4_PWDATA[19], 
        CoreAPB3_0_APBmslave4_PWDATA[18], 
        CoreAPB3_0_APBmslave4_PWDATA[17], 
        CoreAPB3_0_APBmslave4_PWDATA[16], 
        CoreAPB3_0_APBmslave4_PWDATA[15], 
        CoreAPB3_0_APBmslave4_PWDATA[14], 
        CoreAPB3_0_APBmslave4_PWDATA[13], 
        CoreAPB3_0_APBmslave4_PWDATA[12], 
        CoreAPB3_0_APBmslave4_PWDATA[11], 
        CoreAPB3_0_APBmslave4_PWDATA[10], 
        CoreAPB3_0_APBmslave4_PWDATA[9], 
        CoreAPB3_0_APBmslave4_PWDATA[8], 
        CoreAPB3_0_APBmslave4_PWDATA[7], 
        CoreAPB3_0_APBmslave4_PWDATA[6], 
        CoreAPB3_0_APBmslave4_PWDATA[5], 
        CoreAPB3_0_APBmslave4_PWDATA[4], 
        CoreAPB3_0_APBmslave4_PWDATA[3], 
        CoreAPB3_0_APBmslave4_PWDATA[2], 
        CoreAPB3_0_APBmslave4_PWDATA[1], 
        CoreAPB3_0_APBmslave4_PWDATA[0]}), .F_HM0_WRITE(
        CoreAPB3_0_APBmslave4_PWRITE), .FAB_CHRGVBUS(), 
        .FAB_DISCHRGVBUS(), .FAB_DMPULLDOWN(), .FAB_DPPULLDOWN(), 
        .FAB_DRVVBUS(), .FAB_IDPULLUP(), .FAB_OPMODE({nc46, nc47}), 
        .FAB_SUSPENDM(), .FAB_TERMSEL(), .FAB_TXVALID(), .FAB_VCONTROL({
        nc48, nc49, nc50, nc51}), .FAB_VCONTROLLOADM(), .FAB_XCVRSEL({
        nc52, nc53}), .FAB_XDATAOUT({nc54, nc55, nc56, nc57, nc58, 
        nc59, nc60, nc61}), .FACC_GLMUX_SEL(), .FIC32_0_MASTER({nc62, 
        nc63}), .FIC32_1_MASTER({nc64, nc65}), .FPGA_RESET_N(
        FPGA_RESET_N), .GTX_CLK(), .H2F_INTERRUPT({nc66, nc67, nc68, 
        nc69, nc70, nc71, nc72, nc73, nc74, nc75, nc76, nc77, nc78, 
        nc79, nc80, nc81}), .H2F_NMI(), .H2FCALIB(), 
        .I2C0_SCL_MGPIO31B_H2F_A(), .I2C0_SCL_MGPIO31B_H2F_B(), 
        .I2C0_SDA_MGPIO30B_H2F_A(), .I2C0_SDA_MGPIO30B_H2F_B(), 
        .I2C1_SCL_MGPIO1A_H2F_A(), .I2C1_SCL_MGPIO1A_H2F_B(), 
        .I2C1_SDA_MGPIO0A_H2F_A(), .I2C1_SDA_MGPIO0A_H2F_B(), .MDCF(), 
        .MDOENF(), .MDOF(), .MMUART0_CTS_MGPIO19B_H2F_A(), 
        .MMUART0_CTS_MGPIO19B_H2F_B(), .MMUART0_DCD_MGPIO22B_H2F_A(), 
        .MMUART0_DCD_MGPIO22B_H2F_B(), .MMUART0_DSR_MGPIO20B_H2F_A(), 
        .MMUART0_DSR_MGPIO20B_H2F_B(), .MMUART0_DTR_MGPIO18B_H2F_A(), 
        .MMUART0_DTR_MGPIO18B_H2F_B(), .MMUART0_RI_MGPIO21B_H2F_A(), 
        .MMUART0_RI_MGPIO21B_H2F_B(), .MMUART0_RTS_MGPIO17B_H2F_A(), 
        .MMUART0_RTS_MGPIO17B_H2F_B(), .MMUART0_RXD_MGPIO28B_H2F_A(), 
        .MMUART0_RXD_MGPIO28B_H2F_B(), .MMUART0_SCK_MGPIO29B_H2F_A(), 
        .MMUART0_SCK_MGPIO29B_H2F_B(), .MMUART0_TXD_MGPIO27B_H2F_A(), 
        .MMUART0_TXD_MGPIO27B_H2F_B(), .MMUART1_DTR_MGPIO12B_H2F_A(), 
        .MMUART1_RTS_MGPIO11B_H2F_A(), .MMUART1_RTS_MGPIO11B_H2F_B(), 
        .MMUART1_RXD_MGPIO26B_H2F_A(), .MMUART1_RXD_MGPIO26B_H2F_B(), 
        .MMUART1_SCK_MGPIO25B_H2F_A(), .MMUART1_SCK_MGPIO25B_H2F_B(), 
        .MMUART1_TXD_MGPIO24B_H2F_A(), .MMUART1_TXD_MGPIO24B_H2F_B(), 
        .MPLL_LOCK(), .PER2_FABRIC_PADDR({nc82, nc83, nc84, nc85, nc86, 
        nc87, nc88, nc89, nc90, nc91, nc92, nc93, nc94, nc95}), 
        .PER2_FABRIC_PENABLE(), .PER2_FABRIC_PSEL(), 
        .PER2_FABRIC_PWDATA({nc96, nc97, nc98, nc99, nc100, nc101, 
        nc102, nc103, nc104, nc105, nc106, nc107, nc108, nc109, nc110, 
        nc111, nc112, nc113, nc114, nc115, nc116, nc117, nc118, nc119, 
        nc120, nc121, nc122, nc123, nc124, nc125, nc126, nc127}), 
        .PER2_FABRIC_PWRITE(), .RTC_MATCH(), .SLEEPDEEP(), 
        .SLEEPHOLDACK(), .SLEEPING(), .SMBALERT_NO0(), .SMBALERT_NO1(), 
        .SMBSUS_NO0(), .SMBSUS_NO1(), .SPI0_CLK_OUT(), 
        .SPI0_SDI_MGPIO5A_H2F_A(), .SPI0_SDI_MGPIO5A_H2F_B(), 
        .SPI0_SDO_MGPIO6A_H2F_A(), .SPI0_SDO_MGPIO6A_H2F_B(), 
        .SPI0_SS0_MGPIO7A_H2F_A(), .SPI0_SS0_MGPIO7A_H2F_B(), 
        .SPI0_SS1_MGPIO8A_H2F_A(), .SPI0_SS1_MGPIO8A_H2F_B(), 
        .SPI0_SS2_MGPIO9A_H2F_A(), .SPI0_SS2_MGPIO9A_H2F_B(), 
        .SPI0_SS3_MGPIO10A_H2F_A(), .SPI0_SS3_MGPIO10A_H2F_B(), 
        .SPI0_SS4_MGPIO19A_H2F_A(), .SPI0_SS5_MGPIO20A_H2F_A(), 
        .SPI0_SS6_MGPIO21A_H2F_A(), .SPI0_SS7_MGPIO22A_H2F_A(), 
        .SPI1_CLK_OUT(), .SPI1_SDI_MGPIO11A_H2F_A(), 
        .SPI1_SDI_MGPIO11A_H2F_B(), .SPI1_SDO_MGPIO12A_H2F_A(), 
        .SPI1_SDO_MGPIO12A_H2F_B(), .SPI1_SS0_MGPIO13A_H2F_A(), 
        .SPI1_SS0_MGPIO13A_H2F_B(), .SPI1_SS1_MGPIO14A_H2F_A(), 
        .SPI1_SS1_MGPIO14A_H2F_B(), .SPI1_SS2_MGPIO15A_H2F_A(), 
        .SPI1_SS2_MGPIO15A_H2F_B(), .SPI1_SS3_MGPIO16A_H2F_A(), 
        .SPI1_SS3_MGPIO16A_H2F_B(), .SPI1_SS4_MGPIO17A_H2F_A(), 
        .SPI1_SS5_MGPIO18A_H2F_A(), .SPI1_SS6_MGPIO23A_H2F_A(), 
        .SPI1_SS7_MGPIO24A_H2F_A(), .TCGF({nc128, nc129, nc130, nc131, 
        nc132, nc133, nc134, nc135, nc136, nc137}), .TRACECLK(), 
        .TRACEDATA({nc138, nc139, nc140, nc141}), .TX_CLK(), .TX_ENF(), 
        .TX_ERRF(), .TXCTL_EN_RIF(), .TXD_RIF({nc142, nc143, nc144, 
        nc145}), .TXDF({nc146, nc147, nc148, nc149, nc150, nc151, 
        nc152, nc153}), .TXEV(), .WDOGTIMEOUT(), .F_ARREADY_HREADYOUT1(
        ), .F_AWREADY_HREADYOUT0(), .F_BID({nc154, nc155, nc156, nc157})
        , .F_BRESP_HRESP0({nc158, nc159}), .F_BVALID(), 
        .F_RDATA_HRDATA01({nc160, nc161, nc162, nc163, nc164, nc165, 
        nc166, nc167, nc168, nc169, nc170, nc171, nc172, nc173, nc174, 
        nc175, nc176, nc177, nc178, nc179, nc180, nc181, nc182, nc183, 
        nc184, nc185, nc186, nc187, nc188, nc189, nc190, nc191, nc192, 
        nc193, nc194, nc195, nc196, nc197, nc198, nc199, nc200, nc201, 
        nc202, nc203, nc204, nc205, nc206, nc207, nc208, nc209, nc210, 
        nc211, nc212, nc213, nc214, nc215, nc216, nc217, nc218, nc219, 
        nc220, nc221, nc222, nc223}), .F_RID({nc224, nc225, nc226, 
        nc227}), .F_RLAST(), .F_RRESP_HRESP1({nc228, nc229}), 
        .F_RVALID(), .F_WREADY(), .MDDR_FABRIC_PRDATA({nc230, nc231, 
        nc232, nc233, nc234, nc235, nc236, nc237, nc238, nc239, nc240, 
        nc241, nc242, nc243, nc244, nc245}), .MDDR_FABRIC_PREADY(), 
        .MDDR_FABRIC_PSLVERR(), .CAN_RXBUS_F2H_SCP(VCC_net_1), 
        .CAN_TX_EBL_F2H_SCP(VCC_net_1), .CAN_TXBUS_F2H_SCP(VCC_net_1), 
        .COLF(VCC_net_1), .CRSF(VCC_net_1), .F2_DMAREADY({VCC_net_1, 
        VCC_net_1}), .F2H_INTERRUPT({GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1}), .F2HCALIB(VCC_net_1), 
        .F_DMAREADY({VCC_net_1, VCC_net_1}), .F_FM0_ADDR({GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1}), .F_FM0_ENABLE(GND_net_1), .F_FM0_MASTLOCK(
        GND_net_1), .F_FM0_READY(VCC_net_1), .F_FM0_SEL(GND_net_1), 
        .F_FM0_SIZE({GND_net_1, GND_net_1}), .F_FM0_TRANS1(GND_net_1), 
        .F_FM0_WDATA({GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1}), .F_FM0_WRITE(GND_net_1), 
        .F_HM0_RDATA({hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[31], 
        hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[30], 
        hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[29], 
        hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[28], 
        hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[27], 
        hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[26], 
        hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[25], 
        hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[24], 
        hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[23], 
        hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[22], 
        hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[21], 
        hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[20], 
        hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[19], 
        hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[18], 
        hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[17], 
        hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[16], 
        hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[15], 
        hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[14], 
        hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[13], 
        hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[12], 
        hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[11], 
        hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[10], 
        hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[9], 
        hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[8], 
        hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[7], 
        hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[6], 
        hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[5], 
        hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[4], 
        hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[3], 
        hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[2], 
        hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[1], 
        hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[0]}), .F_HM0_READY(
        N_676_i_0), .F_HM0_RESP(GND_net_1), .FAB_AVALID(VCC_net_1), 
        .FAB_HOSTDISCON(VCC_net_1), .FAB_IDDIG(VCC_net_1), 
        .FAB_LINESTATE({VCC_net_1, VCC_net_1}), .FAB_M3_RESET_N(
        VCC_net_1), .FAB_PLL_LOCK(FCCC_0_LOCK), .FAB_RXACTIVE(
        VCC_net_1), .FAB_RXERROR(VCC_net_1), .FAB_RXVALID(VCC_net_1), 
        .FAB_RXVALIDH(GND_net_1), .FAB_SESSEND(VCC_net_1), 
        .FAB_TXREADY(VCC_net_1), .FAB_VBUSVALID(VCC_net_1), 
        .FAB_VSTATUS({VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1}), .FAB_XDATAIN({
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1}), .GTX_CLKPF(VCC_net_1), 
        .I2C0_BCLK(VCC_net_1), .I2C0_SCL_F2H_SCP(VCC_net_1), 
        .I2C0_SDA_F2H_SCP(VCC_net_1), .I2C1_BCLK(VCC_net_1), 
        .I2C1_SCL_F2H_SCP(VCC_net_1), .I2C1_SDA_F2H_SCP(VCC_net_1), 
        .MDIF(VCC_net_1), .MGPIO0A_F2H_GPIN(VCC_net_1), 
        .MGPIO10A_F2H_GPIN(VCC_net_1), .MGPIO11A_F2H_GPIN(VCC_net_1), 
        .MGPIO11B_F2H_GPIN(VCC_net_1), .MGPIO12A_F2H_GPIN(VCC_net_1), 
        .MGPIO13A_F2H_GPIN(VCC_net_1), .MGPIO14A_F2H_GPIN(VCC_net_1), 
        .MGPIO15A_F2H_GPIN(VCC_net_1), .MGPIO16A_F2H_GPIN(VCC_net_1), 
        .MGPIO17B_F2H_GPIN(VCC_net_1), .MGPIO18B_F2H_GPIN(VCC_net_1), 
        .MGPIO19B_F2H_GPIN(VCC_net_1), .MGPIO1A_F2H_GPIN(VCC_net_1), 
        .MGPIO20B_F2H_GPIN(VCC_net_1), .MGPIO21B_F2H_GPIN(VCC_net_1), 
        .MGPIO22B_F2H_GPIN(VCC_net_1), .MGPIO24B_F2H_GPIN(VCC_net_1), 
        .MGPIO25B_F2H_GPIN(VCC_net_1), .MGPIO26B_F2H_GPIN(VCC_net_1), 
        .MGPIO27B_F2H_GPIN(VCC_net_1), .MGPIO28B_F2H_GPIN(VCC_net_1), 
        .MGPIO29B_F2H_GPIN(VCC_net_1), .MGPIO2A_F2H_GPIN(VCC_net_1), 
        .MGPIO30B_F2H_GPIN(VCC_net_1), .MGPIO31B_F2H_GPIN(VCC_net_1), 
        .MGPIO3A_F2H_GPIN(VCC_net_1), .MGPIO4A_F2H_GPIN(VCC_net_1), 
        .MGPIO5A_F2H_GPIN(VCC_net_1), .MGPIO6A_F2H_GPIN(VCC_net_1), 
        .MGPIO7A_F2H_GPIN(VCC_net_1), .MGPIO8A_F2H_GPIN(VCC_net_1), 
        .MGPIO9A_F2H_GPIN(VCC_net_1), .MMUART0_CTS_F2H_SCP(VCC_net_1), 
        .MMUART0_DCD_F2H_SCP(VCC_net_1), .MMUART0_DSR_F2H_SCP(
        VCC_net_1), .MMUART0_DTR_F2H_SCP(VCC_net_1), 
        .MMUART0_RI_F2H_SCP(VCC_net_1), .MMUART0_RTS_F2H_SCP(VCC_net_1)
        , .MMUART0_RXD_F2H_SCP(VCC_net_1), .MMUART0_SCK_F2H_SCP(
        VCC_net_1), .MMUART0_TXD_F2H_SCP(VCC_net_1), 
        .MMUART1_CTS_F2H_SCP(VCC_net_1), .MMUART1_DCD_F2H_SCP(
        VCC_net_1), .MMUART1_DSR_F2H_SCP(VCC_net_1), 
        .MMUART1_RI_F2H_SCP(VCC_net_1), .MMUART1_RTS_F2H_SCP(VCC_net_1)
        , .MMUART1_RXD_F2H_SCP(VCC_net_1), .MMUART1_SCK_F2H_SCP(
        VCC_net_1), .MMUART1_TXD_F2H_SCP(VCC_net_1), 
        .PER2_FABRIC_PRDATA({VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1}), 
        .PER2_FABRIC_PREADY(VCC_net_1), .PER2_FABRIC_PSLVERR(VCC_net_1)
        , .RCGF({VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1}), 
        .RX_CLKPF(VCC_net_1), .RX_DVF(VCC_net_1), .RX_ERRF(VCC_net_1), 
        .RX_EV(VCC_net_1), .RXDF({VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1}), 
        .SLEEPHOLDREQ(GND_net_1), .SMBALERT_NI0(VCC_net_1), 
        .SMBALERT_NI1(VCC_net_1), .SMBSUS_NI0(VCC_net_1), .SMBSUS_NI1(
        VCC_net_1), .SPI0_CLK_IN(VCC_net_1), .SPI0_SDI_F2H_SCP(
        VCC_net_1), .SPI0_SDO_F2H_SCP(VCC_net_1), .SPI0_SS0_F2H_SCP(
        VCC_net_1), .SPI0_SS1_F2H_SCP(VCC_net_1), .SPI0_SS2_F2H_SCP(
        VCC_net_1), .SPI0_SS3_F2H_SCP(VCC_net_1), .SPI1_CLK_IN(
        VCC_net_1), .SPI1_SDI_F2H_SCP(VCC_net_1), .SPI1_SDO_F2H_SCP(
        VCC_net_1), .SPI1_SS0_F2H_SCP(VCC_net_1), .SPI1_SS1_F2H_SCP(
        VCC_net_1), .SPI1_SS2_F2H_SCP(VCC_net_1), .SPI1_SS3_F2H_SCP(
        VCC_net_1), .TX_CLKPF(VCC_net_1), .USER_MSS_GPIO_RESET_N(
        VCC_net_1), .USER_MSS_RESET_N(VCC_net_1), .XCLK_FAB(VCC_net_1), 
        .CLK_BASE(FCCC_0_GL1), .CLK_MDDR_APB(VCC_net_1), 
        .F_ARADDR_HADDR1({VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1}), .F_ARBURST_HTRANS1({
        GND_net_1, GND_net_1}), .F_ARID_HSEL1({GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1}), .F_ARLEN_HBURST1({GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1}), .F_ARLOCK_HMASTLOCK1({GND_net_1, 
        GND_net_1}), .F_ARSIZE_HSIZE1({GND_net_1, GND_net_1}), 
        .F_ARVALID_HWRITE1(GND_net_1), .F_AWADDR_HADDR0({VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1}), .F_AWBURST_HTRANS0({GND_net_1, GND_net_1}), 
        .F_AWID_HSEL0({GND_net_1, GND_net_1, GND_net_1, GND_net_1}), 
        .F_AWLEN_HBURST0({GND_net_1, GND_net_1, GND_net_1, GND_net_1}), 
        .F_AWLOCK_HMASTLOCK0({GND_net_1, GND_net_1}), .F_AWSIZE_HSIZE0({
        GND_net_1, GND_net_1}), .F_AWVALID_HWRITE0(GND_net_1), 
        .F_BREADY(GND_net_1), .F_RMW_AXI(GND_net_1), .F_RREADY(
        GND_net_1), .F_WDATA_HWDATA01({VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1}), .F_WID_HREADY01({GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1}), .F_WLAST(GND_net_1), .F_WSTRB({GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1}), .F_WVALID(GND_net_1), 
        .FPGA_MDDR_ARESET_N(VCC_net_1), .MDDR_FABRIC_PADDR({VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1}), .MDDR_FABRIC_PENABLE(
        VCC_net_1), .MDDR_FABRIC_PSEL(VCC_net_1), .MDDR_FABRIC_PWDATA({
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1}), .MDDR_FABRIC_PWRITE(VCC_net_1), .PRESET_N(
        GND_net_1), .CAN_RXBUS_USBA_DATA1_MGPIO3A_IN(GND_net_1), 
        .CAN_TX_EBL_USBA_DATA2_MGPIO4A_IN(GND_net_1), 
        .CAN_TXBUS_USBA_DATA0_MGPIO2A_IN(GND_net_1), .DM_IN({GND_net_1, 
        GND_net_1, GND_net_1}), .DRAM_DQ_IN({GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1}), .DRAM_DQS_IN({GND_net_1, GND_net_1, GND_net_1}), 
        .DRAM_FIFO_WE_IN({GND_net_1, GND_net_1}), 
        .I2C0_SCL_USBC_DATA1_MGPIO31B_IN(GND_net_1), 
        .I2C0_SDA_USBC_DATA0_MGPIO30B_IN(GND_net_1), 
        .I2C1_SCL_USBA_DATA4_MGPIO1A_IN(GND_net_1), 
        .I2C1_SDA_USBA_DATA3_MGPIO0A_IN(GND_net_1), 
        .MMUART0_CTS_USBC_DATA7_MGPIO19B_IN(GND_net_1), 
        .MMUART0_DCD_MGPIO22B_IN(GND_net_1), .MMUART0_DSR_MGPIO20B_IN(
        GND_net_1), .MMUART0_DTR_USBC_DATA6_MGPIO18B_IN(GND_net_1), 
        .MMUART0_RI_MGPIO21B_IN(GND_net_1), 
        .MMUART0_RTS_USBC_DATA5_MGPIO17B_IN(GND_net_1), 
        .MMUART0_RXD_USBC_STP_MGPIO28B_IN(MMUART_0_RXD_PAD_Y), 
        .MMUART0_SCK_USBC_NXT_MGPIO29B_IN(GND_net_1), 
        .MMUART0_TXD_USBC_DIR_MGPIO27B_IN(GND_net_1), 
        .MMUART1_RXD_USBC_DATA3_MGPIO26B_IN(GND_net_1), 
        .MMUART1_SCK_USBC_DATA4_MGPIO25B_IN(GND_net_1), 
        .MMUART1_TXD_USBC_DATA2_MGPIO24B_IN(GND_net_1), 
        .RGMII_GTX_CLK_RMII_CLK_USBB_XCLK_IN(GND_net_1), 
        .RGMII_MDC_RMII_MDC_IN(GND_net_1), 
        .RGMII_MDIO_RMII_MDIO_USBB_DATA7_IN(GND_net_1), 
        .RGMII_RX_CLK_IN(GND_net_1), 
        .RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_IN(GND_net_1), 
        .RGMII_RXD0_RMII_RXD0_USBB_DATA0_IN(GND_net_1), 
        .RGMII_RXD1_RMII_RXD1_USBB_DATA1_IN(GND_net_1), 
        .RGMII_RXD2_RMII_RX_ER_USBB_DATA3_IN(GND_net_1), 
        .RGMII_RXD3_USBB_DATA4_IN(GND_net_1), .RGMII_TX_CLK_IN(
        GND_net_1), .RGMII_TX_CTL_RMII_TX_EN_USBB_NXT_IN(GND_net_1), 
        .RGMII_TXD0_RMII_TXD0_USBB_DIR_IN(GND_net_1), 
        .RGMII_TXD1_RMII_TXD1_USBB_STP_IN(GND_net_1), 
        .RGMII_TXD2_USBB_DATA5_IN(GND_net_1), 
        .RGMII_TXD3_USBB_DATA6_IN(GND_net_1), .SPI0_SCK_USBA_XCLK_IN(
        GND_net_1), .SPI0_SDI_USBA_DIR_MGPIO5A_IN(GND_net_1), 
        .SPI0_SDO_USBA_STP_MGPIO6A_IN(GND_net_1), 
        .SPI0_SS0_USBA_NXT_MGPIO7A_IN(GND_net_1), 
        .SPI0_SS1_USBA_DATA5_MGPIO8A_IN(GND_net_1), 
        .SPI0_SS2_USBA_DATA6_MGPIO9A_IN(GND_net_1), 
        .SPI0_SS3_USBA_DATA7_MGPIO10A_IN(GND_net_1), .SPI1_SCK_IN(
        GND_net_1), .SPI1_SDI_MGPIO11A_IN(GND_net_1), 
        .SPI1_SDO_MGPIO12A_IN(GND_net_1), .SPI1_SS0_MGPIO13A_IN(
        GND_net_1), .SPI1_SS1_MGPIO14A_IN(GND_net_1), 
        .SPI1_SS2_MGPIO15A_IN(GND_net_1), .SPI1_SS3_MGPIO16A_IN(
        GND_net_1), .SPI1_SS4_MGPIO17A_IN(GND_net_1), 
        .SPI1_SS5_MGPIO18A_IN(GND_net_1), .SPI1_SS6_MGPIO23A_IN(
        GND_net_1), .SPI1_SS7_MGPIO24A_IN(GND_net_1), .USBC_XCLK_IN(
        GND_net_1), .CAN_RXBUS_USBA_DATA1_MGPIO3A_OUT(), 
        .CAN_TX_EBL_USBA_DATA2_MGPIO4A_OUT(), 
        .CAN_TXBUS_USBA_DATA0_MGPIO2A_OUT(), .DRAM_ADDR({nc246, nc247, 
        nc248, nc249, nc250, nc251, nc252, nc253, nc254, nc255, nc256, 
        nc257, nc258, nc259, nc260, nc261}), .DRAM_BA({nc262, nc263, 
        nc264}), .DRAM_CASN(), .DRAM_CKE(), .DRAM_CLK(), .DRAM_CSN(), 
        .DRAM_DM_RDQS_OUT({nc265, nc266, nc267}), .DRAM_DQ_OUT({nc268, 
        nc269, nc270, nc271, nc272, nc273, nc274, nc275, nc276, nc277, 
        nc278, nc279, nc280, nc281, nc282, nc283, nc284, nc285}), 
        .DRAM_DQS_OUT({nc286, nc287, nc288}), .DRAM_FIFO_WE_OUT({nc289, 
        nc290}), .DRAM_ODT(), .DRAM_RASN(), .DRAM_RSTN(), .DRAM_WEN(), 
        .I2C0_SCL_USBC_DATA1_MGPIO31B_OUT(), 
        .I2C0_SDA_USBC_DATA0_MGPIO30B_OUT(), 
        .I2C1_SCL_USBA_DATA4_MGPIO1A_OUT(), 
        .I2C1_SDA_USBA_DATA3_MGPIO0A_OUT(), 
        .MMUART0_CTS_USBC_DATA7_MGPIO19B_OUT(), 
        .MMUART0_DCD_MGPIO22B_OUT(), .MMUART0_DSR_MGPIO20B_OUT(), 
        .MMUART0_DTR_USBC_DATA6_MGPIO18B_OUT(), 
        .MMUART0_RI_MGPIO21B_OUT(), 
        .MMUART0_RTS_USBC_DATA5_MGPIO17B_OUT(), 
        .MMUART0_RXD_USBC_STP_MGPIO28B_OUT(), 
        .MMUART0_SCK_USBC_NXT_MGPIO29B_OUT(), 
        .MMUART0_TXD_USBC_DIR_MGPIO27B_OUT(
        MSS_ADLIB_INST_MMUART0_TXD_USBC_DIR_MGPIO27B_OUT), 
        .MMUART1_RXD_USBC_DATA3_MGPIO26B_OUT(), 
        .MMUART1_SCK_USBC_DATA4_MGPIO25B_OUT(), 
        .MMUART1_TXD_USBC_DATA2_MGPIO24B_OUT(), 
        .RGMII_GTX_CLK_RMII_CLK_USBB_XCLK_OUT(), 
        .RGMII_MDC_RMII_MDC_OUT(), 
        .RGMII_MDIO_RMII_MDIO_USBB_DATA7_OUT(), .RGMII_RX_CLK_OUT(), 
        .RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_OUT(), 
        .RGMII_RXD0_RMII_RXD0_USBB_DATA0_OUT(), 
        .RGMII_RXD1_RMII_RXD1_USBB_DATA1_OUT(), 
        .RGMII_RXD2_RMII_RX_ER_USBB_DATA3_OUT(), 
        .RGMII_RXD3_USBB_DATA4_OUT(), .RGMII_TX_CLK_OUT(), 
        .RGMII_TX_CTL_RMII_TX_EN_USBB_NXT_OUT(), 
        .RGMII_TXD0_RMII_TXD0_USBB_DIR_OUT(), 
        .RGMII_TXD1_RMII_TXD1_USBB_STP_OUT(), 
        .RGMII_TXD2_USBB_DATA5_OUT(), .RGMII_TXD3_USBB_DATA6_OUT(), 
        .SPI0_SCK_USBA_XCLK_OUT(), .SPI0_SDI_USBA_DIR_MGPIO5A_OUT(), 
        .SPI0_SDO_USBA_STP_MGPIO6A_OUT(), 
        .SPI0_SS0_USBA_NXT_MGPIO7A_OUT(), 
        .SPI0_SS1_USBA_DATA5_MGPIO8A_OUT(), 
        .SPI0_SS2_USBA_DATA6_MGPIO9A_OUT(), 
        .SPI0_SS3_USBA_DATA7_MGPIO10A_OUT(), .SPI1_SCK_OUT(), 
        .SPI1_SDI_MGPIO11A_OUT(), .SPI1_SDO_MGPIO12A_OUT(), 
        .SPI1_SS0_MGPIO13A_OUT(), .SPI1_SS1_MGPIO14A_OUT(), 
        .SPI1_SS2_MGPIO15A_OUT(), .SPI1_SS3_MGPIO16A_OUT(), 
        .SPI1_SS4_MGPIO17A_OUT(), .SPI1_SS5_MGPIO18A_OUT(), 
        .SPI1_SS6_MGPIO23A_OUT(), .SPI1_SS7_MGPIO24A_OUT(), 
        .USBC_XCLK_OUT(), .CAN_RXBUS_USBA_DATA1_MGPIO3A_OE(), 
        .CAN_TX_EBL_USBA_DATA2_MGPIO4A_OE(), 
        .CAN_TXBUS_USBA_DATA0_MGPIO2A_OE(), .DM_OE({nc291, nc292, 
        nc293}), .DRAM_DQ_OE({nc294, nc295, nc296, nc297, nc298, nc299, 
        nc300, nc301, nc302, nc303, nc304, nc305, nc306, nc307, nc308, 
        nc309, nc310, nc311}), .DRAM_DQS_OE({nc312, nc313, nc314}), 
        .I2C0_SCL_USBC_DATA1_MGPIO31B_OE(), 
        .I2C0_SDA_USBC_DATA0_MGPIO30B_OE(), 
        .I2C1_SCL_USBA_DATA4_MGPIO1A_OE(), 
        .I2C1_SDA_USBA_DATA3_MGPIO0A_OE(), 
        .MMUART0_CTS_USBC_DATA7_MGPIO19B_OE(), 
        .MMUART0_DCD_MGPIO22B_OE(), .MMUART0_DSR_MGPIO20B_OE(), 
        .MMUART0_DTR_USBC_DATA6_MGPIO18B_OE(), .MMUART0_RI_MGPIO21B_OE(
        ), .MMUART0_RTS_USBC_DATA5_MGPIO17B_OE(), 
        .MMUART0_RXD_USBC_STP_MGPIO28B_OE(), 
        .MMUART0_SCK_USBC_NXT_MGPIO29B_OE(), 
        .MMUART0_TXD_USBC_DIR_MGPIO27B_OE(
        MSS_ADLIB_INST_MMUART0_TXD_USBC_DIR_MGPIO27B_OE), 
        .MMUART1_RXD_USBC_DATA3_MGPIO26B_OE(), 
        .MMUART1_SCK_USBC_DATA4_MGPIO25B_OE(), 
        .MMUART1_TXD_USBC_DATA2_MGPIO24B_OE(), 
        .RGMII_GTX_CLK_RMII_CLK_USBB_XCLK_OE(), .RGMII_MDC_RMII_MDC_OE(
        ), .RGMII_MDIO_RMII_MDIO_USBB_DATA7_OE(), .RGMII_RX_CLK_OE(), 
        .RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_OE(), 
        .RGMII_RXD0_RMII_RXD0_USBB_DATA0_OE(), 
        .RGMII_RXD1_RMII_RXD1_USBB_DATA1_OE(), 
        .RGMII_RXD2_RMII_RX_ER_USBB_DATA3_OE(), 
        .RGMII_RXD3_USBB_DATA4_OE(), .RGMII_TX_CLK_OE(), 
        .RGMII_TX_CTL_RMII_TX_EN_USBB_NXT_OE(), 
        .RGMII_TXD0_RMII_TXD0_USBB_DIR_OE(), 
        .RGMII_TXD1_RMII_TXD1_USBB_STP_OE(), .RGMII_TXD2_USBB_DATA5_OE(
        ), .RGMII_TXD3_USBB_DATA6_OE(), .SPI0_SCK_USBA_XCLK_OE(), 
        .SPI0_SDI_USBA_DIR_MGPIO5A_OE(), .SPI0_SDO_USBA_STP_MGPIO6A_OE(
        ), .SPI0_SS0_USBA_NXT_MGPIO7A_OE(), 
        .SPI0_SS1_USBA_DATA5_MGPIO8A_OE(), 
        .SPI0_SS2_USBA_DATA6_MGPIO9A_OE(), 
        .SPI0_SS3_USBA_DATA7_MGPIO10A_OE(), .SPI1_SCK_OE(), 
        .SPI1_SDI_MGPIO11A_OE(), .SPI1_SDO_MGPIO12A_OE(), 
        .SPI1_SS0_MGPIO13A_OE(), .SPI1_SS1_MGPIO14A_OE(), 
        .SPI1_SS2_MGPIO15A_OE(), .SPI1_SS3_MGPIO16A_OE(), 
        .SPI1_SS4_MGPIO17A_OE(), .SPI1_SS5_MGPIO18A_OE(), 
        .SPI1_SS6_MGPIO23A_OE(), .SPI1_SS7_MGPIO24A_OE(), 
        .USBC_XCLK_OE());
    GND GND (.Y(GND_net_1));
    TRIBUFF MMUART_0_TXD_PAD (.D(
        MSS_ADLIB_INST_MMUART0_TXD_USBC_DIR_MGPIO27B_OUT), .E(
        MSS_ADLIB_INST_MMUART0_TXD_USBC_DIR_MGPIO27B_OE), .PAD(
        MMUART_0_TXD));
    
endmodule


module hello_regs_FCCC_0_FCCC(
       FCCC_0_GL1,
       FCCC_0_LOCK,
       OSC_0_RCOSC_25_50MHZ_CCC_OUT_RCOSC_25_50MHZ_CCC
    );
output FCCC_0_GL1;
output FCCC_0_LOCK;
input  OSC_0_RCOSC_25_50MHZ_CCC_OUT_RCOSC_25_50MHZ_CCC;

    wire GL1_net, VCC_net_1, GND_net_1;
    
    CLKINT GL1_INST (.A(GL1_net), .Y(FCCC_0_GL1));
    VCC VCC (.Y(VCC_net_1));
    GND GND (.Y(GND_net_1));
    CCC #( .INIT(210'h0000007FB8000044D64000318C6307C6318C61EC0404040400301)
        , .VCOFREQUENCY(800.0) )  CCC_INST (.Y0(), .Y1(), .Y2(), .Y3(), 
        .PRDATA({nc0, nc1, nc2, nc3, nc4, nc5, nc6, nc7}), .LOCK(
        FCCC_0_LOCK), .BUSY(), .CLK0(VCC_net_1), .CLK1(VCC_net_1), 
        .CLK2(VCC_net_1), .CLK3(VCC_net_1), .NGMUX0_SEL(GND_net_1), 
        .NGMUX1_SEL(GND_net_1), .NGMUX2_SEL(GND_net_1), .NGMUX3_SEL(
        GND_net_1), .NGMUX0_HOLD_N(VCC_net_1), .NGMUX1_HOLD_N(
        VCC_net_1), .NGMUX2_HOLD_N(VCC_net_1), .NGMUX3_HOLD_N(
        VCC_net_1), .NGMUX0_ARST_N(VCC_net_1), .NGMUX1_ARST_N(
        VCC_net_1), .NGMUX2_ARST_N(VCC_net_1), .NGMUX3_ARST_N(
        VCC_net_1), .PLL_BYPASS_N(VCC_net_1), .PLL_ARST_N(VCC_net_1), 
        .PLL_POWERDOWN_N(VCC_net_1), .GPD0_ARST_N(VCC_net_1), 
        .GPD1_ARST_N(VCC_net_1), .GPD2_ARST_N(VCC_net_1), .GPD3_ARST_N(
        VCC_net_1), .PRESET_N(GND_net_1), .PCLK(VCC_net_1), .PSEL(
        VCC_net_1), .PENABLE(VCC_net_1), .PWRITE(VCC_net_1), .PADDR({
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1}), .PWDATA({VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1}), 
        .CLK0_PAD(GND_net_1), .CLK1_PAD(GND_net_1), .CLK2_PAD(
        GND_net_1), .CLK3_PAD(GND_net_1), .GL0(), .GL1(GL1_net), .GL2()
        , .GL3(), .RCOSC_25_50MHZ(
        OSC_0_RCOSC_25_50MHZ_CCC_OUT_RCOSC_25_50MHZ_CCC), .RCOSC_1MHZ(
        GND_net_1), .XTLOSC(GND_net_1));
    
endmodule


module reg16x8(
       CoreAPB3_0_APBmslave5_PRDATA,
       CoreAPB3_0_APBmslave4_PWDATA,
       CoreAPB3_0_APBmslave4_PADDR,
       mem_8__2_i_0_0_a2,
       mem_0__2_i_0_0_a2,
       PRDATA_0_iv_0_0_a2_1,
       MSS_RESET_N_M2F_c,
       FCCC_0_GL1,
       rd_enable,
       CoreAPB3_0_APBmslave4_PENABLE,
       CoreAPB3_0_APBmslave4_PWRITE
    );
output [7:0] CoreAPB3_0_APBmslave5_PRDATA;
input  [7:0] CoreAPB3_0_APBmslave4_PWDATA;
input  [5:2] CoreAPB3_0_APBmslave4_PADDR;
output [2:2] mem_8__2_i_0_0_a2;
output [0:0] mem_0__2_i_0_0_a2;
input  [3:3] PRDATA_0_iv_0_0_a2_1;
input  MSS_RESET_N_M2F_c;
input  FCCC_0_GL1;
input  rd_enable;
input  CoreAPB3_0_APBmslave4_PENABLE;
input  CoreAPB3_0_APBmslave4_PWRITE;

    wire un1_data_out8_121_net_1, un1_data_out8_121_i, 
        un1_data_out8_25_net_1, un1_data_out8_25_i, 
        un1_data_out8_9_net_1, un1_data_out8_9_i, 
        un1_data_out8_80_net_1, un1_data_out8_80_i, 
        un1_data_out8_27_net_1, un1_data_out8_27_i, 
        un1_data_out8_11_net_1, un1_data_out8_11_i, 
        un1_data_out8_81_net_1, un1_data_out8_81_i, 
        un1_data_out8_57_net_1, un1_data_out8_57_i, 
        un1_data_out8_112_net_1, un1_data_out8_112_i, 
        un1_data_out8_104_net_1, un1_data_out8_104_i, 
        un1_data_out8_16_net_1, un1_data_out8_16_i, 
        un1_data_out8_88_net_1, un1_data_out8_88_i, 
        un1_data_out8_97_net_1, un1_data_out8_97_i, 
        un1_data_out8_72_net_1, un1_data_out8_72_i, 
        un1_data_out8_7_net_1, un1_data_out8_7_i, 
        un1_data_out8_124_net_1, un1_data_out8_124_i, 
        un1_data_out8_28_net_1, un1_data_out8_28_i, 
        un1_data_out8_12_net_1, un1_data_out8_12_i, 
        un1_data_out8_net_1, un1_data_out8_i, un1_data_out8_13_net_1, 
        un1_data_out8_13_i, un1_data_out8_82_net_1, un1_data_out8_82_i, 
        un1_data_out8_58_net_1, un1_data_out8_58_i, 
        un1_data_out8_113_net_1, un1_data_out8_113_i, 
        un1_data_out8_105_net_1, un1_data_out8_105_i, 
        un1_data_out8_17_net_1, un1_data_out8_17_i, 
        un1_data_out8_89_net_1, un1_data_out8_89_i, 
        un1_data_out8_98_net_1, un1_data_out8_98_i, 
        un1_data_out8_73_net_1, un1_data_out8_73_i, 
        un1_data_out8_5_net_1, un1_data_out8_5_i, 
        un1_data_out8_126_net_1, un1_data_out8_126_i, 
        un1_data_out8_30_net_1, un1_data_out8_30_i, 
        un1_data_out8_14_net_1, un1_data_out8_14_i, 
        un1_data_out8_2_net_1, un1_data_out8_2_i, 
        un1_data_out8_123_net_1, un1_data_out8_123_i, 
        un1_data_out8_83_net_1, un1_data_out8_83_i, 
        un1_data_out8_59_net_1, un1_data_out8_59_i, 
        un1_data_out8_114_net_1, un1_data_out8_114_i, 
        un1_data_out8_106_net_1, un1_data_out8_106_i, 
        un1_data_out8_18_net_1, un1_data_out8_18_i, 
        un1_data_out8_90_net_1, un1_data_out8_90_i, 
        un1_data_out8_99_net_1, un1_data_out8_99_i, 
        un1_data_out8_74_net_1, un1_data_out8_74_i, 
        un1_data_out8_64_net_1, un1_data_out8_64_i, 
        un1_data_out8_48_net_1, un1_data_out8_48_i, 
        un1_data_out8_32_net_1, un1_data_out8_32_i, 
        un1_data_out8_43_net_1, un1_data_out8_43_i, 
        un1_data_out8_4_net_1, un1_data_out8_4_i, 
        un1_data_out8_125_net_1, un1_data_out8_125_i, 
        un1_data_out8_29_net_1, un1_data_out8_29_i, 
        un1_data_out8_56_net_1, un1_data_out8_56_i, 
        un1_data_out8_115_net_1, un1_data_out8_115_i, 
        un1_data_out8_107_net_1, un1_data_out8_107_i, 
        un1_data_out8_19_net_1, un1_data_out8_19_i, 
        un1_data_out8_91_net_1, un1_data_out8_91_i, 
        un1_data_out8_96_net_1, un1_data_out8_96_i, 
        un1_data_out8_75_net_1, un1_data_out8_75_i, 
        un1_data_out8_66_net_1, un1_data_out8_66_i, 
        un1_data_out8_50_net_1, un1_data_out8_50_i, 
        un1_data_out8_34_net_1, un1_data_out8_34_i, 
        un1_data_out8_41_net_1, un1_data_out8_41_i, 
        un1_data_out8_6_net_1, un1_data_out8_6_i, 
        un1_data_out8_127_net_1, un1_data_out8_127_i, 
        un1_data_out8_31_net_1, un1_data_out8_31_i, 
        un1_data_out8_15_net_1, un1_data_out8_15_i, 
        un1_data_out8_116_net_1, un1_data_out8_116_i, 
        un1_data_out8_108_net_1, un1_data_out8_108_i, 
        un1_data_out8_20_net_1, un1_data_out8_20_i, 
        un1_data_out8_92_net_1, un1_data_out8_92_i, 
        un1_data_out8_101_net_1, un1_data_out8_101_i, 
        un1_data_out8_76_net_1, un1_data_out8_76_i, 
        un1_data_out8_68_net_1, un1_data_out8_68_i, 
        un1_data_out8_52_net_1, un1_data_out8_52_i, 
        un1_data_out8_36_net_1, un1_data_out8_36_i, 
        un1_data_out8_47_net_1, un1_data_out8_47_i, 
        un1_data_out8_65_net_1, un1_data_out8_65_i, 
        un1_data_out8_49_net_1, un1_data_out8_49_i, 
        un1_data_out8_33_net_1, un1_data_out8_33_i, 
        un1_data_out8_40_net_1, un1_data_out8_40_i, 
        un1_data_out8_84_net_1, un1_data_out8_84_i, 
        un1_data_out8_109_net_1, un1_data_out8_109_i, 
        un1_data_out8_21_net_1, un1_data_out8_21_i, 
        un1_data_out8_93_net_1, un1_data_out8_93_i, 
        un1_data_out8_102_net_1, un1_data_out8_102_i, 
        un1_data_out8_77_net_1, un1_data_out8_77_i, 
        un1_data_out8_69_net_1, un1_data_out8_69_i, 
        un1_data_out8_54_net_1, un1_data_out8_54_i, 
        un1_data_out8_38_net_1, un1_data_out8_38_i, 
        un1_data_out8_45_net_1, un1_data_out8_45_i, 
        un1_data_out8_67_net_1, un1_data_out8_67_i, 
        un1_data_out8_51_net_1, un1_data_out8_51_i, 
        un1_data_out8_35_net_1, un1_data_out8_35_i, 
        un1_data_out8_42_net_1, un1_data_out8_42_i, 
        un1_data_out8_85_net_1, un1_data_out8_85_i, 
        un1_data_out8_61_net_1, un1_data_out8_61_i, 
        un1_data_out8_22_net_1, un1_data_out8_22_i, 
        un1_data_out8_94_net_1, un1_data_out8_94_i, 
        un1_data_out8_103_net_1, un1_data_out8_103_i, 
        un1_data_out8_78_net_1, un1_data_out8_78_i, 
        un1_data_out8_70_net_1, un1_data_out8_70_i, 
        un1_data_out8_3_net_1, un1_data_out8_3_i, 
        un1_data_out8_120_net_1, un1_data_out8_120_i, 
        un1_data_out8_24_net_1, un1_data_out8_24_i, 
        un1_data_out8_8_net_1, un1_data_out8_8_i, 
        un1_data_out8_53_net_1, un1_data_out8_53_i, 
        un1_data_out8_37_net_1, un1_data_out8_37_i, 
        un1_data_out8_44_net_1, un1_data_out8_44_i, 
        un1_data_out8_86_net_1, un1_data_out8_86_i, 
        un1_data_out8_62_net_1, un1_data_out8_62_i, 
        un1_data_out8_117_net_1, un1_data_out8_117_i, 
        un1_data_out8_95_net_1, un1_data_out8_95_i, 
        un1_data_out8_100_net_1, un1_data_out8_100_i, 
        un1_data_out8_79_net_1, un1_data_out8_79_i, 
        un1_data_out8_71_net_1, un1_data_out8_71_i, 
        un1_data_out8_1_net_1, un1_data_out8_1_i, 
        un1_data_out8_122_net_1, un1_data_out8_122_i, 
        un1_data_out8_26_net_1, un1_data_out8_26_i, 
        un1_data_out8_10_net_1, un1_data_out8_10_i, 
        un1_data_out8_55_net_1, un1_data_out8_55_i, 
        un1_data_out8_39_net_1, un1_data_out8_39_i, 
        un1_data_out8_46_net_1, un1_data_out8_46_i, 
        un1_data_out8_87_net_1, un1_data_out8_87_i, 
        un1_data_out8_63_net_1, un1_data_out8_63_i, 
        un1_data_out8_118_net_1, un1_data_out8_118_i, 
        un1_data_out8_110_net_1, un1_data_out8_110_i, 
        un1_data_out8_60_net_1, un1_data_out8_60_i, 
        un1_data_out8_119_net_1, un1_data_out8_119_i, 
        un1_data_out8_111_net_1, un1_data_out8_111_i, 
        un1_data_out8_23_net_1, un1_data_out8_23_i, VCC_net_1, N_11, 
        GND_net_1, N_9, N_13, N_7, N_15, N_17, N_19, N_5, 
        un1_data_out8_23_set_net_1, un1_data_out8_247_rs_net_1, 
        \mem_12_rs[7] , \mem_12_[7]_net_1 , un1_data_out8_247_i, 
        mem_12__1_sqmuxa, un1_data_out8_111_set_net_1, 
        un1_data_out8_215_rs_net_1, \mem_13_rs[7] , \mem_13_[7]_net_1 , 
        un1_data_out8_215_i, mem_13__1_sqmuxa, 
        un1_data_out8_119_set_net_1, un1_data_out8_223_rs_net_1, 
        \mem_14_rs[7] , \mem_14_[7]_net_1 , un1_data_out8_223_i, 
        mem_14__1_sqmuxa, un1_data_out8_60_set_net_1, 
        un1_data_out8_254_rs_net_1, \mem_15_rs[7] , \mem_15_[7]_net_1 , 
        un1_data_out8_254_i, mem_15__1_sqmuxa, 
        un1_data_out8_110_set_net_1, un1_data_out8_214_rs_net_1, 
        \mem_13_rs[6] , \mem_13_[6]_net_1 , un1_data_out8_214_i, 
        un1_data_out8_118_set_net_1, un1_data_out8_222_rs_net_1, 
        \mem_14_rs[6] , \mem_14_[6]_net_1 , un1_data_out8_222_i, 
        un1_data_out8_63_set_net_1, un1_data_out8_253_rs_net_1, 
        \mem_15_rs[6] , \mem_15_[6]_net_1 , un1_data_out8_253_i, 
        un1_data_out8_87_set_net_1, un1_data_out8_151_rs_net_1, 
        \mem_0_rs[7] , \mem_0_[7]_net_1 , un1_data_out8_151_i, 
        mem_0__1_sqmuxa, un1_data_out8_46_set_net_1, 
        un1_data_out8_159_rs_net_1, \mem_1_rs[7] , \mem_1_[7]_net_1 , 
        un1_data_out8_159_i, mem_1__1_sqmuxa, 
        un1_data_out8_39_set_net_1, un1_data_out8_167_rs_net_1, 
        \mem_2_rs[7] , \mem_2_[7]_net_1 , un1_data_out8_167_i, 
        mem_2__1_sqmuxa, un1_data_out8_55_set_net_1, 
        un1_data_out8_135_rs_net_1, \mem_3_rs[7] , \mem_3_[7]_net_1 , 
        un1_data_out8_135_i, mem_3__1_sqmuxa, 
        un1_data_out8_10_set_net_1, un1_data_out8_185_rs_net_1, 
        \mem_4_rs[7] , \mem_4_[7]_net_1 , un1_data_out8_185_i, 
        mem_4__1_sqmuxa, un1_data_out8_26_set_net_1, 
        un1_data_out8_201_rs_net_1, \mem_5_rs[7] , \mem_5_[7]_net_1 , 
        un1_data_out8_201_i, mem_5__1_sqmuxa, 
        un1_data_out8_122_set_net_1, un1_data_out8_177_rs_net_1, 
        \mem_6_rs[7] , \mem_6_[7]_net_1 , un1_data_out8_177_i, 
        mem_6__1_sqmuxa, un1_data_out8_1_set_net_1, 
        un1_data_out8_233_rs_net_1, \mem_7_rs[7] , \mem_7_[7]_net_1 , 
        un1_data_out8_233_i, mem_7__1_sqmuxa, 
        un1_data_out8_71_set_net_1, un1_data_out8_188_rs_net_1, 
        \mem_8_rs[7] , \mem_8_[7]_net_1 , un1_data_out8_188_i, 
        mem_8__1_sqmuxa, un1_data_out8_79_set_net_1, 
        un1_data_out8_204_rs_net_1, \mem_9_rs[7] , \mem_9_[7]_net_1 , 
        un1_data_out8_204_i, mem_9__1_sqmuxa, 
        un1_data_out8_100_set_net_1, un1_data_out8_180_rs_net_1, 
        \mem_10_rs[7] , \mem_10_[7]_net_1 , un1_data_out8_180_i, 
        mem_10__1_sqmuxa, un1_data_out8_95_set_net_1, 
        un1_data_out8_236_rs_net_1, \mem_11_rs[7] , \mem_11_[7]_net_1 , 
        un1_data_out8_236_i, mem_11__1_sqmuxa, 
        un1_data_out8_117_set_net_1, un1_data_out8_221_rs_net_1, 
        \mem_14_rs[5] , \mem_14_[5]_net_1 , un1_data_out8_221_i, 
        un1_data_out8_62_set_net_1, un1_data_out8_252_rs_net_1, 
        \mem_15_rs[5] , \mem_15_[5]_net_1 , un1_data_out8_252_i, 
        un1_data_out8_86_set_net_1, un1_data_out8_150_rs_net_1, 
        \mem_0_rs[6] , \mem_0_[6]_net_1 , un1_data_out8_150_i, 
        un1_data_out8_44_set_net_1, un1_data_out8_158_rs_net_1, 
        \mem_1_rs[6] , \mem_1_[6]_net_1 , un1_data_out8_158_i, 
        un1_data_out8_37_set_net_1, un1_data_out8_166_rs_net_1, 
        \mem_2_rs[6] , \mem_2_[6]_net_1 , un1_data_out8_166_i, 
        un1_data_out8_53_set_net_1, un1_data_out8_134_rs_net_1, 
        \mem_3_rs[6] , \mem_3_[6]_net_1 , un1_data_out8_134_i, 
        un1_data_out8_8_set_net_1, un1_data_out8_143_rs_net_1, 
        \mem_4_rs[6] , \mem_4_[6]_net_1 , un1_data_out8_143_i, 
        un1_data_out8_24_set_net_1, un1_data_out8_199_rs_net_1, 
        \mem_5_rs[6] , \mem_5_[6]_net_1 , un1_data_out8_199_i, 
        un1_data_out8_120_set_net_1, un1_data_out8_175_rs_net_1, 
        \mem_6_rs[6] , \mem_6_[6]_net_1 , un1_data_out8_175_i, 
        un1_data_out8_3_set_net_1, un1_data_out8_231_rs_net_1, 
        \mem_7_rs[6] , \mem_7_[6]_net_1 , un1_data_out8_231_i, 
        un1_data_out8_70_set_net_1, un1_data_out8_186_rs_net_1, 
        \mem_8_rs[6] , \mem_8_[6]_net_1 , un1_data_out8_186_i, 
        un1_data_out8_78_set_net_1, un1_data_out8_202_rs_net_1, 
        \mem_9_rs[6] , \mem_9_[6]_net_1 , un1_data_out8_202_i, 
        un1_data_out8_103_set_net_1, un1_data_out8_178_rs_net_1, 
        \mem_10_rs[6] , \mem_10_[6]_net_1 , un1_data_out8_178_i, 
        un1_data_out8_94_set_net_1, un1_data_out8_234_rs_net_1, 
        \mem_11_rs[6] , \mem_11_[6]_net_1 , un1_data_out8_234_i, 
        un1_data_out8_22_set_net_1, un1_data_out8_246_rs_net_1, 
        \mem_12_rs[6] , \mem_12_[6]_net_1 , un1_data_out8_246_i, 
        un1_data_out8_61_set_net_1, un1_data_out8_255_rs_net_1, 
        \mem_15_rs[4] , \mem_15_[4]_net_1 , un1_data_out8_255_i, 
        un1_data_out8_85_set_net_1, un1_data_out8_149_rs_net_1, 
        \mem_0_rs[5] , \mem_0_[5]_net_1 , un1_data_out8_149_i, 
        un1_data_out8_42_set_net_1, un1_data_out8_157_rs_net_1, 
        \mem_1_rs[5] , \mem_1_[5]_net_1 , un1_data_out8_157_i, 
        un1_data_out8_35_set_net_1, un1_data_out8_165_rs_net_1, 
        \mem_2_rs[5] , \mem_2_[5]_net_1 , un1_data_out8_165_i, 
        un1_data_out8_51_set_net_1, un1_data_out8_133_rs_net_1, 
        \mem_3_rs[5] , \mem_3_[5]_net_1 , un1_data_out8_133_i, 
        un1_data_out8_67_set_net_1, un1_data_out8_141_rs_net_1, 
        \mem_4_rs[5] , \mem_4_[5]_net_1 , un1_data_out8_141_i, 
        un1_data_out8_45_set_net_1, un1_data_out8_197_rs_net_1, 
        \mem_5_rs[5] , \mem_5_[5]_net_1 , un1_data_out8_197_i, 
        un1_data_out8_38_set_net_1, un1_data_out8_173_rs_net_1, 
        \mem_6_rs[5] , \mem_6_[5]_net_1 , un1_data_out8_173_i, 
        un1_data_out8_54_set_net_1, un1_data_out8_229_rs_net_1, 
        \mem_7_rs[5] , \mem_7_[5]_net_1 , un1_data_out8_229_i, 
        un1_data_out8_69_set_net_1, un1_data_out8_184_rs_net_1, 
        \mem_8_rs[5] , \mem_8_[5]_net_1 , un1_data_out8_184_i, 
        un1_data_out8_77_set_net_1, un1_data_out8_200_rs_net_1, 
        \mem_9_rs[5] , \mem_9_[5]_net_1 , un1_data_out8_200_i, 
        un1_data_out8_102_set_net_1, un1_data_out8_176_rs_net_1, 
        \mem_10_rs[5] , \mem_10_[5]_net_1 , un1_data_out8_176_i, 
        un1_data_out8_93_set_net_1, un1_data_out8_232_rs_net_1, 
        \mem_11_rs[5] , \mem_11_[5]_net_1 , un1_data_out8_232_i, 
        un1_data_out8_21_set_net_1, un1_data_out8_245_rs_net_1, 
        \mem_12_rs[5] , \mem_12_[5]_net_1 , un1_data_out8_245_i, 
        un1_data_out8_109_set_net_1, un1_data_out8_213_rs_net_1, 
        \mem_13_rs[5] , \mem_13_[5]_net_1 , un1_data_out8_213_i, 
        un1_data_out8_84_set_net_1, un1_data_out8_148_rs_net_1, 
        \mem_0_rs[4] , \mem_0_[4]_net_1 , un1_data_out8_148_i, 
        un1_data_out8_40_set_net_1, un1_data_out8_156_rs_net_1, 
        \mem_1_rs[4] , \mem_1_[4]_net_1 , un1_data_out8_156_i, 
        un1_data_out8_33_set_net_1, un1_data_out8_164_rs_net_1, 
        \mem_2_rs[4] , \mem_2_[4]_net_1 , un1_data_out8_164_i, 
        un1_data_out8_49_set_net_1, un1_data_out8_132_rs_net_1, 
        \mem_3_rs[4] , \mem_3_[4]_net_1 , un1_data_out8_132_i, 
        un1_data_out8_65_set_net_1, un1_data_out8_140_rs_net_1, 
        \mem_4_rs[4] , \mem_4_[4]_net_1 , un1_data_out8_140_i, 
        un1_data_out8_47_set_net_1, un1_data_out8_195_rs_net_1, 
        \mem_5_rs[4] , \mem_5_[4]_net_1 , un1_data_out8_195_i, 
        un1_data_out8_36_set_net_1, un1_data_out8_171_rs_net_1, 
        \mem_6_rs[4] , \mem_6_[4]_net_1 , un1_data_out8_171_i, 
        un1_data_out8_52_set_net_1, un1_data_out8_227_rs_net_1, 
        \mem_7_rs[4] , \mem_7_[4]_net_1 , un1_data_out8_227_i, 
        un1_data_out8_68_set_net_1, un1_data_out8_142_rs_net_1, 
        \mem_8_rs[4] , \mem_8_[4]_net_1 , un1_data_out8_142_i, 
        un1_data_out8_76_set_net_1, un1_data_out8_198_rs_net_1, 
        \mem_9_rs[4] , \mem_9_[4]_net_1 , un1_data_out8_198_i, 
        un1_data_out8_101_set_net_1, un1_data_out8_174_rs_net_1, 
        \mem_10_rs[4] , \mem_10_[4]_net_1 , un1_data_out8_174_i, 
        un1_data_out8_92_set_net_1, un1_data_out8_230_rs_net_1, 
        \mem_11_rs[4] , \mem_11_[4]_net_1 , un1_data_out8_230_i, 
        un1_data_out8_20_set_net_1, un1_data_out8_244_rs_net_1, 
        \mem_12_rs[4] , \mem_12_[4]_net_1 , un1_data_out8_244_i, 
        un1_data_out8_108_set_net_1, un1_data_out8_212_rs_net_1, 
        \mem_13_rs[4] , \mem_13_[4]_net_1 , un1_data_out8_212_i, 
        un1_data_out8_116_set_net_1, un1_data_out8_220_rs_net_1, 
        \mem_14_rs[4] , \mem_14_[4]_net_1 , un1_data_out8_220_i, 
        un1_data_out8_15_set_net_1, un1_data_out8_155_rs_net_1, 
        \mem_1_rs[3] , \mem_1_[3]_net_1 , un1_data_out8_155_i, 
        un1_data_out8_31_set_net_1, un1_data_out8_163_rs_net_1, 
        \mem_2_rs[3] , \mem_2_[3]_net_1 , un1_data_out8_163_i, 
        un1_data_out8_127_set_net_1, un1_data_out8_131_rs_net_1, 
        \mem_3_rs[3] , \mem_3_[3]_net_1 , un1_data_out8_131_i, 
        un1_data_out8_6_set_net_1, un1_data_out8_139_rs_net_1, 
        \mem_4_rs[3] , \mem_4_[3]_net_1 , un1_data_out8_139_i, 
        un1_data_out8_41_set_net_1, un1_data_out8_193_rs_net_1, 
        \mem_5_rs[3] , \mem_5_[3]_net_1 , un1_data_out8_193_i, 
        un1_data_out8_34_set_net_1, un1_data_out8_169_rs_net_1, 
        \mem_6_rs[3] , \mem_6_[3]_net_1 , un1_data_out8_169_i, 
        un1_data_out8_50_set_net_1, un1_data_out8_225_rs_net_1, 
        \mem_7_rs[3] , \mem_7_[3]_net_1 , un1_data_out8_225_i, 
        un1_data_out8_66_set_net_1, un1_data_out8_241_rs_net_1, 
        \mem_8_rs[3] , \mem_8_[3]_net_1 , un1_data_out8_241_i, 
        un1_data_out8_75_set_net_1, un1_data_out8_196_rs_net_1, 
        \mem_9_rs[3] , \mem_9_[3]_net_1 , un1_data_out8_196_i, 
        un1_data_out8_96_set_net_1, un1_data_out8_172_rs_net_1, 
        \mem_10_rs[3] , \mem_10_[3]_net_1 , un1_data_out8_172_i, 
        un1_data_out8_91_set_net_1, un1_data_out8_228_rs_net_1, 
        \mem_11_rs[3] , \mem_11_[3]_net_1 , un1_data_out8_228_i, 
        un1_data_out8_19_set_net_1, un1_data_out8_243_rs_net_1, 
        \mem_12_rs[3] , \mem_12_[3]_net_1 , un1_data_out8_243_i, 
        un1_data_out8_107_set_net_1, un1_data_out8_211_rs_net_1, 
        \mem_13_rs[3] , \mem_13_[3]_net_1 , un1_data_out8_211_i, 
        un1_data_out8_115_set_net_1, un1_data_out8_219_rs_net_1, 
        \mem_14_rs[3] , \mem_14_[3]_net_1 , un1_data_out8_219_i, 
        un1_data_out8_56_set_net_1, un1_data_out8_250_rs_net_1, 
        \mem_15_rs[3] , \mem_15_[3]_net_1 , un1_data_out8_250_i, 
        un1_data_out8_29_set_net_1, un1_data_out8_162_rs_net_1, 
        \mem_2_rs[2] , \mem_2_[2]_net_1 , un1_data_out8_162_i, 
        un1_data_out8_125_set_net_1, un1_data_out8_130_rs_net_1, 
        \mem_3_rs[2] , \mem_3_[2]_net_1 , un1_data_out8_130_i, 
        un1_data_out8_4_set_net_1, un1_data_out8_138_rs_net_1, 
        \mem_4_rs[2] , \mem_4_[2]_net_1 , un1_data_out8_138_i, 
        un1_data_out8_43_set_net_1, un1_data_out8_191_rs_net_1, 
        \mem_5_rs[2] , \mem_5_[2]_net_1 , un1_data_out8_191_i, 
        un1_data_out8_32_set_net_1, un1_data_out8_207_rs_net_1, 
        \mem_6_rs[2] , \mem_6_[2]_net_1 , un1_data_out8_207_i, 
        un1_data_out8_48_set_net_1, un1_data_out8_183_rs_net_1, 
        \mem_7_rs[2] , \mem_7_[2]_net_1 , un1_data_out8_183_i, 
        un1_data_out8_64_set_net_1, un1_data_out8_239_rs_net_1, 
        \mem_8_rs[2] , \mem_8_[2]_net_1 , un1_data_out8_239_i, 
        un1_data_out8_74_set_net_1, un1_data_out8_194_rs_net_1, 
        \mem_9_rs[2] , \mem_9_[2]_net_1 , un1_data_out8_194_i, 
        un1_data_out8_99_set_net_1, un1_data_out8_170_rs_net_1, 
        \mem_10_rs[2] , \mem_10_[2]_net_1 , un1_data_out8_170_i, 
        un1_data_out8_90_set_net_1, un1_data_out8_226_rs_net_1, 
        \mem_11_rs[2] , \mem_11_[2]_net_1 , un1_data_out8_226_i, 
        un1_data_out8_18_set_net_1, un1_data_out8_242_rs_net_1, 
        \mem_12_rs[2] , \mem_12_[2]_net_1 , un1_data_out8_242_i, 
        un1_data_out8_106_set_net_1, un1_data_out8_210_rs_net_1, 
        \mem_13_rs[2] , \mem_13_[2]_net_1 , un1_data_out8_210_i, 
        un1_data_out8_114_set_net_1, un1_data_out8_218_rs_net_1, 
        \mem_14_rs[2] , \mem_14_[2]_net_1 , un1_data_out8_218_i, 
        un1_data_out8_59_set_net_1, un1_data_out8_249_rs_net_1, 
        \mem_15_rs[2] , \mem_15_[2]_net_1 , un1_data_out8_249_i, 
        un1_data_out8_83_set_net_1, un1_data_out8_146_rs_net_1, 
        \mem_0_rs[3] , \mem_0_[3]_net_1 , un1_data_out8_146_i, 
        un1_data_out8_123_set_net_1, un1_data_out8_129_rs_net_1, 
        \mem_3_rs[1] , \mem_3_[1]_net_1 , un1_data_out8_129_i, 
        un1_data_out8_2_set_net_1, un1_data_out8_137_rs_net_1, 
        \mem_4_rs[1] , \mem_4_[1]_net_1 , un1_data_out8_137_i, 
        un1_data_out8_14_set_net_1, un1_data_out8_189_rs_net_1, 
        \mem_5_rs[1] , \mem_5_[1]_net_1 , un1_data_out8_189_i, 
        un1_data_out8_30_set_net_1, un1_data_out8_205_rs_net_1, 
        \mem_6_rs[1] , \mem_6_[1]_net_1 , un1_data_out8_205_i, 
        un1_data_out8_126_set_net_1, un1_data_out8_181_rs_net_1, 
        \mem_7_rs[1] , \mem_7_[1]_net_1 , un1_data_out8_181_i, 
        un1_data_out8_5_set_net_1, un1_data_out8_237_rs_net_1, 
        \mem_8_rs[1] , \mem_8_[1]_net_1 , un1_data_out8_237_i, 
        un1_data_out8_73_set_net_1, un1_data_out8_192_rs_net_1, 
        \mem_9_rs[1] , \mem_9_[1]_net_1 , un1_data_out8_192_i, 
        un1_data_out8_98_set_net_1, un1_data_out8_168_rs_net_1, 
        \mem_10_rs[1] , \mem_10_[1]_net_1 , un1_data_out8_168_i, 
        un1_data_out8_89_set_net_1, un1_data_out8_224_rs_net_1, 
        \mem_11_rs[1] , \mem_11_[1]_net_1 , un1_data_out8_224_i, 
        un1_data_out8_17_set_net_1, un1_data_out8_240_rs_net_1, 
        \mem_12_rs[1] , \mem_12_[1]_net_1 , un1_data_out8_240_i, 
        un1_data_out8_105_set_net_1, un1_data_out8_209_rs_net_1, 
        \mem_13_rs[1] , \mem_13_[1]_net_1 , un1_data_out8_209_i, 
        un1_data_out8_113_set_net_1, un1_data_out8_217_rs_net_1, 
        \mem_14_rs[1] , \mem_14_[1]_net_1 , un1_data_out8_217_i, 
        un1_data_out8_58_set_net_1, un1_data_out8_248_rs_net_1, 
        \mem_15_rs[1] , \mem_15_[1]_net_1 , un1_data_out8_248_i, 
        un1_data_out8_82_set_net_1, un1_data_out8_145_rs_net_1, 
        \mem_0_rs[2] , \mem_0_[2]_net_1 , un1_data_out8_145_i, 
        un1_data_out8_13_set_net_1, un1_data_out8_154_rs_net_1, 
        \mem_1_rs[2] , \mem_1_[2]_net_1 , un1_data_out8_154_i, 
        un1_data_out8_set_net_1, un1_data_out8_136_rs_net_1, 
        \mem_4_rs[0] , \mem_4_[0]_net_1 , un1_data_out8_136_i, 
        un1_data_out8_12_set_net_1, un1_data_out8_187_rs_net_1, 
        \mem_5_rs[0] , \mem_5_[0]_net_1 , un1_data_out8_187_i, 
        un1_data_out8_28_set_net_1, un1_data_out8_203_rs_net_1, 
        \mem_6_rs[0] , \mem_6_[0]_net_1 , un1_data_out8_203_i, 
        un1_data_out8_124_set_net_1, un1_data_out8_179_rs_net_1, 
        \mem_7_rs[0] , \mem_7_[0]_net_1 , un1_data_out8_179_i, 
        un1_data_out8_7_set_net_1, un1_data_out8_235_rs_net_1, 
        \mem_8_rs[0] , \mem_8_[0]_net_1 , un1_data_out8_235_i, 
        un1_data_out8_72_set_net_1, un1_data_out8_190_rs_net_1, 
        \mem_9_rs[0] , \mem_9_[0]_net_1 , un1_data_out8_190_i, 
        un1_data_out8_97_set_net_1, un1_data_out8_206_rs_net_1, 
        \mem_10_rs[0] , \mem_10_[0]_net_1 , un1_data_out8_206_i, 
        un1_data_out8_88_set_net_1, un1_data_out8_182_rs_net_1, 
        \mem_11_rs[0] , \mem_11_[0]_net_1 , un1_data_out8_182_i, 
        un1_data_out8_16_set_net_1, un1_data_out8_238_rs_net_1, 
        \mem_12_rs[0] , \mem_12_[0]_net_1 , un1_data_out8_238_i, 
        un1_data_out8_104_set_net_1, un1_data_out8_208_rs_net_1, 
        \mem_13_rs[0] , \mem_13_[0]_net_1 , un1_data_out8_208_i, 
        un1_data_out8_112_set_net_1, un1_data_out8_216_rs_net_1, 
        \mem_14_rs[0] , \mem_14_[0]_net_1 , un1_data_out8_216_i, 
        un1_data_out8_57_set_net_1, un1_data_out8_251_rs_net_1, 
        \mem_15_rs[0] , \mem_15_[0]_net_1 , un1_data_out8_251_i, 
        un1_data_out8_81_set_net_1, un1_data_out8_144_rs_net_1, 
        \mem_0_rs[1] , \mem_0_[1]_net_1 , un1_data_out8_144_i, 
        un1_data_out8_11_set_net_1, un1_data_out8_153_rs_net_1, 
        \mem_1_rs[1] , \mem_1_[1]_net_1 , un1_data_out8_153_i, 
        un1_data_out8_27_set_net_1, un1_data_out8_161_rs_net_1, 
        \mem_2_rs[1] , \mem_2_[1]_net_1 , un1_data_out8_161_i, 
        un1_data_out8_80_set_net_1, un1_data_out8_147_rs_net_1, 
        \mem_0_rs[0] , \mem_0_[0]_net_1 , un1_data_out8_147_i, 
        un1_data_out8_9_set_net_1, un1_data_out8_152_rs_net_1, 
        \mem_1_rs[0] , \mem_1_[0]_net_1 , un1_data_out8_152_i, 
        un1_data_out8_25_set_net_1, un1_data_out8_160_rs_net_1, 
        \mem_2_rs[0] , \mem_2_[0]_net_1 , un1_data_out8_160_i, 
        un1_data_out8_121_set_net_1, un1_data_out8_128_rs_net_1, 
        \mem_3_rs[0] , \mem_3_[0]_net_1 , un1_data_out8_128_i, 
        \mem_5__2_i_0_0_a2[0] , \mem_14__2_i_0_0_a2[2] , 
        \mem_11__2_i_0_0_a2[2] , \mem_3__2_i_0_0_a2[0] , 
        \mem_6__2_i_0_0_a2[2] , \mem_13__2_i_0_0_a2[0] , 
        \mem_12__2_i_0_0_a2[0] , \mem_10__2_i_0_0_a2[0] , 
        \mem_1__2_i_0_0_a2[0] , \mem_7__2_i_0_0_a2[1] , 
        \mem_2__2_i_0_0_a2[0] , \mem_9__2_i_0_0_a2[0] , 
        \mem_4__2_i_0_0_a2[0] , \mem_15__2_i_0_0_a2[0] , 
        \data_out_2_15_i_i_a3_8[6]_net_1 , 
        \data_out_2_15_i_i_a3_8[5]_net_1 , 
        \data_out_2_15_i_i_a3_8[4]_net_1 , 
        \data_out_2_15_i_i_a3_8[2]_net_1 , N_641, N_413, N_397, N_381, 
        \data_out_2_15_i_i_7[2]_net_1 , \data_out_2_15_i_i_5[2]_net_1 , 
        \data_out_2_15_i_i_4[2]_net_1 , \data_out_2_15_i_i_3[2]_net_1 , 
        \data_out_2_15_i_i_2[2]_net_1 , \data_out_2_15_i_i_1[2]_net_1 , 
        \data_out_2_15_i_i_0[2]_net_1 , 
        \data_out_2_15_i_0_i_7[0]_net_1 , 
        \data_out_2_15_i_0_i_5[0]_net_1 , 
        \data_out_2_15_i_0_i_4[0]_net_1 , 
        \data_out_2_15_i_0_i_3[0]_net_1 , 
        \data_out_2_15_i_0_i_2[0]_net_1 , 
        \data_out_2_15_i_0_i_1[0]_net_1 , 
        \data_out_2_15_i_0_i_0[0]_net_1 , 
        \data_out_2_15_i_i_7[4]_net_1 , \data_out_2_15_i_i_5[4]_net_1 , 
        \data_out_2_15_i_i_4[4]_net_1 , \data_out_2_15_i_i_3[4]_net_1 , 
        \data_out_2_15_i_i_2[4]_net_1 , \data_out_2_15_i_i_1[4]_net_1 , 
        \data_out_2_15_i_i_0[4]_net_1 , 
        \data_out_2_15_i_0_i_7[7]_net_1 , 
        \data_out_2_15_i_0_i_5[7]_net_1 , 
        \data_out_2_15_i_0_i_4[7]_net_1 , 
        \data_out_2_15_i_0_i_3[7]_net_1 , 
        \data_out_2_15_i_0_i_2[7]_net_1 , 
        \data_out_2_15_i_0_i_1[7]_net_1 , 
        \data_out_2_15_i_0_i_0[7]_net_1 , 
        \data_out_2_15_i_i_7[5]_net_1 , \data_out_2_15_i_i_5[5]_net_1 , 
        \data_out_2_15_i_i_4[5]_net_1 , \data_out_2_15_i_i_3[5]_net_1 , 
        \data_out_2_15_i_i_2[5]_net_1 , \data_out_2_15_i_i_1[5]_net_1 , 
        \data_out_2_15_i_i_0[5]_net_1 , 
        \data_out_2_15_i_0_i_7[3]_net_1 , 
        \data_out_2_15_i_0_i_5[3]_net_1 , 
        \data_out_2_15_i_0_i_4[3]_net_1 , 
        \data_out_2_15_i_0_i_3[3]_net_1 , 
        \data_out_2_15_i_0_i_2[3]_net_1 , 
        \data_out_2_15_i_0_i_1[3]_net_1 , 
        \data_out_2_15_i_0_i_0[3]_net_1 , 
        \data_out_2_15_i_i_7[6]_net_1 , \data_out_2_15_i_i_5[6]_net_1 , 
        \data_out_2_15_i_i_4[6]_net_1 , \data_out_2_15_i_i_3[6]_net_1 , 
        \data_out_2_15_i_i_2[6]_net_1 , \data_out_2_15_i_i_1[6]_net_1 , 
        \data_out_2_15_i_i_0[6]_net_1 , 
        \data_out_2_15_i_0_i_7[1]_net_1 , 
        \data_out_2_15_i_0_i_5[1]_net_1 , 
        \data_out_2_15_i_0_i_4[1]_net_1 , 
        \data_out_2_15_i_0_i_3[1]_net_1 , 
        \data_out_2_15_i_0_i_2[1]_net_1 , 
        \data_out_2_15_i_0_i_1[1]_net_1 , 
        \data_out_2_15_i_0_i_0[1]_net_1 , 
        mem_14__1_sqmuxa_0_a2_0_a3_0_a2_net_1, 
        \data_out_2_15_i_i_11[2]_net_1 , 
        \data_out_2_15_i_0_i_11[0]_net_1 , 
        \data_out_2_15_i_i_11[4]_net_1 , 
        \data_out_2_15_i_0_i_11[7]_net_1 , 
        \data_out_2_15_i_i_11[5]_net_1 , 
        \data_out_2_15_i_0_i_11[3]_net_1 , 
        \data_out_2_15_i_i_11[6]_net_1 , 
        \data_out_2_15_i_0_i_11[1]_net_1 , 
        \data_out_2_15_i_i_12[2]_net_1 , 
        \data_out_2_15_i_0_i_12[0]_net_1 , 
        \data_out_2_15_i_i_12[4]_net_1 , 
        \data_out_2_15_i_0_i_12[7]_net_1 , 
        \data_out_2_15_i_i_12[5]_net_1 , 
        \data_out_2_15_i_0_i_12[3]_net_1 , 
        \data_out_2_15_i_i_12[6]_net_1 , 
        \data_out_2_15_i_0_i_12[1]_net_1 ;
    
    SLE un1_data_out8_2_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_4__1_sqmuxa), .ALn(un1_data_out8_2_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_data_out8_2_set_net_1));
    CFG3 #( .INIT(8'hF8) )  un1_data_out8_195_rs_RNIIQQ11 (.A(
        un1_data_out8_47_set_net_1), .B(un1_data_out8_195_rs_net_1), 
        .C(\mem_5_rs[4] ), .Y(\mem_5_[4]_net_1 ));
    SLE \mem_13_[4]  (.D(CoreAPB3_0_APBmslave4_PWDATA[4]), .CLK(
        FCCC_0_GL1), .EN(mem_13__1_sqmuxa), .ALn(un1_data_out8_212_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_13_rs[4] ));
    CFG3 #( .INIT(8'hF8) )  \mem_10__RNI19QJ[1]  (.A(
        un1_data_out8_98_set_net_1), .B(un1_data_out8_168_rs_net_1), 
        .C(\mem_10_rs[1] ), .Y(\mem_10_[1]_net_1 ));
    CFG1 #( .INIT(2'h1) )  un1_data_out8_88_set_RNO (.A(
        un1_data_out8_88_net_1), .Y(un1_data_out8_88_i));
    CFG1 #( .INIT(2'h1) )  un1_data_out8_117_set_RNO (.A(
        un1_data_out8_117_net_1), .Y(un1_data_out8_117_i));
    CFG3 #( .INIT(8'h02) )  un1_data_out8_88 (.A(\mem_11_[0]_net_1 ), 
        .B(\mem_11__2_i_0_0_a2[2] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_88_net_1));
    SLE \mem_4_[5]  (.D(CoreAPB3_0_APBmslave4_PWDATA[5]), .CLK(
        FCCC_0_GL1), .EN(mem_4__1_sqmuxa), .ALn(un1_data_out8_141_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_4_rs[5] ));
    SLE \mem_12_[2]  (.D(CoreAPB3_0_APBmslave4_PWDATA[2]), .CLK(
        FCCC_0_GL1), .EN(mem_12__1_sqmuxa), .ALn(un1_data_out8_242_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_12_rs[2] ));
    CFG3 #( .INIT(8'h02) )  un1_data_out8_59 (.A(\mem_15_[2]_net_1 ), 
        .B(\mem_15__2_i_0_0_a2[0] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_59_net_1));
    SLE un1_data_out8_11_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_1__1_sqmuxa), .ALn(un1_data_out8_11_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_data_out8_11_set_net_1));
    CFG4 #( .INIT(16'hEAC0) )  \data_out_2_15_i_0_i_0[3]  (.A(
        \mem_10_[3]_net_1 ), .B(\mem_12_[3]_net_1 ), .C(
        \mem_12__2_i_0_0_a2[0] ), .D(\mem_10__2_i_0_0_a2[0] ), .Y(
        \data_out_2_15_i_0_i_0[3]_net_1 ));
    SLE un1_data_out8_7_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_8__1_sqmuxa), .ALn(un1_data_out8_7_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_data_out8_7_set_net_1));
    CFG3 #( .INIT(8'hF2) )  un1_data_out8_184 (.A(\mem_8_[5]_net_1 ), 
        .B(mem_8__2_i_0_0_a2[2]), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_184_i));
    SLE un1_data_out8_70_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_8__1_sqmuxa), .ALn(un1_data_out8_70_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_data_out8_70_set_net_1));
    SLE un1_data_out8_219_rs (.D(VCC_net_1), .CLK(
        un1_data_out8_115_net_1), .EN(VCC_net_1), .ALn(
        un1_data_out8_219_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(VCC_net_1), .Q(un1_data_out8_219_rs_net_1));
    SLE un1_data_out8_241_rs (.D(VCC_net_1), .CLK(
        un1_data_out8_66_net_1), .EN(VCC_net_1), .ALn(
        un1_data_out8_241_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(VCC_net_1), .Q(un1_data_out8_241_rs_net_1));
    CFG3 #( .INIT(8'hF2) )  un1_data_out8_235 (.A(\mem_8_[0]_net_1 ), 
        .B(mem_8__2_i_0_0_a2[2]), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_235_i));
    SLE un1_data_out8_134_rs (.D(VCC_net_1), .CLK(
        un1_data_out8_53_net_1), .EN(VCC_net_1), .ALn(
        un1_data_out8_134_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(VCC_net_1), .Q(un1_data_out8_134_rs_net_1));
    SLE un1_data_out8_131_rs (.D(VCC_net_1), .CLK(
        un1_data_out8_127_net_1), .EN(VCC_net_1), .ALn(
        un1_data_out8_131_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(VCC_net_1), .Q(un1_data_out8_131_rs_net_1));
    SLE \mem_11_[4]  (.D(CoreAPB3_0_APBmslave4_PWDATA[4]), .CLK(
        FCCC_0_GL1), .EN(mem_11__1_sqmuxa), .ALn(un1_data_out8_230_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_11_rs[4] ));
    CFG3 #( .INIT(8'h02) )  un1_data_out8_32 (.A(\mem_6_[2]_net_1 ), 
        .B(\mem_6__2_i_0_0_a2[2] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_32_net_1));
    SLE \mem_13_[6]  (.D(CoreAPB3_0_APBmslave4_PWDATA[6]), .CLK(
        FCCC_0_GL1), .EN(mem_13__1_sqmuxa), .ALn(un1_data_out8_214_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_13_rs[6] ));
    SLE \mem_1_[2]  (.D(CoreAPB3_0_APBmslave4_PWDATA[2]), .CLK(
        FCCC_0_GL1), .EN(mem_1__1_sqmuxa), .ALn(un1_data_out8_154_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_1_rs[2] ));
    CFG3 #( .INIT(8'h02) )  un1_data_out8_83 (.A(\mem_0_[3]_net_1 ), 
        .B(mem_0__2_i_0_0_a2[0]), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_83_net_1));
    CFG3 #( .INIT(8'h02) )  un1_data_out8_78 (.A(\mem_9_[6]_net_1 ), 
        .B(\mem_9__2_i_0_0_a2[0] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_78_net_1));
    SLE \mem_9_[2]  (.D(CoreAPB3_0_APBmslave4_PWDATA[2]), .CLK(
        FCCC_0_GL1), .EN(mem_9__1_sqmuxa), .ALn(un1_data_out8_194_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_9_rs[2] ));
    SLE \mem_6_[1]  (.D(CoreAPB3_0_APBmslave4_PWDATA[1]), .CLK(
        FCCC_0_GL1), .EN(mem_6__1_sqmuxa), .ALn(un1_data_out8_205_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_6_rs[1] ));
    CFG3 #( .INIT(8'hF8) )  un1_data_out8_6_set_RNIPDKE (.A(
        un1_data_out8_6_set_net_1), .B(un1_data_out8_139_rs_net_1), .C(
        \mem_4_rs[3] ), .Y(\mem_4_[3]_net_1 ));
    CFG3 #( .INIT(8'hF2) )  un1_data_out8_134 (.A(\mem_3_[6]_net_1 ), 
        .B(\mem_3__2_i_0_0_a2[0] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_134_i));
    CFG3 #( .INIT(8'hF8) )  \mem_14__RNI42QK[4]  (.A(
        un1_data_out8_116_set_net_1), .B(un1_data_out8_220_rs_net_1), 
        .C(\mem_14_rs[4] ), .Y(\mem_14_[4]_net_1 ));
    CFG3 #( .INIT(8'hF8) )  un1_data_out8_222_rs_RNIAICF (.A(
        un1_data_out8_118_set_net_1), .B(un1_data_out8_222_rs_net_1), 
        .C(\mem_14_rs[6] ), .Y(\mem_14_[6]_net_1 ));
    CFG4 #( .INIT(16'hFFFE) )  \data_out_2_15_i_i_12[6]  (.A(
        \data_out_2_15_i_i_2[6]_net_1 ), .B(
        \data_out_2_15_i_i_1[6]_net_1 ), .C(
        \data_out_2_15_i_i_3[6]_net_1 ), .D(
        \data_out_2_15_i_i_0[6]_net_1 ), .Y(
        \data_out_2_15_i_i_12[6]_net_1 ));
    CFG3 #( .INIT(8'h02) )  un1_data_out8_125 (.A(\mem_3_[2]_net_1 ), 
        .B(\mem_3__2_i_0_0_a2[0] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_125_net_1));
    SLE un1_data_out8_36_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_6__1_sqmuxa), .ALn(un1_data_out8_36_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_data_out8_36_set_net_1));
    CFG4 #( .INIT(16'hECA0) )  \data_out_2_15_i_0_i_4[0]  (.A(
        \mem_6_[0]_net_1 ), .B(\mem_4_[0]_net_1 ), .C(
        \mem_6__2_i_0_0_a2[2] ), .D(\mem_4__2_i_0_0_a2[0] ), .Y(
        \data_out_2_15_i_0_i_4[0]_net_1 ));
    CFG2 #( .INIT(4'h8) )  \data_out_2_15_i_0_i_a3_8[3]  (.A(
        \mem_3__2_i_0_0_a2[0] ), .B(\mem_3_[3]_net_1 ), .Y(N_397));
    SLE un1_data_out8_252_rs (.D(VCC_net_1), .CLK(
        un1_data_out8_62_net_1), .EN(VCC_net_1), .ALn(
        un1_data_out8_252_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(VCC_net_1), .Q(un1_data_out8_252_rs_net_1));
    CFG3 #( .INIT(8'hF2) )  un1_data_out8_206 (.A(\mem_10_[0]_net_1 ), 
        .B(\mem_10__2_i_0_0_a2[0] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_206_i));
    CFG3 #( .INIT(8'h02) )  un1_data_out8_35 (.A(\mem_2_[5]_net_1 ), 
        .B(\mem_2__2_i_0_0_a2[0] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_35_net_1));
    SLE un1_data_out8_9_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_1__1_sqmuxa), .ALn(un1_data_out8_9_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_data_out8_9_set_net_1));
    SLE \mem_11_[6]  (.D(CoreAPB3_0_APBmslave4_PWDATA[6]), .CLK(
        FCCC_0_GL1), .EN(mem_11__1_sqmuxa), .ALn(un1_data_out8_234_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_11_rs[6] ));
    SLE un1_data_out8_43_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_5__1_sqmuxa), .ALn(un1_data_out8_43_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_data_out8_43_set_net_1));
    CFG1 #( .INIT(2'h1) )  un1_data_out8_118_set_RNO (.A(
        un1_data_out8_118_net_1), .Y(un1_data_out8_118_i));
    SLE \mem_0_[1]  (.D(CoreAPB3_0_APBmslave4_PWDATA[1]), .CLK(
        FCCC_0_GL1), .EN(mem_0__1_sqmuxa), .ALn(un1_data_out8_144_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_0_rs[1] ));
    CFG3 #( .INIT(8'h02) )  un1_data_out8_73 (.A(\mem_9_[1]_net_1 ), 
        .B(\mem_9__2_i_0_0_a2[0] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_73_net_1));
    CFG3 #( .INIT(8'hF8) )  \mem_2__RNIE2FF[6]  (.A(
        un1_data_out8_37_set_net_1), .B(un1_data_out8_166_rs_net_1), 
        .C(\mem_2_rs[6] ), .Y(\mem_2_[6]_net_1 ));
    CFG3 #( .INIT(8'h02) )  un1_data_out8_117 (.A(\mem_14_[5]_net_1 ), 
        .B(\mem_14__2_i_0_0_a2[2] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_117_net_1));
    CFG3 #( .INIT(8'hF2) )  un1_data_out8_155 (.A(\mem_1_[3]_net_1 ), 
        .B(\mem_1__2_i_0_0_a2[0] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_155_i));
    CFG2 #( .INIT(4'h8) )  mem_6__1_sqmuxa_0_a2_0_a3_0_a3 (.A(
        mem_14__1_sqmuxa_0_a2_0_a3_0_a2_net_1), .B(
        \mem_6__2_i_0_0_a2[2] ), .Y(mem_6__1_sqmuxa));
    CFG1 #( .INIT(2'h1) )  un1_data_out8_12_set_RNO (.A(
        un1_data_out8_12_net_1), .Y(un1_data_out8_12_i));
    CFG3 #( .INIT(8'h02) )  un1_data_out8_34 (.A(\mem_6_[3]_net_1 ), 
        .B(\mem_6__2_i_0_0_a2[2] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_34_net_1));
    CFG2 #( .INIT(4'h8) )  \data_out_2_15_i_0_i_a3_8[7]  (.A(
        \mem_3__2_i_0_0_a2[0] ), .B(\mem_3_[7]_net_1 ), .Y(N_381));
    SLE un1_data_out8_230_rs (.D(VCC_net_1), .CLK(
        un1_data_out8_92_net_1), .EN(VCC_net_1), .ALn(
        un1_data_out8_230_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(VCC_net_1), .Q(un1_data_out8_230_rs_net_1));
    SLE un1_data_out8_160_rs (.D(VCC_net_1), .CLK(
        un1_data_out8_25_net_1), .EN(VCC_net_1), .ALn(
        un1_data_out8_160_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(VCC_net_1), .Q(un1_data_out8_160_rs_net_1));
    CFG3 #( .INIT(8'h02) )  un1_data_out8_87 (.A(\mem_0_[7]_net_1 ), 
        .B(mem_0__2_i_0_0_a2[0]), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_87_net_1));
    SLE un1_data_out8_44_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_1__1_sqmuxa), .ALn(un1_data_out8_44_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_data_out8_44_set_net_1));
    SLE un1_data_out8_205_rs (.D(VCC_net_1), .CLK(
        un1_data_out8_30_net_1), .EN(VCC_net_1), .ALn(
        un1_data_out8_205_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(VCC_net_1), .Q(un1_data_out8_205_rs_net_1));
    CFG1 #( .INIT(2'h1) )  un1_data_out8_104_set_RNO (.A(
        un1_data_out8_104_net_1), .Y(un1_data_out8_104_i));
    CFG3 #( .INIT(8'hF2) )  un1_data_out8_174 (.A(\mem_10_[4]_net_1 ), 
        .B(\mem_10__2_i_0_0_a2[0] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_174_i));
    CFG3 #( .INIT(8'hF2) )  un1_data_out8_228 (.A(\mem_11_[3]_net_1 ), 
        .B(\mem_11__2_i_0_0_a2[2] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_228_i));
    CFG3 #( .INIT(8'hF2) )  un1_data_out8_145 (.A(\mem_0_[2]_net_1 ), 
        .B(mem_0__2_i_0_0_a2[0]), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_145_i));
    CFG3 #( .INIT(8'hF8) )  un1_data_out8_137_rs_RNIHLLB (.A(
        un1_data_out8_2_set_net_1), .B(un1_data_out8_137_rs_net_1), .C(
        \mem_4_rs[1] ), .Y(\mem_4_[1]_net_1 ));
    CFG1 #( .INIT(2'h1) )  un1_data_out8_82_set_RNO (.A(
        un1_data_out8_82_net_1), .Y(un1_data_out8_82_i));
    SLE un1_data_out8_220_rs (.D(VCC_net_1), .CLK(
        un1_data_out8_116_net_1), .EN(VCC_net_1), .ALn(
        un1_data_out8_220_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(VCC_net_1), .Q(un1_data_out8_220_rs_net_1));
    SLE un1_data_out8_242_rs (.D(VCC_net_1), .CLK(
        un1_data_out8_18_net_1), .EN(VCC_net_1), .ALn(
        un1_data_out8_242_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(VCC_net_1), .Q(un1_data_out8_242_rs_net_1));
    CFG3 #( .INIT(8'hF8) )  un1_data_out8_216_rs_RNI1SD6 (.A(
        un1_data_out8_112_set_net_1), .B(un1_data_out8_216_rs_net_1), 
        .C(\mem_14_rs[0] ), .Y(\mem_14_[0]_net_1 ));
    SLE \mem_8_[3]  (.D(CoreAPB3_0_APBmslave4_PWDATA[3]), .CLK(
        FCCC_0_GL1), .EN(mem_8__1_sqmuxa), .ALn(un1_data_out8_241_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_8_rs[3] ));
    SLE un1_data_out8_13_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_1__1_sqmuxa), .ALn(un1_data_out8_13_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_data_out8_13_set_net_1));
    CFG3 #( .INIT(8'hF2) )  un1_data_out8_231 (.A(\mem_7_[6]_net_1 ), 
        .B(\mem_7__2_i_0_0_a2[1] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_231_i));
    CFG4 #( .INIT(16'hFFFE) )  \data_out_2_15_i_i_12[2]  (.A(
        \data_out_2_15_i_i_2[2]_net_1 ), .B(
        \data_out_2_15_i_i_1[2]_net_1 ), .C(
        \data_out_2_15_i_i_3[2]_net_1 ), .D(
        \data_out_2_15_i_i_0[2]_net_1 ), .Y(
        \data_out_2_15_i_i_12[2]_net_1 ));
    CFG4 #( .INIT(16'hEAC0) )  \data_out_2_15_i_0_i_2[0]  (.A(
        \mem_13_[0]_net_1 ), .B(\mem_11_[0]_net_1 ), .C(
        \mem_11__2_i_0_0_a2[2] ), .D(\mem_13__2_i_0_0_a2[0] ), .Y(
        \data_out_2_15_i_0_i_2[0]_net_1 ));
    CFG1 #( .INIT(2'h1) )  un1_data_out8_64_set_RNO (.A(
        un1_data_out8_64_net_1), .Y(un1_data_out8_64_i));
    CFG3 #( .INIT(8'h02) )  un1_data_out8_77 (.A(\mem_9_[5]_net_1 ), 
        .B(\mem_9__2_i_0_0_a2[0] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_77_net_1));
    CFG4 #( .INIT(16'hFFFE) )  \data_out_2_15_i_i[4]  (.A(
        \data_out_2_15_i_i_4[4]_net_1 ), .B(
        \data_out_2_15_i_i_5[4]_net_1 ), .C(
        \data_out_2_15_i_i_12[4]_net_1 ), .D(
        \data_out_2_15_i_i_11[4]_net_1 ), .Y(N_15));
    SLE un1_data_out8_97_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_10__1_sqmuxa), .ALn(un1_data_out8_97_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_data_out8_97_set_net_1));
    CFG3 #( .INIT(8'hF8) )  un1_data_out8_14_set_RNIC4GM (.A(
        un1_data_out8_14_set_net_1), .B(un1_data_out8_189_rs_net_1), 
        .C(\mem_5_rs[1] ), .Y(\mem_5_[1]_net_1 ));
    CFG2 #( .INIT(4'h8) )  mem_8__1_sqmuxa_0_a2_0_a3_0_a3 (.A(
        mem_14__1_sqmuxa_0_a2_0_a3_0_a2_net_1), .B(
        mem_8__2_i_0_0_a2[2]), .Y(mem_8__1_sqmuxa));
    SLE \mem_1_[1]  (.D(CoreAPB3_0_APBmslave4_PWDATA[1]), .CLK(
        FCCC_0_GL1), .EN(mem_1__1_sqmuxa), .ALn(un1_data_out8_153_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_1_rs[1] ));
    SLE \mem_9_[1]  (.D(CoreAPB3_0_APBmslave4_PWDATA[1]), .CLK(
        FCCC_0_GL1), .EN(mem_9__1_sqmuxa), .ALn(un1_data_out8_192_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_9_rs[1] ));
    CFG4 #( .INIT(16'hEAC0) )  \data_out_2_15_i_i_0[5]  (.A(
        \mem_10_[5]_net_1 ), .B(\mem_12_[5]_net_1 ), .C(
        \mem_12__2_i_0_0_a2[0] ), .D(\mem_10__2_i_0_0_a2[0] ), .Y(
        \data_out_2_15_i_i_0[5]_net_1 ));
    SLE \mem_12_[7]  (.D(CoreAPB3_0_APBmslave4_PWDATA[7]), .CLK(
        FCCC_0_GL1), .EN(mem_12__1_sqmuxa), .ALn(un1_data_out8_247_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_12_rs[7] ));
    CFG3 #( .INIT(8'hF8) )  un1_data_out8_152_rs_RNIHTAV (.A(
        un1_data_out8_9_set_net_1), .B(un1_data_out8_152_rs_net_1), .C(
        \mem_1_rs[0] ), .Y(\mem_1_[0]_net_1 ));
    CFG3 #( .INIT(8'hF2) )  un1_data_out8_129 (.A(\mem_3_[1]_net_1 ), 
        .B(\mem_3__2_i_0_0_a2[0] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_129_i));
    CFG4 #( .INIT(16'hFFF8) )  \data_out_2_15_i_i_11[4]  (.A(
        \mem_5__2_i_0_0_a2[0] ), .B(\mem_5_[4]_net_1 ), .C(
        \data_out_2_15_i_i_7[4]_net_1 ), .D(
        \data_out_2_15_i_i_a3_8[4]_net_1 ), .Y(
        \data_out_2_15_i_i_11[4]_net_1 ));
    SLE un1_data_out8_14_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_5__1_sqmuxa), .ALn(un1_data_out8_14_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_data_out8_14_set_net_1));
    SLE \mem_14_[0]  (.D(CoreAPB3_0_APBmslave4_PWDATA[0]), .CLK(
        FCCC_0_GL1), .EN(mem_14__1_sqmuxa), .ALn(un1_data_out8_216_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_14_rs[0] ));
    CFG3 #( .INIT(8'hF8) )  un1_data_out8_119_set_RNIDQL4 (.A(
        un1_data_out8_119_set_net_1), .B(un1_data_out8_223_rs_net_1), 
        .C(\mem_14_rs[7] ), .Y(\mem_14_[7]_net_1 ));
    CFG3 #( .INIT(8'hF8) )  un1_data_out8_60_set_RNIT81Q (.A(
        un1_data_out8_60_set_net_1), .B(un1_data_out8_254_rs_net_1), 
        .C(\mem_15_rs[7] ), .Y(\mem_15_[7]_net_1 ));
    CFG3 #( .INIT(8'hF2) )  un1_data_out8_248 (.A(\mem_15_[1]_net_1 ), 
        .B(\mem_15__2_i_0_0_a2[0] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_248_i));
    CFG3 #( .INIT(8'hF8) )  un1_data_out8_100_set_RNI1BDF (.A(
        un1_data_out8_100_set_net_1), .B(un1_data_out8_180_rs_net_1), 
        .C(\mem_10_rs[7] ), .Y(\mem_10_[7]_net_1 ));
    SLE \mem_10_[5]  (.D(CoreAPB3_0_APBmslave4_PWDATA[5]), .CLK(
        FCCC_0_GL1), .EN(mem_10__1_sqmuxa), .ALn(un1_data_out8_176_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_10_rs[5] ));
    CFG3 #( .INIT(8'hF8) )  un1_data_out8_110_set_RNI2GL71 (.A(
        un1_data_out8_110_set_net_1), .B(un1_data_out8_214_rs_net_1), 
        .C(\mem_13_rs[6] ), .Y(\mem_13_[6]_net_1 ));
    CFG3 #( .INIT(8'hF2) )  un1_data_out8_180 (.A(\mem_10_[7]_net_1 ), 
        .B(\mem_10__2_i_0_0_a2[0] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_180_i));
    SLE un1_data_out8_4_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_4__1_sqmuxa), .ALn(un1_data_out8_4_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_data_out8_4_set_net_1));
    SLE \data_out[5]  (.D(N_17), .CLK(FCCC_0_GL1), .EN(rd_enable), 
        .ALn(MSS_RESET_N_M2F_c), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(
        CoreAPB3_0_APBmslave5_PRDATA[5]));
    CFG4 #( .INIT(16'h0020) )  \WRITE_GEN.mem_5__2_i_0_0_a2[0]  (.A(
        CoreAPB3_0_APBmslave4_PADDR[2]), .B(
        CoreAPB3_0_APBmslave4_PADDR[5]), .C(
        CoreAPB3_0_APBmslave4_PADDR[4]), .D(
        CoreAPB3_0_APBmslave4_PADDR[3]), .Y(\mem_5__2_i_0_0_a2[0] ));
    SLE \mem_5_[2]  (.D(CoreAPB3_0_APBmslave4_PWDATA[2]), .CLK(
        FCCC_0_GL1), .EN(mem_5__1_sqmuxa), .ALn(un1_data_out8_191_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_5_rs[2] ));
    CFG3 #( .INIT(8'hF8) )  un1_data_out8_10_set_RNI9A5D (.A(
        un1_data_out8_10_set_net_1), .B(un1_data_out8_185_rs_net_1), 
        .C(\mem_4_rs[7] ), .Y(\mem_4_[7]_net_1 ));
    CFG1 #( .INIT(2'h1) )  un1_data_out8_34_set_RNO (.A(
        un1_data_out8_34_net_1), .Y(un1_data_out8_34_i));
    CFG3 #( .INIT(8'hF2) )  un1_data_out8_159 (.A(\mem_1_[7]_net_1 ), 
        .B(\mem_1__2_i_0_0_a2[0] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_159_i));
    CFG3 #( .INIT(8'hF8) )  un1_data_out8_231_rs_RNILT5G (.A(
        un1_data_out8_3_set_net_1), .B(un1_data_out8_231_rs_net_1), .C(
        \mem_7_rs[6] ), .Y(\mem_7_[6]_net_1 ));
    CFG3 #( .INIT(8'hF8) )  un1_data_out8_22_set_RNIOHIQ (.A(
        un1_data_out8_22_set_net_1), .B(un1_data_out8_246_rs_net_1), 
        .C(\mem_12_rs[6] ), .Y(\mem_12_[6]_net_1 ));
    CFG1 #( .INIT(2'h1) )  un1_data_out8_67_set_RNO (.A(
        un1_data_out8_67_net_1), .Y(un1_data_out8_67_i));
    CFG1 #( .INIT(2'h1) )  un1_data_out8_54_set_RNO (.A(
        un1_data_out8_54_net_1), .Y(un1_data_out8_54_i));
    CFG3 #( .INIT(8'hF8) )  un1_data_out8_202_rs_RNIHN171 (.A(
        un1_data_out8_78_set_net_1), .B(un1_data_out8_202_rs_net_1), 
        .C(\mem_9_rs[6] ), .Y(\mem_9_[6]_net_1 ));
    SLE \mem_6_[6]  (.D(CoreAPB3_0_APBmslave4_PWDATA[6]), .CLK(
        FCCC_0_GL1), .EN(mem_6__1_sqmuxa), .ALn(un1_data_out8_175_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_6_rs[6] ));
    SLE un1_data_out8_48_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_7__1_sqmuxa), .ALn(un1_data_out8_48_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_data_out8_48_set_net_1));
    SLE \mem_10_[1]  (.D(CoreAPB3_0_APBmslave4_PWDATA[1]), .CLK(
        FCCC_0_GL1), .EN(mem_10__1_sqmuxa), .ALn(un1_data_out8_168_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_10_rs[1] ));
    CFG3 #( .INIT(8'hF8) )  \mem_15__RNIPFOP[0]  (.A(
        un1_data_out8_57_set_net_1), .B(un1_data_out8_251_rs_net_1), 
        .C(\mem_15_rs[0] ), .Y(\mem_15_[0]_net_1 ));
    CFG3 #( .INIT(8'hF2) )  un1_data_out8_237 (.A(\mem_8_[1]_net_1 ), 
        .B(mem_8__2_i_0_0_a2[2]), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_237_i));
    CFG3 #( .INIT(8'hF2) )  un1_data_out8_162 (.A(\mem_2_[2]_net_1 ), 
        .B(\mem_2__2_i_0_0_a2[0] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_162_i));
    CFG1 #( .INIT(2'h1) )  un1_data_out8_44_set_RNO (.A(
        un1_data_out8_44_net_1), .Y(un1_data_out8_44_i));
    CFG3 #( .INIT(8'hF2) )  un1_data_out8_130 (.A(\mem_3_[2]_net_1 ), 
        .B(\mem_3__2_i_0_0_a2[0] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_130_i));
    CFG3 #( .INIT(8'hF2) )  un1_data_out8_149 (.A(\mem_0_[5]_net_1 ), 
        .B(mem_0__2_i_0_0_a2[0]), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_149_i));
    CFG4 #( .INIT(16'hECA0) )  \data_out_2_15_i_0_i_1[7]  (.A(
        \mem_14_[7]_net_1 ), .B(\mem_9_[7]_net_1 ), .C(
        \mem_14__2_i_0_0_a2[2] ), .D(\mem_9__2_i_0_0_a2[0] ), .Y(
        \data_out_2_15_i_0_i_1[7]_net_1 ));
    SLE un1_data_out8_194_rs (.D(VCC_net_1), .CLK(
        un1_data_out8_74_net_1), .EN(VCC_net_1), .ALn(
        un1_data_out8_194_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(VCC_net_1), .Q(un1_data_out8_194_rs_net_1));
    CFG4 #( .INIT(16'hEAC0) )  \data_out_2_15_i_0_i_2[7]  (.A(
        \mem_13_[7]_net_1 ), .B(\mem_11_[7]_net_1 ), .C(
        \mem_11__2_i_0_0_a2[2] ), .D(\mem_13__2_i_0_0_a2[0] ), .Y(
        \data_out_2_15_i_0_i_2[7]_net_1 ));
    SLE un1_data_out8_191_rs (.D(VCC_net_1), .CLK(
        un1_data_out8_43_net_1), .EN(VCC_net_1), .ALn(
        un1_data_out8_191_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(VCC_net_1), .Q(un1_data_out8_191_rs_net_1));
    SLE \mem_0_[6]  (.D(CoreAPB3_0_APBmslave4_PWDATA[6]), .CLK(
        FCCC_0_GL1), .EN(mem_0__1_sqmuxa), .ALn(un1_data_out8_150_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_0_rs[6] ));
    SLE un1_data_out8_8_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_4__1_sqmuxa), .ALn(un1_data_out8_8_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_data_out8_8_set_net_1));
    CFG3 #( .INIT(8'hF2) )  un1_data_out8_128 (.A(\mem_3_[0]_net_1 ), 
        .B(\mem_3__2_i_0_0_a2[0] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_128_i));
    CFG3 #( .INIT(8'hF2) )  un1_data_out8_214 (.A(\mem_13_[6]_net_1 ), 
        .B(\mem_13__2_i_0_0_a2[0] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_214_i));
    CFG1 #( .INIT(2'h1) )  un1_data_out8_20_set_RNO (.A(
        un1_data_out8_20_net_1), .Y(un1_data_out8_20_i));
    CFG3 #( .INIT(8'h02) )  un1_data_out8_12 (.A(\mem_5_[0]_net_1 ), 
        .B(\mem_5__2_i_0_0_a2[0] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_12_net_1));
    CFG3 #( .INIT(8'hF8) )  \mem_14__RNI44NB[1]  (.A(
        un1_data_out8_113_set_net_1), .B(un1_data_out8_217_rs_net_1), 
        .C(\mem_14_rs[1] ), .Y(\mem_14_[1]_net_1 ));
    CFG4 #( .INIT(16'hEAC0) )  \data_out_2_15_i_i_0[4]  (.A(
        \mem_10_[4]_net_1 ), .B(\mem_12_[4]_net_1 ), .C(
        \mem_12__2_i_0_0_a2[0] ), .D(\mem_10__2_i_0_0_a2[0] ), .Y(
        \data_out_2_15_i_i_0[4]_net_1 ));
    SLE un1_data_out8_154_rs (.D(VCC_net_1), .CLK(
        un1_data_out8_13_net_1), .EN(VCC_net_1), .ALn(
        un1_data_out8_154_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(VCC_net_1), .Q(un1_data_out8_154_rs_net_1));
    SLE un1_data_out8_151_rs (.D(VCC_net_1), .CLK(
        un1_data_out8_87_net_1), .EN(VCC_net_1), .ALn(
        un1_data_out8_151_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(VCC_net_1), .Q(un1_data_out8_151_rs_net_1));
    SLE un1_data_out8_95_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_11__1_sqmuxa), .ALn(un1_data_out8_95_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_data_out8_95_set_net_1));
    CFG1 #( .INIT(2'h1) )  un1_data_out8_37_set_RNO (.A(
        un1_data_out8_37_net_1), .Y(un1_data_out8_37_i));
    CFG3 #( .INIT(8'hF2) )  un1_data_out8_183 (.A(\mem_7_[2]_net_1 ), 
        .B(\mem_7__2_i_0_0_a2[1] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_183_i));
    CFG4 #( .INIT(16'hECA0) )  \data_out_2_15_i_i_1[6]  (.A(
        \mem_14_[6]_net_1 ), .B(\mem_9_[6]_net_1 ), .C(
        \mem_14__2_i_0_0_a2[2] ), .D(\mem_9__2_i_0_0_a2[0] ), .Y(
        \data_out_2_15_i_i_1[6]_net_1 ));
    SLE un1_data_out8_236_rs (.D(VCC_net_1), .CLK(
        un1_data_out8_95_net_1), .EN(VCC_net_1), .ALn(
        un1_data_out8_236_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(VCC_net_1), .Q(un1_data_out8_236_rs_net_1));
    SLE un1_data_out8_170_rs (.D(VCC_net_1), .CLK(
        un1_data_out8_99_net_1), .EN(VCC_net_1), .ALn(
        un1_data_out8_170_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(VCC_net_1), .Q(un1_data_out8_170_rs_net_1));
    SLE un1_data_out8_39_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_2__1_sqmuxa), .ALn(un1_data_out8_39_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_data_out8_39_set_net_1));
    CFG1 #( .INIT(2'h1) )  un1_data_out8_28_set_RNO (.A(
        un1_data_out8_28_net_1), .Y(un1_data_out8_28_i));
    CFG3 #( .INIT(8'hF2) )  un1_data_out8_233 (.A(\mem_7_[7]_net_1 ), 
        .B(\mem_7__2_i_0_0_a2[1] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_233_i));
    CFG1 #( .INIT(2'h1) )  un1_data_out8_57_set_RNO (.A(
        un1_data_out8_57_net_1), .Y(un1_data_out8_57_i));
    CFG3 #( .INIT(8'hF8) )  un1_data_out8_230_rs_RNILOQJ (.A(
        un1_data_out8_92_set_net_1), .B(un1_data_out8_230_rs_net_1), 
        .C(\mem_11_rs[4] ), .Y(\mem_11_[4]_net_1 ));
    CFG3 #( .INIT(8'hF8) )  un1_data_out8_123_set_RNILUEL (.A(
        un1_data_out8_123_set_net_1), .B(un1_data_out8_129_rs_net_1), 
        .C(\mem_3_rs[1] ), .Y(\mem_3_[1]_net_1 ));
    SLE un1_data_out8_211_rs (.D(VCC_net_1), .CLK(
        un1_data_out8_107_net_1), .EN(VCC_net_1), .ALn(
        un1_data_out8_211_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(VCC_net_1), .Q(un1_data_out8_211_rs_net_1));
    CFG4 #( .INIT(16'hEAC0) )  \data_out_2_15_i_i_3[2]  (.A(
        \mem_15_[2]_net_1 ), .B(\mem_7_[2]_net_1 ), .C(
        \mem_7__2_i_0_0_a2[1] ), .D(\mem_15__2_i_0_0_a2[0] ), .Y(
        \data_out_2_15_i_i_3[2]_net_1 ));
    SLE un1_data_out8_208_rs (.D(VCC_net_1), .CLK(
        un1_data_out8_104_net_1), .EN(VCC_net_1), .ALn(
        un1_data_out8_208_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(VCC_net_1), .Q(un1_data_out8_208_rs_net_1));
    SLE un1_data_out8_18_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_12__1_sqmuxa), .ALn(un1_data_out8_18_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_data_out8_18_set_net_1));
    CFG3 #( .INIT(8'hF2) )  un1_data_out8_158 (.A(\mem_1_[6]_net_1 ), 
        .B(\mem_1__2_i_0_0_a2[0] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_158_i));
    CFG4 #( .INIT(16'hEAC0) )  \data_out_2_15_i_0_i_2[1]  (.A(
        \mem_13_[1]_net_1 ), .B(\mem_11_[1]_net_1 ), .C(
        \mem_11__2_i_0_0_a2[2] ), .D(\mem_13__2_i_0_0_a2[0] ), .Y(
        \data_out_2_15_i_0_i_2[1]_net_1 ));
    CFG3 #( .INIT(8'h02) )  un1_data_out8_15 (.A(\mem_1_[3]_net_1 ), 
        .B(\mem_1__2_i_0_0_a2[0] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_15_net_1));
    CFG1 #( .INIT(2'h1) )  un1_data_out8_47_set_RNO (.A(
        un1_data_out8_47_net_1), .Y(un1_data_out8_47_i));
    CFG3 #( .INIT(8'hF8) )  \mem_3__RNIHIVR[0]  (.A(
        un1_data_out8_121_set_net_1), .B(un1_data_out8_128_rs_net_1), 
        .C(\mem_3_rs[0] ), .Y(\mem_3_[0]_net_1 ));
    SLE un1_data_out8_226_rs (.D(VCC_net_1), .CLK(
        un1_data_out8_90_net_1), .EN(VCC_net_1), .ALn(
        un1_data_out8_226_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(VCC_net_1), .Q(un1_data_out8_226_rs_net_1));
    CFG1 #( .INIT(2'h1) )  un1_data_out8_66_set_RNO (.A(
        un1_data_out8_66_net_1), .Y(un1_data_out8_66_i));
    CFG3 #( .INIT(8'hF2) )  un1_data_out8_170 (.A(\mem_10_[2]_net_1 ), 
        .B(\mem_10__2_i_0_0_a2[0] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_170_i));
    CFG3 #( .INIT(8'h02) )  un1_data_out8_102 (.A(\mem_10_[5]_net_1 ), 
        .B(\mem_10__2_i_0_0_a2[0] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_102_net_1));
    CFG3 #( .INIT(8'hF2) )  un1_data_out8_133 (.A(\mem_3_[5]_net_1 ), 
        .B(\mem_3__2_i_0_0_a2[0] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_133_i));
    SLE un1_data_out8_31_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_2__1_sqmuxa), .ALn(un1_data_out8_31_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_data_out8_31_set_net_1));
    CFG3 #( .INIT(8'hF8) )  un1_data_out8_82_set_RNI5G7C (.A(
        un1_data_out8_82_set_net_1), .B(un1_data_out8_145_rs_net_1), 
        .C(\mem_0_rs[2] ), .Y(\mem_0_[2]_net_1 ));
    CFG3 #( .INIT(8'hF2) )  un1_data_out8_148 (.A(\mem_0_[4]_net_1 ), 
        .B(mem_0__2_i_0_0_a2[0]), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_148_i));
    CFG3 #( .INIT(8'h02) )  un1_data_out8_14 (.A(\mem_5_[1]_net_1 ), 
        .B(\mem_5__2_i_0_0_a2[0] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_14_net_1));
    SLE \mem_5_[1]  (.D(CoreAPB3_0_APBmslave4_PWDATA[1]), .CLK(
        FCCC_0_GL1), .EN(mem_5__1_sqmuxa), .ALn(un1_data_out8_189_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_5_rs[1] ));
    CFG3 #( .INIT(8'h02) )  un1_data_out8_89 (.A(\mem_11_[1]_net_1 ), 
        .B(\mem_11__2_i_0_0_a2[2] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_89_net_1));
    SLE un1_data_out8_144_rs (.D(VCC_net_1), .CLK(
        un1_data_out8_81_net_1), .EN(VCC_net_1), .ALn(
        un1_data_out8_144_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(VCC_net_1), .Q(un1_data_out8_144_rs_net_1));
    SLE un1_data_out8_141_rs (.D(VCC_net_1), .CLK(
        un1_data_out8_67_net_1), .EN(VCC_net_1), .ALn(
        un1_data_out8_141_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(VCC_net_1), .Q(un1_data_out8_141_rs_net_1));
    CFG3 #( .INIT(8'hF8) )  un1_data_out8_16_set_RNIMO0V (.A(
        un1_data_out8_16_set_net_1), .B(un1_data_out8_238_rs_net_1), 
        .C(\mem_12_rs[0] ), .Y(\mem_12_[0]_net_1 ));
    CFG3 #( .INIT(8'hF2) )  un1_data_out8_167 (.A(\mem_2_[7]_net_1 ), 
        .B(\mem_2__2_i_0_0_a2[0] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_167_i));
    GND GND (.Y(GND_net_1));
    SLE un1_data_out8_250_rs (.D(VCC_net_1), .CLK(
        un1_data_out8_56_net_1), .EN(VCC_net_1), .ALn(
        un1_data_out8_250_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(VCC_net_1), .Q(un1_data_out8_250_rs_net_1));
    CFG3 #( .INIT(8'hF2) )  un1_data_out8_194 (.A(\mem_9_[2]_net_1 ), 
        .B(\mem_9__2_i_0_0_a2[0] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_194_i));
    SLE \mem_15_[2]  (.D(CoreAPB3_0_APBmslave4_PWDATA[2]), .CLK(
        FCCC_0_GL1), .EN(mem_15__1_sqmuxa), .ALn(un1_data_out8_249_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_15_rs[2] ));
    SLE un1_data_out8_184_rs (.D(VCC_net_1), .CLK(
        un1_data_out8_69_net_1), .EN(VCC_net_1), .ALn(
        un1_data_out8_184_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(VCC_net_1), .Q(un1_data_out8_184_rs_net_1));
    SLE \mem_1_[6]  (.D(CoreAPB3_0_APBmslave4_PWDATA[6]), .CLK(
        FCCC_0_GL1), .EN(mem_1__1_sqmuxa), .ALn(un1_data_out8_158_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_1_rs[6] ));
    CFG4 #( .INIT(16'hEAC0) )  \data_out_2_15_i_i_4[6]  (.A(
        \mem_4_[6]_net_1 ), .B(\mem_2_[6]_net_1 ), .C(
        \mem_2__2_i_0_0_a2[0] ), .D(\mem_4__2_i_0_0_a2[0] ), .Y(
        \data_out_2_15_i_i_4[6]_net_1 ));
    SLE un1_data_out8_181_rs (.D(VCC_net_1), .CLK(
        un1_data_out8_126_net_1), .EN(VCC_net_1), .ALn(
        un1_data_out8_181_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(VCC_net_1), .Q(un1_data_out8_181_rs_net_1));
    CFG4 #( .INIT(16'hEAC0) )  \data_out_2_15_i_0_i_4[3]  (.A(
        \mem_4_[3]_net_1 ), .B(\mem_2_[3]_net_1 ), .C(
        \mem_2__2_i_0_0_a2[0] ), .D(\mem_4__2_i_0_0_a2[0] ), .Y(
        \data_out_2_15_i_0_i_4[3]_net_1 ));
    SLE \mem_9_[6]  (.D(CoreAPB3_0_APBmslave4_PWDATA[6]), .CLK(
        FCCC_0_GL1), .EN(mem_9__1_sqmuxa), .ALn(un1_data_out8_202_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_9_rs[6] ));
    CFG4 #( .INIT(16'hFFF8) )  \data_out_2_15_i_0_i_11[3]  (.A(
        \mem_5__2_i_0_0_a2[0] ), .B(\mem_5_[3]_net_1 ), .C(
        \data_out_2_15_i_0_i_7[3]_net_1 ), .D(N_397), .Y(
        \data_out_2_15_i_0_i_11[3]_net_1 ));
    SLE un1_data_out8_92_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_11__1_sqmuxa), .ALn(un1_data_out8_92_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_data_out8_92_set_net_1));
    SLE \mem_8_[4]  (.D(CoreAPB3_0_APBmslave4_PWDATA[4]), .CLK(
        FCCC_0_GL1), .EN(mem_8__1_sqmuxa), .ALn(un1_data_out8_142_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_8_rs[4] ));
    CFG4 #( .INIT(16'hEAC0) )  \data_out_2_15_i_0_i_2[3]  (.A(
        \mem_13_[3]_net_1 ), .B(\mem_11_[3]_net_1 ), .C(
        \mem_11__2_i_0_0_a2[2] ), .D(\mem_13__2_i_0_0_a2[0] ), .Y(
        \data_out_2_15_i_0_i_2[3]_net_1 ));
    CFG3 #( .INIT(8'hF8) )  un1_data_out8_106_set_RNIVI321 (.A(
        un1_data_out8_106_set_net_1), .B(un1_data_out8_210_rs_net_1), 
        .C(\mem_13_rs[2] ), .Y(\mem_13_[2]_net_1 ));
    SLE \mem_13_[3]  (.D(CoreAPB3_0_APBmslave4_PWDATA[3]), .CLK(
        FCCC_0_GL1), .EN(mem_13__1_sqmuxa), .ALn(un1_data_out8_211_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_13_rs[3] ));
    CFG1 #( .INIT(2'h1) )  un1_data_out8_90_set_RNO (.A(
        un1_data_out8_90_net_1), .Y(un1_data_out8_90_i));
    CFG1 #( .INIT(2'h1) )  un1_data_out8_36_set_RNO (.A(
        un1_data_out8_36_net_1), .Y(un1_data_out8_36_i));
    CFG3 #( .INIT(8'h02) )  un1_data_out8_28 (.A(\mem_6_[0]_net_1 ), 
        .B(\mem_6__2_i_0_0_a2[2] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_28_net_1));
    CFG3 #( .INIT(8'hF8) )  \mem_2__RNI6AGC[4]  (.A(
        un1_data_out8_33_set_net_1), .B(un1_data_out8_164_rs_net_1), 
        .C(\mem_2_rs[4] ), .Y(\mem_2_[4]_net_1 ));
    CFG1 #( .INIT(2'h1) )  un1_data_out8_56_set_RNO (.A(
        un1_data_out8_56_net_1), .Y(un1_data_out8_56_i));
    CFG1 #( .INIT(2'h1) )  un1_data_out8_98_set_RNO (.A(
        un1_data_out8_98_net_1), .Y(un1_data_out8_98_i));
    CFG3 #( .INIT(8'hF8) )  un1_data_out8_97_set_RNIOAJE (.A(
        un1_data_out8_97_set_net_1), .B(un1_data_out8_206_rs_net_1), 
        .C(\mem_10_rs[0] ), .Y(\mem_10_[0]_net_1 ));
    CFG3 #( .INIT(8'h02) )  un1_data_out8_79 (.A(\mem_9_[7]_net_1 ), 
        .B(\mem_9__2_i_0_0_a2[0] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_79_net_1));
    SLE un1_data_out8_137_rs (.D(VCC_net_1), .CLK(
        un1_data_out8_2_net_1), .EN(VCC_net_1), .ALn(
        un1_data_out8_137_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(VCC_net_1), .Q(un1_data_out8_137_rs_net_1));
    CFG4 #( .INIT(16'hEAC0) )  \data_out_2_15_i_i_3[5]  (.A(
        \mem_15_[5]_net_1 ), .B(\mem_7_[5]_net_1 ), .C(
        \mem_7__2_i_0_0_a2[1] ), .D(\mem_15__2_i_0_0_a2[0] ), .Y(
        \data_out_2_15_i_i_3[5]_net_1 ));
    CFG3 #( .INIT(8'h02) )  un1_data_out8_92 (.A(\mem_11_[4]_net_1 ), 
        .B(\mem_11__2_i_0_0_a2[2] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_92_net_1));
    CFG3 #( .INIT(8'h02) )  un1_data_out8_48 (.A(\mem_7_[2]_net_1 ), 
        .B(\mem_7__2_i_0_0_a2[1] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_48_net_1));
    CFG3 #( .INIT(8'hF2) )  un1_data_out8_173 (.A(\mem_6_[5]_net_1 ), 
        .B(\mem_6__2_i_0_0_a2[2] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_173_i));
    CFG1 #( .INIT(2'h1) )  un1_data_out8_46_set_RNO (.A(
        un1_data_out8_46_net_1), .Y(un1_data_out8_46_i));
    CFG3 #( .INIT(8'h02) )  un1_data_out8_31 (.A(\mem_2_[3]_net_1 ), 
        .B(\mem_2__2_i_0_0_a2[0] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_31_net_1));
    SLE \mem_11_[3]  (.D(CoreAPB3_0_APBmslave4_PWDATA[3]), .CLK(
        FCCC_0_GL1), .EN(mem_11__1_sqmuxa), .ALn(un1_data_out8_228_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_11_rs[3] ));
    CFG4 #( .INIT(16'hFFF8) )  \data_out_2_15_i_i_11[5]  (.A(
        \mem_5__2_i_0_0_a2[0] ), .B(\mem_5_[5]_net_1 ), .C(
        \data_out_2_15_i_i_7[5]_net_1 ), .D(
        \data_out_2_15_i_i_a3_8[5]_net_1 ), .Y(
        \data_out_2_15_i_i_11[5]_net_1 ));
    CFG3 #( .INIT(8'hF2) )  un1_data_out8_239 (.A(\mem_8_[2]_net_1 ), 
        .B(mem_8__2_i_0_0_a2[2]), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_239_i));
    SLE un1_data_out8_212_rs (.D(VCC_net_1), .CLK(
        un1_data_out8_108_net_1), .EN(VCC_net_1), .ALn(
        un1_data_out8_212_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(VCC_net_1), .Q(un1_data_out8_212_rs_net_1));
    SLE \mem_7_[3]  (.D(CoreAPB3_0_APBmslave4_PWDATA[3]), .CLK(
        FCCC_0_GL1), .EN(mem_7__1_sqmuxa), .ALn(un1_data_out8_225_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_7_rs[3] ));
    SLE un1_data_out8_204_rs (.D(VCC_net_1), .CLK(
        un1_data_out8_79_net_1), .EN(VCC_net_1), .ALn(
        un1_data_out8_204_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(VCC_net_1), .Q(un1_data_out8_204_rs_net_1));
    CFG3 #( .INIT(8'hF8) )  un1_data_out8_187_rs_RNI7LTR (.A(
        un1_data_out8_12_set_net_1), .B(un1_data_out8_187_rs_net_1), 
        .C(\mem_5_rs[0] ), .Y(\mem_5_[0]_net_1 ));
    CFG4 #( .INIT(16'hEAC0) )  \data_out_2_15_i_0_i_4[1]  (.A(
        \mem_4_[1]_net_1 ), .B(\mem_2_[1]_net_1 ), .C(
        \mem_2__2_i_0_0_a2[0] ), .D(\mem_4__2_i_0_0_a2[0] ), .Y(
        \data_out_2_15_i_0_i_4[1]_net_1 ));
    SLE un1_data_out8_240_rs (.D(VCC_net_1), .CLK(
        un1_data_out8_17_net_1), .EN(VCC_net_1), .ALn(
        un1_data_out8_240_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(VCC_net_1), .Q(un1_data_out8_240_rs_net_1));
    CFG3 #( .INIT(8'h02) )  un1_data_out8_23 (.A(\mem_12_[7]_net_1 ), 
        .B(\mem_12__2_i_0_0_a2[0] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_23_net_1));
    CFG2 #( .INIT(4'h8) )  mem_4__1_sqmuxa_0_a3_0_a3 (.A(
        mem_14__1_sqmuxa_0_a2_0_a3_0_a2_net_1), .B(
        \mem_4__2_i_0_0_a2[0] ), .Y(mem_4__1_sqmuxa));
    CFG1 #( .INIT(2'h1) )  un1_data_out8_22_set_RNO (.A(
        un1_data_out8_22_net_1), .Y(un1_data_out8_22_i));
    CFG3 #( .INIT(8'hF8) )  un1_data_out8_184_rs_RNIOI4M (.A(
        un1_data_out8_69_set_net_1), .B(un1_data_out8_184_rs_net_1), 
        .C(\mem_8_rs[5] ), .Y(\mem_8_[5]_net_1 ));
    CFG3 #( .INIT(8'h02) )  un1_data_out8_115 (.A(\mem_14_[3]_net_1 ), 
        .B(\mem_14__2_i_0_0_a2[2] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_115_net_1));
    SLE \mem_2_[3]  (.D(CoreAPB3_0_APBmslave4_PWDATA[3]), .CLK(
        FCCC_0_GL1), .EN(mem_2__1_sqmuxa), .ALn(un1_data_out8_163_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_2_rs[3] ));
    CFG4 #( .INIT(16'hECA0) )  \data_out_2_15_i_0_i_1[3]  (.A(
        \mem_14_[3]_net_1 ), .B(\mem_9_[3]_net_1 ), .C(
        \mem_14__2_i_0_0_a2[2] ), .D(\mem_9__2_i_0_0_a2[0] ), .Y(
        \data_out_2_15_i_0_i_1[3]_net_1 ));
    CFG3 #( .INIT(8'h02) )  un1_data_out8_107 (.A(\mem_13_[3]_net_1 ), 
        .B(\mem_13__2_i_0_0_a2[0] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_107_net_1));
    CFG4 #( .INIT(16'h0800) )  \WRITE_GEN.mem_11__2_i_0_0_a2[2]  (.A(
        CoreAPB3_0_APBmslave4_PADDR[2]), .B(
        CoreAPB3_0_APBmslave4_PADDR[5]), .C(
        CoreAPB3_0_APBmslave4_PADDR[4]), .D(
        CoreAPB3_0_APBmslave4_PADDR[3]), .Y(\mem_11__2_i_0_0_a2[2] ));
    CFG3 #( .INIT(8'h02) )  un1_data_out8_95 (.A(\mem_11_[7]_net_1 ), 
        .B(\mem_11__2_i_0_0_a2[2] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_95_net_1));
    CFG3 #( .INIT(8'hF8) )  un1_data_out8_41_set_RNI9RFM (.A(
        un1_data_out8_41_set_net_1), .B(un1_data_out8_193_rs_net_1), 
        .C(\mem_5_rs[3] ), .Y(\mem_5_[3]_net_1 ));
    CFG3 #( .INIT(8'h02) )  un1_data_out8_43 (.A(\mem_5_[2]_net_1 ), 
        .B(\mem_5__2_i_0_0_a2[0] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_43_net_1));
    SLE \mem_8_[0]  (.D(CoreAPB3_0_APBmslave4_PWDATA[0]), .CLK(
        FCCC_0_GL1), .EN(mem_8__1_sqmuxa), .ALn(un1_data_out8_235_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_8_rs[0] ));
    SLE \mem_4_[3]  (.D(CoreAPB3_0_APBmslave4_PWDATA[3]), .CLK(
        FCCC_0_GL1), .EN(mem_4__1_sqmuxa), .ALn(un1_data_out8_139_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_4_rs[3] ));
    CFG3 #( .INIT(8'hF8) )  \mem_10__RNISPDJ[2]  (.A(
        un1_data_out8_99_set_net_1), .B(un1_data_out8_170_rs_net_1), 
        .C(\mem_10_rs[2] ), .Y(\mem_10_[2]_net_1 ));
    CFG3 #( .INIT(8'h02) )  un1_data_out8_94 (.A(\mem_11_[6]_net_1 ), 
        .B(\mem_11__2_i_0_0_a2[2] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_94_net_1));
    CFG3 #( .INIT(8'h02) )  un1_data_out8_121 (.A(\mem_3_[0]_net_1 ), 
        .B(\mem_3__2_i_0_0_a2[0] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_121_net_1));
    CFG4 #( .INIT(16'hECA0) )  \data_out_2_15_i_i_1[2]  (.A(
        \mem_14_[2]_net_1 ), .B(\mem_9_[2]_net_1 ), .C(
        \mem_14__2_i_0_0_a2[2] ), .D(\mem_9__2_i_0_0_a2[0] ), .Y(
        \data_out_2_15_i_i_1[2]_net_1 ));
    SLE un1_data_out8_33_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_2__1_sqmuxa), .ALn(un1_data_out8_33_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_data_out8_33_set_net_1));
    CFG1 #( .INIT(2'h1) )  un1_data_out8_123_set_RNO (.A(
        un1_data_out8_123_net_1), .Y(un1_data_out8_123_i));
    CFG4 #( .INIT(16'hECA0) )  \data_out_2_15_i_i_5[6]  (.A(
        \mem_6_[6]_net_1 ), .B(\mem_1_[6]_net_1 ), .C(
        \mem_6__2_i_0_0_a2[2] ), .D(\mem_1__2_i_0_0_a2[0] ), .Y(
        \data_out_2_15_i_i_5[6]_net_1 ));
    CFG3 #( .INIT(8'h02) )  un1_data_out8_27 (.A(\mem_2_[1]_net_1 ), 
        .B(\mem_2__2_i_0_0_a2[0] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_27_net_1));
    CFG3 #( .INIT(8'hF2) )  un1_data_out8_218 (.A(\mem_14_[2]_net_1 ), 
        .B(\mem_14__2_i_0_0_a2[2] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_218_i));
    CFG1 #( .INIT(2'h1) )  un1_data_out8_63_set_RNO (.A(
        un1_data_out8_63_net_1), .Y(un1_data_out8_63_i));
    CFG3 #( .INIT(8'hF8) )  \mem_3__RNI8EOO[6]  (.A(
        un1_data_out8_53_set_net_1), .B(un1_data_out8_134_rs_net_1), 
        .C(\mem_3_rs[6] ), .Y(\mem_3_[6]_net_1 ));
    SLE un1_data_out8_57_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_15__1_sqmuxa), .ALn(un1_data_out8_57_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_data_out8_57_set_net_1));
    CFG1 #( .INIT(2'h1) )  un1_data_out8_101_set_RNO (.A(
        un1_data_out8_101_net_1), .Y(un1_data_out8_101_i));
    CFG3 #( .INIT(8'hF8) )  un1_data_out8_29_set_RNI7L49 (.A(
        un1_data_out8_29_set_net_1), .B(un1_data_out8_162_rs_net_1), 
        .C(\mem_2_rs[2] ), .Y(\mem_2_[2]_net_1 ));
    CFG3 #( .INIT(8'hF2) )  un1_data_out8_151 (.A(\mem_0_[7]_net_1 ), 
        .B(mem_0__2_i_0_0_a2[0]), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_151_i));
    CFG1 #( .INIT(2'h1) )  un1_data_out8_125_set_RNO (.A(
        un1_data_out8_125_net_1), .Y(un1_data_out8_125_i));
    SLE un1_data_out8_34_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_6__1_sqmuxa), .ALn(un1_data_out8_34_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_data_out8_34_set_net_1));
    CFG3 #( .INIT(8'h02) )  un1_data_out8_126 (.A(\mem_7_[1]_net_1 ), 
        .B(\mem_7__2_i_0_0_a2[1] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_126_net_1));
    CFG3 #( .INIT(8'h02) )  un1_data_out8_47 (.A(\mem_5_[4]_net_1 ), 
        .B(\mem_5__2_i_0_0_a2[0] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_47_net_1));
    CFG4 #( .INIT(16'hEAC0) )  \data_out_2_15_i_0_i_3[0]  (.A(
        \mem_15_[0]_net_1 ), .B(\mem_7_[0]_net_1 ), .C(
        \mem_7__2_i_0_0_a2[1] ), .D(\mem_15__2_i_0_0_a2[0] ), .Y(
        \data_out_2_15_i_0_i_3[0]_net_1 ));
    CFG3 #( .INIT(8'hF8) )  \mem_8__RNIPMA31[1]  (.A(
        un1_data_out8_5_set_net_1), .B(un1_data_out8_237_rs_net_1), .C(
        \mem_8_rs[1] ), .Y(\mem_8_[1]_net_1 ));
    CFG1 #( .INIT(2'h1) )  un1_data_out8_92_set_RNO (.A(
        un1_data_out8_92_net_1), .Y(un1_data_out8_92_i));
    SLE \mem_5_[6]  (.D(CoreAPB3_0_APBmslave4_PWDATA[6]), .CLK(
        FCCC_0_GL1), .EN(mem_5__1_sqmuxa), .ALn(un1_data_out8_199_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_5_rs[6] ));
    CFG1 #( .INIT(2'h1) )  un1_data_out8_127_set_RNO (.A(
        un1_data_out8_127_net_1), .Y(un1_data_out8_127_i));
    CFG3 #( .INIT(8'hF8) )  un1_data_out8_64_set_RNIHR0S (.A(
        un1_data_out8_64_set_net_1), .B(un1_data_out8_239_rs_net_1), 
        .C(\mem_8_rs[2] ), .Y(\mem_8_[2]_net_1 ));
    CFG3 #( .INIT(8'hF8) )  un1_data_out8_156_rs_RNI41241 (.A(
        un1_data_out8_40_set_net_1), .B(un1_data_out8_156_rs_net_1), 
        .C(\mem_1_rs[4] ), .Y(\mem_1_[4]_net_1 ));
    SLE un1_data_out8_164_rs (.D(VCC_net_1), .CLK(
        un1_data_out8_33_net_1), .EN(VCC_net_1), .ALn(
        un1_data_out8_164_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(VCC_net_1), .Q(un1_data_out8_164_rs_net_1));
    SLE \mem_15_[7]  (.D(CoreAPB3_0_APBmslave4_PWDATA[7]), .CLK(
        FCCC_0_GL1), .EN(mem_15__1_sqmuxa), .ALn(un1_data_out8_254_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_15_rs[7] ));
    SLE un1_data_out8_161_rs (.D(VCC_net_1), .CLK(
        un1_data_out8_27_net_1), .EN(VCC_net_1), .ALn(
        un1_data_out8_161_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(VCC_net_1), .Q(un1_data_out8_161_rs_net_1));
    CFG3 #( .INIT(8'hF8) )  un1_data_out8_240_rs_RNIH9KU (.A(
        un1_data_out8_17_set_net_1), .B(un1_data_out8_240_rs_net_1), 
        .C(\mem_12_rs[1] ), .Y(\mem_12_[1]_net_1 ));
    CFG3 #( .INIT(8'hF2) )  un1_data_out8_141 (.A(\mem_4_[5]_net_1 ), 
        .B(\mem_4__2_i_0_0_a2[0] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_141_i));
    CFG3 #( .INIT(8'hF8) )  \mem_14__RNI7C0H[2]  (.A(
        un1_data_out8_114_set_net_1), .B(un1_data_out8_218_rs_net_1), 
        .C(\mem_14_rs[2] ), .Y(\mem_14_[2]_net_1 ));
    CFG3 #( .INIT(8'hF2) )  un1_data_out8_190 (.A(\mem_9_[0]_net_1 ), 
        .B(\mem_9__2_i_0_0_a2[0] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_190_i));
    CFG3 #( .INIT(8'hF8) )  un1_data_out8_94_set_RNITEJG (.A(
        un1_data_out8_94_set_net_1), .B(un1_data_out8_234_rs_net_1), 
        .C(\mem_11_rs[6] ), .Y(\mem_11_[6]_net_1 ));
    CFG1 #( .INIT(2'h1) )  un1_data_out8_106_set_RNO (.A(
        un1_data_out8_106_net_1), .Y(un1_data_out8_106_i));
    CFG3 #( .INIT(8'h02) )  un1_data_out8_119 (.A(\mem_14_[7]_net_1 ), 
        .B(\mem_14__2_i_0_0_a2[2] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_119_net_1));
    CFG1 #( .INIT(2'h1) )  un1_data_out8_33_set_RNO (.A(
        un1_data_out8_33_net_1), .Y(un1_data_out8_33_i));
    CFG3 #( .INIT(8'hF2) )  un1_data_out8_156 (.A(\mem_1_[4]_net_1 ), 
        .B(\mem_1__2_i_0_0_a2[0] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_156_i));
    CFG3 #( .INIT(8'hF8) )  un1_data_out8_18_set_RNILK0L (.A(
        un1_data_out8_18_set_net_1), .B(un1_data_out8_242_rs_net_1), 
        .C(\mem_12_rs[2] ), .Y(\mem_12_[2]_net_1 ));
    CFG2 #( .INIT(4'h8) )  mem_12__1_sqmuxa_0_a3_0_a3 (.A(
        mem_14__1_sqmuxa_0_a2_0_a3_0_a2_net_1), .B(
        \mem_12__2_i_0_0_a2[0] ), .Y(mem_12__1_sqmuxa));
    SLE un1_data_out8_96_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_10__1_sqmuxa), .ALn(un1_data_out8_96_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_data_out8_96_set_net_1));
    CFG3 #( .INIT(8'hF2) )  un1_data_out8_236 (.A(\mem_11_[7]_net_1 ), 
        .B(\mem_11__2_i_0_0_a2[2] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_236_i));
    CFG1 #( .INIT(2'h1) )  un1_data_out8_53_set_RNO (.A(
        un1_data_out8_53_net_1), .Y(un1_data_out8_53_i));
    SLE \mem_12_[5]  (.D(CoreAPB3_0_APBmslave4_PWDATA[5]), .CLK(
        FCCC_0_GL1), .EN(mem_12__1_sqmuxa), .ALn(un1_data_out8_245_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_12_rs[5] ));
    SLE \mem_13_[0]  (.D(CoreAPB3_0_APBmslave4_PWDATA[0]), .CLK(
        FCCC_0_GL1), .EN(mem_13__1_sqmuxa), .ALn(un1_data_out8_208_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_13_rs[0] ));
    SLE un1_data_out8_40_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_1__1_sqmuxa), .ALn(un1_data_out8_40_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_data_out8_40_set_net_1));
    CFG1 #( .INIT(2'h1) )  un1_data_out8_43_set_RNO (.A(
        un1_data_out8_43_net_1), .Y(un1_data_out8_43_i));
    CFG3 #( .INIT(8'hF2) )  un1_data_out8_146 (.A(\mem_0_[3]_net_1 ), 
        .B(mem_0__2_i_0_0_a2[0]), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_146_i));
    CFG4 #( .INIT(16'hFFFE) )  \data_out_2_15_i_i[6]  (.A(
        \data_out_2_15_i_i_4[6]_net_1 ), .B(
        \data_out_2_15_i_i_5[6]_net_1 ), .C(
        \data_out_2_15_i_i_12[6]_net_1 ), .D(
        \data_out_2_15_i_i_11[6]_net_1 ), .Y(N_19));
    SLE un1_data_out8_246_rs (.D(VCC_net_1), .CLK(
        un1_data_out8_22_net_1), .EN(VCC_net_1), .ALn(
        un1_data_out8_246_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(VCC_net_1), .Q(un1_data_out8_246_rs_net_1));
    SLE un1_data_out8_203_rs (.D(VCC_net_1), .CLK(
        un1_data_out8_28_net_1), .EN(VCC_net_1), .ALn(
        un1_data_out8_203_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(VCC_net_1), .Q(un1_data_out8_203_rs_net_1));
    CFG3 #( .INIT(8'h02) )  un1_data_out8_3 (.A(\mem_7_[6]_net_1 ), .B(
        \mem_7__2_i_0_0_a2[1] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_3_net_1));
    CFG3 #( .INIT(8'hF8) )  un1_data_out8_19_set_RNIOS9Q (.A(
        un1_data_out8_19_set_net_1), .B(un1_data_out8_243_rs_net_1), 
        .C(\mem_12_rs[3] ), .Y(\mem_12_[3]_net_1 ));
    CFG1 #( .INIT(2'h1) )  un1_data_out8_100_set_RNO (.A(
        un1_data_out8_100_net_1), .Y(un1_data_out8_100_i));
    CFG2 #( .INIT(4'h8) )  mem_14__1_sqmuxa_0_a2_0_a3_0_a3 (.A(
        mem_14__1_sqmuxa_0_a2_0_a3_0_a2_net_1), .B(
        \mem_14__2_i_0_0_a2[2] ), .Y(mem_14__1_sqmuxa));
    SLE \mem_12_[1]  (.D(CoreAPB3_0_APBmslave4_PWDATA[1]), .CLK(
        FCCC_0_GL1), .EN(mem_12__1_sqmuxa), .ALn(un1_data_out8_240_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_12_rs[1] ));
    CFG3 #( .INIT(8'hF2) )  un1_data_out8_204 (.A(\mem_9_[7]_net_1 ), 
        .B(\mem_9__2_i_0_0_a2[0] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_204_i));
    SLE un1_data_out8_136_rs (.D(VCC_net_1), .CLK(un1_data_out8_net_1), 
        .EN(VCC_net_1), .ALn(un1_data_out8_136_i), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(VCC_net_1), .Q(
        un1_data_out8_136_rs_net_1));
    SLE \mem_11_[0]  (.D(CoreAPB3_0_APBmslave4_PWDATA[0]), .CLK(
        FCCC_0_GL1), .EN(mem_11__1_sqmuxa), .ALn(un1_data_out8_182_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_11_rs[0] ));
    SLE un1_data_out8_55_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_3__1_sqmuxa), .ALn(un1_data_out8_55_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_data_out8_55_set_net_1));
    CFG3 #( .INIT(8'h02) )  un1_data_out8_62 (.A(\mem_15_[5]_net_1 ), 
        .B(\mem_15__2_i_0_0_a2[0] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_62_net_1));
    SLE un1_data_out8_197_rs (.D(VCC_net_1), .CLK(
        un1_data_out8_45_net_1), .EN(VCC_net_1), .ALn(
        un1_data_out8_197_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(VCC_net_1), .Q(un1_data_out8_197_rs_net_1));
    CFG4 #( .INIT(16'hECA0) )  \data_out_2_15_i_i_5[2]  (.A(
        \mem_6_[2]_net_1 ), .B(\mem_1_[2]_net_1 ), .C(
        \mem_6__2_i_0_0_a2[2] ), .D(\mem_1__2_i_0_0_a2[0] ), .Y(
        \data_out_2_15_i_i_5[2]_net_1 ));
    CFG3 #( .INIT(8'hF2) )  un1_data_out8_193 (.A(\mem_5_[3]_net_1 ), 
        .B(\mem_5__2_i_0_0_a2[0] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_193_i));
    SLE \mem_3_[7]  (.D(CoreAPB3_0_APBmslave4_PWDATA[7]), .CLK(
        FCCC_0_GL1), .EN(mem_3__1_sqmuxa), .ALn(un1_data_out8_135_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_3_rs[7] ));
    SLE un1_data_out8_38_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_6__1_sqmuxa), .ALn(un1_data_out8_38_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_data_out8_38_set_net_1));
    SLE \mem_7_[4]  (.D(CoreAPB3_0_APBmslave4_PWDATA[4]), .CLK(
        FCCC_0_GL1), .EN(mem_7__1_sqmuxa), .ALn(un1_data_out8_227_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_7_rs[4] ));
    SLE un1_data_out8_113_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_14__1_sqmuxa), .ALn(un1_data_out8_113_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_data_out8_113_set_net_1));
    SLE un1_data_out8_67_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_4__1_sqmuxa), .ALn(un1_data_out8_67_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_data_out8_67_set_net_1));
    SLE un1_data_out8_157_rs (.D(VCC_net_1), .CLK(
        un1_data_out8_42_net_1), .EN(VCC_net_1), .ALn(
        un1_data_out8_157_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(VCC_net_1), .Q(un1_data_out8_157_rs_net_1));
    CFG3 #( .INIT(8'hF8) )  \mem_11__RNIQ77K[3]  (.A(
        un1_data_out8_91_set_net_1), .B(un1_data_out8_228_rs_net_1), 
        .C(\mem_11_rs[3] ), .Y(\mem_11_[3]_net_1 ));
    CFG3 #( .INIT(8'h02) )  un1_data_out8_118 (.A(\mem_14_[6]_net_1 ), 
        .B(\mem_14__2_i_0_0_a2[2] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_118_net_1));
    CFG3 #( .INIT(8'hF8) )  un1_data_out8_108_set_RNI53MS (.A(
        un1_data_out8_108_set_net_1), .B(un1_data_out8_212_rs_net_1), 
        .C(\mem_13_rs[4] ), .Y(\mem_13_[4]_net_1 ));
    CFG3 #( .INIT(8'h02) )  un1_data_out8_11 (.A(\mem_1_[1]_net_1 ), 
        .B(\mem_1__2_i_0_0_a2[0] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_11_net_1));
    SLE un1_data_out8_123_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_3__1_sqmuxa), .ALn(un1_data_out8_123_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_data_out8_123_set_net_1));
    CFG2 #( .INIT(4'h8) )  mem_5__1_sqmuxa_0_a3_0_a3 (.A(
        mem_14__1_sqmuxa_0_a2_0_a3_0_a2_net_1), .B(
        \mem_5__2_i_0_0_a2[0] ), .Y(mem_5__1_sqmuxa));
    SLE \mem_2_[4]  (.D(CoreAPB3_0_APBmslave4_PWDATA[4]), .CLK(
        FCCC_0_GL1), .EN(mem_2__1_sqmuxa), .ALn(un1_data_out8_164_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_2_rs[4] ));
    SLE \mem_3_[5]  (.D(CoreAPB3_0_APBmslave4_PWDATA[5]), .CLK(
        FCCC_0_GL1), .EN(mem_3__1_sqmuxa), .ALn(un1_data_out8_133_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_3_rs[5] ));
    CFG3 #( .INIT(8'hF8) )  un1_data_out8_7_set_RNIONGP (.A(
        un1_data_out8_7_set_net_1), .B(un1_data_out8_235_rs_net_1), .C(
        \mem_8_rs[0] ), .Y(\mem_8_[0]_net_1 ));
    SLE un1_data_out8_10_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_4__1_sqmuxa), .ALn(un1_data_out8_10_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_data_out8_10_set_net_1));
    SLE un1_data_out8_103_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_10__1_sqmuxa), .ALn(un1_data_out8_103_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_data_out8_103_set_net_1));
    SLE un1_data_out8_139_rs (.D(VCC_net_1), .CLK(
        un1_data_out8_6_net_1), .EN(VCC_net_1), .ALn(
        un1_data_out8_139_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(VCC_net_1), .Q(un1_data_out8_139_rs_net_1));
    CFG3 #( .INIT(8'h02) )  un1_data_out8_65 (.A(\mem_4_[4]_net_1 ), 
        .B(\mem_4__2_i_0_0_a2[0] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_65_net_1));
    CFG4 #( .INIT(16'hFFFE) )  \data_out_2_15_i_0_i[1]  (.A(
        \data_out_2_15_i_0_i_4[1]_net_1 ), .B(
        \data_out_2_15_i_0_i_5[1]_net_1 ), .C(
        \data_out_2_15_i_0_i_12[1]_net_1 ), .D(
        \data_out_2_15_i_0_i_11[1]_net_1 ), .Y(N_9));
    CFG3 #( .INIT(8'h02) )  un1_data_out8_36 (.A(\mem_6_[4]_net_1 ), 
        .B(\mem_6__2_i_0_0_a2[2] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_36_net_1));
    SLE \mem_4_[4]  (.D(CoreAPB3_0_APBmslave4_PWDATA[4]), .CLK(
        FCCC_0_GL1), .EN(mem_4__1_sqmuxa), .ALn(un1_data_out8_140_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_4_rs[4] ));
    CFG2 #( .INIT(4'h8) )  mem_3__1_sqmuxa_0_a3_0_a3 (.A(
        mem_14__1_sqmuxa_0_a2_0_a3_0_a2_net_1), .B(
        \mem_3__2_i_0_0_a2[0] ), .Y(mem_3__1_sqmuxa));
    CFG3 #( .INIT(8'hF2) )  un1_data_out8_165 (.A(\mem_2_[5]_net_1 ), 
        .B(\mem_2__2_i_0_0_a2[0] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_165_i));
    SLE un1_data_out8_129_rs (.D(VCC_net_1), .CLK(
        un1_data_out8_123_net_1), .EN(VCC_net_1), .ALn(
        un1_data_out8_129_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(VCC_net_1), .Q(un1_data_out8_129_rs_net_1));
    CFG1 #( .INIT(2'h1) )  un1_data_out8_119_set_RNO (.A(
        un1_data_out8_119_net_1), .Y(un1_data_out8_119_i));
    CFG3 #( .INIT(8'h02) )  un1_data_out8_64 (.A(\mem_8_[2]_net_1 ), 
        .B(mem_8__2_i_0_0_a2[2]), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_64_net_1));
    SLE un1_data_out8_210_rs (.D(VCC_net_1), .CLK(
        un1_data_out8_106_net_1), .EN(VCC_net_1), .ALn(
        un1_data_out8_210_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(VCC_net_1), .Q(un1_data_out8_210_rs_net_1));
    CFG3 #( .INIT(8'hF8) )  \mem_12__RNIL9951[5]  (.A(
        un1_data_out8_21_set_net_1), .B(un1_data_out8_245_rs_net_1), 
        .C(\mem_12_rs[5] ), .Y(\mem_12_[5]_net_1 ));
    SLE un1_data_out8_52_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_7__1_sqmuxa), .ALn(un1_data_out8_52_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_data_out8_52_set_net_1));
    SLE un1_data_out8_207_rs (.D(VCC_net_1), .CLK(
        un1_data_out8_32_net_1), .EN(VCC_net_1), .ALn(
        un1_data_out8_207_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(VCC_net_1), .Q(un1_data_out8_207_rs_net_1));
    CFG3 #( .INIT(8'h02) )  un1_data_out8_52 (.A(\mem_7_[4]_net_1 ), 
        .B(\mem_7__2_i_0_0_a2[1] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_52_net_1));
    CFG3 #( .INIT(8'hF8) )  \mem_14__RNI7A3Q[5]  (.A(
        un1_data_out8_117_set_net_1), .B(un1_data_out8_221_rs_net_1), 
        .C(\mem_14_rs[5] ), .Y(\mem_14_[5]_net_1 ));
    SLE un1_data_out8_147_rs (.D(VCC_net_1), .CLK(
        un1_data_out8_80_net_1), .EN(VCC_net_1), .ALn(
        un1_data_out8_147_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(VCC_net_1), .Q(un1_data_out8_147_rs_net_1));
    SLE \mem_10_[4]  (.D(CoreAPB3_0_APBmslave4_PWDATA[4]), .CLK(
        FCCC_0_GL1), .EN(mem_10__1_sqmuxa), .ALn(un1_data_out8_174_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_10_rs[4] ));
    CFG4 #( .INIT(16'hEAC0) )  \data_out_2_15_i_i_2[2]  (.A(
        \mem_13_[2]_net_1 ), .B(\mem_11_[2]_net_1 ), .C(
        \mem_11__2_i_0_0_a2[2] ), .D(\mem_13__2_i_0_0_a2[0] ), .Y(
        \data_out_2_15_i_i_2[2]_net_1 ));
    SLE un1_data_out8_187_rs (.D(VCC_net_1), .CLK(
        un1_data_out8_12_net_1), .EN(VCC_net_1), .ALn(
        un1_data_out8_187_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(VCC_net_1), .Q(un1_data_out8_187_rs_net_1));
    SLE un1_data_out8_174_rs (.D(VCC_net_1), .CLK(
        un1_data_out8_101_net_1), .EN(VCC_net_1), .ALn(
        un1_data_out8_174_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(VCC_net_1), .Q(un1_data_out8_174_rs_net_1));
    SLE \mem_7_[0]  (.D(CoreAPB3_0_APBmslave4_PWDATA[0]), .CLK(
        FCCC_0_GL1), .EN(mem_7__1_sqmuxa), .ALn(un1_data_out8_179_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_7_rs[0] ));
    SLE un1_data_out8_171_rs (.D(VCC_net_1), .CLK(
        un1_data_out8_36_net_1), .EN(VCC_net_1), .ALn(
        un1_data_out8_171_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(VCC_net_1), .Q(un1_data_out8_171_rs_net_1));
    CFG4 #( .INIT(16'hEAC0) )  \data_out_2_15_i_0_i_0[0]  (.A(
        \mem_10_[0]_net_1 ), .B(\mem_12_[0]_net_1 ), .C(
        \mem_12__2_i_0_0_a2[0] ), .D(\mem_10__2_i_0_0_a2[0] ), .Y(
        \data_out_2_15_i_0_i_0[0]_net_1 ));
    CFG3 #( .INIT(8'h02) )  un1_data_out8_29 (.A(\mem_2_[2]_net_1 ), 
        .B(\mem_2__2_i_0_0_a2[0] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_29_net_1));
    SLE \mem_14_[2]  (.D(CoreAPB3_0_APBmslave4_PWDATA[2]), .CLK(
        FCCC_0_GL1), .EN(mem_14__1_sqmuxa), .ALn(un1_data_out8_218_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_14_rs[2] ));
    SLE \mem_2_[0]  (.D(CoreAPB3_0_APBmslave4_PWDATA[0]), .CLK(
        FCCC_0_GL1), .EN(mem_2__1_sqmuxa), .ALn(un1_data_out8_160_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_2_rs[0] ));
    CFG3 #( .INIT(8'h02) )  un1_data_out8_55 (.A(\mem_3_[7]_net_1 ), 
        .B(\mem_3__2_i_0_0_a2[0] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_55_net_1));
    CFG3 #( .INIT(8'h02) )  un1_data_out8_30 (.A(\mem_6_[1]_net_1 ), 
        .B(\mem_6__2_i_0_0_a2[2] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_30_net_1));
    CFG3 #( .INIT(8'hF2) )  un1_data_out8_220 (.A(\mem_14_[4]_net_1 ), 
        .B(\mem_14__2_i_0_0_a2[2] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_220_i));
    SLE un1_data_out8_65_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_4__1_sqmuxa), .ALn(un1_data_out8_65_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_data_out8_65_set_net_1));
    CFG3 #( .INIT(8'h02) )  un1_data_out8_49 (.A(\mem_3_[4]_net_1 ), 
        .B(\mem_3__2_i_0_0_a2[0] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_49_net_1));
    CFG2 #( .INIT(4'h8) )  mem_7__1_sqmuxa_0_a3_0_a3 (.A(
        mem_14__1_sqmuxa_0_a2_0_a3_0_a2_net_1), .B(
        \mem_7__2_i_0_0_a2[1] ), .Y(mem_7__1_sqmuxa));
    SLE \mem_4_[0]  (.D(CoreAPB3_0_APBmslave4_PWDATA[0]), .CLK(
        FCCC_0_GL1), .EN(mem_4__1_sqmuxa), .ALn(un1_data_out8_136_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_4_rs[0] ));
    CFG3 #( .INIT(8'hF8) )  \mem_3__RNICQ721[7]  (.A(
        un1_data_out8_55_set_net_1), .B(un1_data_out8_135_rs_net_1), 
        .C(\mem_3_rs[7] ), .Y(\mem_3_[7]_net_1 ));
    CFG2 #( .INIT(4'h8) )  \data_out_2_15_i_i_a3_8[6]  (.A(
        \mem_3__2_i_0_0_a2[0] ), .B(\mem_3_[6]_net_1 ), .Y(
        \data_out_2_15_i_i_a3_8[6]_net_1 ));
    SLE \mem_10_[6]  (.D(CoreAPB3_0_APBmslave4_PWDATA[6]), .CLK(
        FCCC_0_GL1), .EN(mem_10__1_sqmuxa), .ALn(un1_data_out8_178_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_10_rs[6] ));
    SLE un1_data_out8_133_rs (.D(VCC_net_1), .CLK(
        un1_data_out8_51_net_1), .EN(VCC_net_1), .ALn(
        un1_data_out8_133_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(VCC_net_1), .Q(un1_data_out8_133_rs_net_1));
    CFG3 #( .INIT(8'h02) )  un1_data_out8_105 (.A(\mem_13_[1]_net_1 ), 
        .B(\mem_13__2_i_0_0_a2[0] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_105_net_1));
    CFG3 #( .INIT(8'h02) )  un1_data_out8_91 (.A(\mem_11_[3]_net_1 ), 
        .B(\mem_11__2_i_0_0_a2[2] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_91_net_1));
    CFG3 #( .INIT(8'hF2) )  un1_data_out8_182 (.A(\mem_11_[0]_net_1 ), 
        .B(\mem_11__2_i_0_0_a2[2] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_182_i));
    CFG1 #( .INIT(2'h1) )  un1_data_out8_65_set_RNO (.A(
        un1_data_out8_65_net_1), .Y(un1_data_out8_65_i));
    CFG3 #( .INIT(8'h02) )  un1_data_out8_54 (.A(\mem_7_[5]_net_1 ), 
        .B(\mem_7__2_i_0_0_a2[1] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_54_net_1));
    CFG4 #( .INIT(16'hFFF8) )  \data_out_2_15_i_i_11[2]  (.A(
        \mem_5__2_i_0_0_a2[0] ), .B(\mem_5_[2]_net_1 ), .C(
        \data_out_2_15_i_i_7[2]_net_1 ), .D(
        \data_out_2_15_i_i_a3_8[2]_net_1 ), .Y(
        \data_out_2_15_i_i_11[2]_net_1 ));
    CFG4 #( .INIT(16'hECA0) )  \data_out_2_15_i_0_i_7[7]  (.A(
        \mem_8_[7]_net_1 ), .B(\mem_0_[7]_net_1 ), .C(
        mem_8__2_i_0_0_a2[2]), .D(mem_0__2_i_0_0_a2[0]), .Y(
        \data_out_2_15_i_0_i_7[7]_net_1 ));
    CFG1 #( .INIT(2'h1) )  un1_data_out8_set_RNO (.A(
        un1_data_out8_net_1), .Y(un1_data_out8_i));
    CFG4 #( .INIT(16'hECA0) )  \data_out_2_15_i_i_5[4]  (.A(
        \mem_6_[4]_net_1 ), .B(\mem_1_[4]_net_1 ), .C(
        \mem_6__2_i_0_0_a2[2] ), .D(\mem_1__2_i_0_0_a2[0] ), .Y(
        \data_out_2_15_i_i_5[4]_net_1 ));
    SLE un1_data_out8_235_rs (.D(VCC_net_1), .CLK(
        un1_data_out8_7_net_1), .EN(VCC_net_1), .ALn(
        un1_data_out8_235_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(VCC_net_1), .Q(un1_data_out8_235_rs_net_1));
    CFG3 #( .INIT(8'hF2) )  un1_data_out8_250 (.A(\mem_15_[3]_net_1 ), 
        .B(\mem_15__2_i_0_0_a2[0] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_250_i));
    CFG3 #( .INIT(8'hF8) )  un1_data_out8_147_rs_RNI3C1M (.A(
        un1_data_out8_80_set_net_1), .B(un1_data_out8_147_rs_net_1), 
        .C(\mem_0_rs[0] ), .Y(\mem_0_[0]_net_1 ));
    CFG3 #( .INIT(8'hF8) )  un1_data_out8_150_rs_RNI9PMB (.A(
        un1_data_out8_86_set_net_1), .B(un1_data_out8_150_rs_net_1), 
        .C(\mem_0_rs[6] ), .Y(\mem_0_[6]_net_1 ));
    CFG3 #( .INIT(8'hF8) )  \mem_2__RNIAMVL[5]  (.A(
        un1_data_out8_35_set_net_1), .B(un1_data_out8_165_rs_net_1), 
        .C(\mem_2_rs[5] ), .Y(\mem_2_[5]_net_1 ));
    SLE un1_data_out8_99_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_10__1_sqmuxa), .ALn(un1_data_out8_99_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_data_out8_99_set_net_1));
    CFG1 #( .INIT(2'h1) )  un1_data_out8_4_set_RNO (.A(
        un1_data_out8_4_net_1), .Y(un1_data_out8_4_i));
    CFG1 #( .INIT(2'h1) )  un1_data_out8_61_set_RNO (.A(
        un1_data_out8_61_net_1), .Y(un1_data_out8_61_i));
    CFG3 #( .INIT(8'hF2) )  un1_data_out8_169 (.A(\mem_6_[3]_net_1 ), 
        .B(\mem_6__2_i_0_0_a2[2] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_169_i));
    SLE un1_data_out8_225_rs (.D(VCC_net_1), .CLK(
        un1_data_out8_50_net_1), .EN(VCC_net_1), .ALn(
        un1_data_out8_225_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(VCC_net_1), .Q(un1_data_out8_225_rs_net_1));
    CFG3 #( .INIT(8'hF8) )  \mem_7__RNIQQ531[1]  (.A(
        un1_data_out8_126_set_net_1), .B(un1_data_out8_181_rs_net_1), 
        .C(\mem_7_rs[1] ), .Y(\mem_7_[1]_net_1 ));
    CFG3 #( .INIT(8'hF2) )  un1_data_out8_240 (.A(\mem_12_[1]_net_1 ), 
        .B(\mem_12__2_i_0_0_a2[0] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_240_i));
    CFG3 #( .INIT(8'hF2) )  un1_data_out8_132 (.A(\mem_3_[4]_net_1 ), 
        .B(\mem_3__2_i_0_0_a2[0] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_132_i));
    CFG1 #( .INIT(2'h1) )  un1_data_out8_5_set_RNO (.A(
        un1_data_out8_5_net_1), .Y(un1_data_out8_5_i));
    CFG3 #( .INIT(8'hF8) )  un1_data_out8_232_rs_RNIP37Q (.A(
        un1_data_out8_93_set_net_1), .B(un1_data_out8_232_rs_net_1), 
        .C(\mem_11_rs[5] ), .Y(\mem_11_[5]_net_1 ));
    CFG3 #( .INIT(8'hF8) )  \mem_3__RNIGG5O[2]  (.A(
        un1_data_out8_125_set_net_1), .B(un1_data_out8_130_rs_net_1), 
        .C(\mem_3_rs[2] ), .Y(\mem_3_[2]_net_1 ));
    SLE un1_data_out8_138_rs (.D(VCC_net_1), .CLK(
        un1_data_out8_4_net_1), .EN(VCC_net_1), .ALn(
        un1_data_out8_138_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(VCC_net_1), .Q(un1_data_out8_138_rs_net_1));
    CFG3 #( .INIT(8'hF8) )  un1_data_out8_42_set_RNI8DHT (.A(
        un1_data_out8_42_set_net_1), .B(un1_data_out8_157_rs_net_1), 
        .C(\mem_1_rs[5] ), .Y(\mem_1_[5]_net_1 ));
    SLE \data_out[4]  (.D(N_15), .CLK(FCCC_0_GL1), .EN(rd_enable), 
        .ALn(MSS_RESET_N_M2F_c), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(
        CoreAPB3_0_APBmslave5_PRDATA[4]));
    CFG4 #( .INIT(16'h0008) )  \WRITE_GEN.mem_9__2_i_0_0_a2[0]  (.A(
        CoreAPB3_0_APBmslave4_PADDR[2]), .B(
        CoreAPB3_0_APBmslave4_PADDR[5]), .C(
        CoreAPB3_0_APBmslave4_PADDR[4]), .D(
        CoreAPB3_0_APBmslave4_PADDR[3]), .Y(\mem_9__2_i_0_0_a2[0] ));
    SLE un1_data_out8_62_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_15__1_sqmuxa), .ALn(un1_data_out8_62_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_data_out8_62_set_net_1));
    CFG1 #( .INIT(2'h1) )  un1_data_out8_35_set_RNO (.A(
        un1_data_out8_35_net_1), .Y(un1_data_out8_35_i));
    SLE un1_data_out8_91_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_11__1_sqmuxa), .ALn(un1_data_out8_91_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_data_out8_91_set_net_1));
    CFG3 #( .INIT(8'hF2) )  un1_data_out8_208 (.A(\mem_13_[0]_net_1 ), 
        .B(\mem_13__2_i_0_0_a2[0] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_208_i));
    CFG1 #( .INIT(2'h1) )  un1_data_out8_55_set_RNO (.A(
        un1_data_out8_55_net_1), .Y(un1_data_out8_55_i));
    CFG3 #( .INIT(8'h02) )  un1_data_out8_1 (.A(\mem_7_[7]_net_1 ), .B(
        \mem_7__2_i_0_0_a2[1] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_1_net_1));
    SLE un1_data_out8_196_rs (.D(VCC_net_1), .CLK(
        un1_data_out8_75_net_1), .EN(VCC_net_1), .ALn(
        un1_data_out8_196_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(VCC_net_1), .Q(un1_data_out8_196_rs_net_1));
    CFG3 #( .INIT(8'h02) )  un1_data_out8_111 (.A(\mem_13_[7]_net_1 ), 
        .B(\mem_13__2_i_0_0_a2[0] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_111_net_1));
    CFG1 #( .INIT(2'h1) )  un1_data_out8_74_set_RNO (.A(
        un1_data_out8_74_net_1), .Y(un1_data_out8_74_i));
    CFG3 #( .INIT(8'hF2) )  un1_data_out8_222 (.A(\mem_14_[6]_net_1 ), 
        .B(\mem_14__2_i_0_0_a2[2] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_222_i));
    SLE un1_data_out8_128_rs (.D(VCC_net_1), .CLK(
        un1_data_out8_121_net_1), .EN(VCC_net_1), .ALn(
        un1_data_out8_128_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(VCC_net_1), .Q(un1_data_out8_128_rs_net_1));
    CFG4 #( .INIT(16'hFFFE) )  \data_out_2_15_i_i_12[5]  (.A(
        \data_out_2_15_i_i_2[5]_net_1 ), .B(
        \data_out_2_15_i_i_1[5]_net_1 ), .C(
        \data_out_2_15_i_i_3[5]_net_1 ), .D(
        \data_out_2_15_i_i_0[5]_net_1 ), .Y(
        \data_out_2_15_i_i_12[5]_net_1 ));
    SLE \data_out[3]  (.D(N_7), .CLK(FCCC_0_GL1), .EN(rd_enable), .ALn(
        MSS_RESET_N_M2F_c), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(
        CoreAPB3_0_APBmslave5_PRDATA[3]));
    SLE un1_data_out8_156_rs (.D(VCC_net_1), .CLK(
        un1_data_out8_40_net_1), .EN(VCC_net_1), .ALn(
        un1_data_out8_156_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(VCC_net_1), .Q(un1_data_out8_156_rs_net_1));
    CFG3 #( .INIT(8'hF8) )  un1_data_out8_46_set_RNIG5G01 (.A(
        un1_data_out8_46_set_net_1), .B(un1_data_out8_159_rs_net_1), 
        .C(\mem_1_rs[7] ), .Y(\mem_1_[7]_net_1 ));
    CFG1 #( .INIT(2'h1) )  un1_data_out8_45_set_RNO (.A(
        un1_data_out8_45_net_1), .Y(un1_data_out8_45_i));
    CFG1 #( .INIT(2'h1) )  un1_data_out8_112_set_RNO (.A(
        un1_data_out8_112_net_1), .Y(un1_data_out8_112_i));
    SLE un1_data_out8_27_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_2__1_sqmuxa), .ALn(un1_data_out8_27_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_data_out8_27_set_net_1));
    SLE un1_data_out8_87_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_0__1_sqmuxa), .ALn(un1_data_out8_87_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_data_out8_87_set_net_1));
    CFG1 #( .INIT(2'h1) )  un1_data_out8_31_set_RNO (.A(
        un1_data_out8_31_net_1), .Y(un1_data_out8_31_i));
    CFG1 #( .INIT(2'h1) )  un1_data_out8_51_set_RNO (.A(
        un1_data_out8_51_net_1), .Y(un1_data_out8_51_i));
    SLE un1_data_out8_115_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_14__1_sqmuxa), .ALn(un1_data_out8_115_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_data_out8_115_set_net_1));
    SLE un1_data_out8_216_rs (.D(VCC_net_1), .CLK(
        un1_data_out8_112_net_1), .EN(VCC_net_1), .ALn(
        un1_data_out8_216_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(VCC_net_1), .Q(un1_data_out8_216_rs_net_1));
    CFG4 #( .INIT(16'hEAC0) )  \data_out_2_15_i_i_0[6]  (.A(
        \mem_10_[6]_net_1 ), .B(\mem_12_[6]_net_1 ), .C(
        \mem_12__2_i_0_0_a2[0] ), .D(\mem_10__2_i_0_0_a2[0] ), .Y(
        \data_out_2_15_i_i_0[6]_net_1 ));
    CFG3 #( .INIT(8'hF2) )  un1_data_out8_187 (.A(\mem_5_[0]_net_1 ), 
        .B(\mem_5__2_i_0_0_a2[0] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_187_i));
    SLE un1_data_out8_125_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_3__1_sqmuxa), .ALn(un1_data_out8_125_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_data_out8_125_set_net_1));
    CFG3 #( .INIT(8'hF2) )  un1_data_out8_252 (.A(\mem_15_[5]_net_1 ), 
        .B(\mem_15__2_i_0_0_a2[0] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_252_i));
    CFG3 #( .INIT(8'hF8) )  un1_data_out8_241_rs_RNIDGQV (.A(
        un1_data_out8_66_set_net_1), .B(un1_data_out8_241_rs_net_1), 
        .C(\mem_8_rs[3] ), .Y(\mem_8_[3]_net_1 ));
    CFG3 #( .INIT(8'h02) )  un1_data_out8_116 (.A(\mem_14_[4]_net_1 ), 
        .B(\mem_14__2_i_0_0_a2[2] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_116_net_1));
    CFG3 #( .INIT(8'hF2) )  un1_data_out8_172 (.A(\mem_10_[3]_net_1 ), 
        .B(\mem_10__2_i_0_0_a2[0] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_172_i));
    SLE un1_data_out8_199_rs (.D(VCC_net_1), .CLK(
        un1_data_out8_24_net_1), .EN(VCC_net_1), .ALn(
        un1_data_out8_199_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(VCC_net_1), .Q(un1_data_out8_199_rs_net_1));
    CFG1 #( .INIT(2'h1) )  un1_data_out8_41_set_RNO (.A(
        un1_data_out8_41_net_1), .Y(un1_data_out8_41_i));
    CFG3 #( .INIT(8'h02) )  un1_data_out8_109 (.A(\mem_13_[5]_net_1 ), 
        .B(\mem_13__2_i_0_0_a2[0] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_109_net_1));
    SLE un1_data_out8_105_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_13__1_sqmuxa), .ALn(un1_data_out8_105_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_data_out8_105_set_net_1));
    CFG3 #( .INIT(8'hF2) )  un1_data_out8_168 (.A(\mem_10_[1]_net_1 ), 
        .B(\mem_10__2_i_0_0_a2[0] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_168_i));
    SLE \mem_8_[2]  (.D(CoreAPB3_0_APBmslave4_PWDATA[2]), .CLK(
        FCCC_0_GL1), .EN(mem_8__1_sqmuxa), .ALn(un1_data_out8_239_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_8_rs[2] ));
    CFG4 #( .INIT(16'h0010) )  \WRITE_GEN.mem_4__2_i_0_0_a2[0]  (.A(
        CoreAPB3_0_APBmslave4_PADDR[2]), .B(
        CoreAPB3_0_APBmslave4_PADDR[5]), .C(
        CoreAPB3_0_APBmslave4_PADDR[4]), .D(
        CoreAPB3_0_APBmslave4_PADDR[3]), .Y(\mem_4__2_i_0_0_a2[0] ));
    SLE un1_data_out8_167_rs (.D(VCC_net_1), .CLK(
        un1_data_out8_39_net_1), .EN(VCC_net_1), .ALn(
        un1_data_out8_167_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(VCC_net_1), .Q(un1_data_out8_167_rs_net_1));
    CFG3 #( .INIT(8'h02) )  un1_data_out8_16 (.A(\mem_12_[0]_net_1 ), 
        .B(\mem_12__2_i_0_0_a2[0] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_16_net_1));
    SLE un1_data_out8_56_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_15__1_sqmuxa), .ALn(un1_data_out8_56_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_data_out8_56_set_net_1));
    SLE \mem_6_[7]  (.D(CoreAPB3_0_APBmslave4_PWDATA[7]), .CLK(
        FCCC_0_GL1), .EN(mem_6__1_sqmuxa), .ALn(un1_data_out8_177_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_6_rs[7] ));
    SLE un1_data_out8_159_rs (.D(VCC_net_1), .CLK(
        un1_data_out8_46_net_1), .EN(VCC_net_1), .ALn(
        un1_data_out8_159_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(VCC_net_1), .Q(un1_data_out8_159_rs_net_1));
    CFG3 #( .INIT(8'hF8) )  un1_data_out8_192_rs_RNIFTFT (.A(
        un1_data_out8_73_set_net_1), .B(un1_data_out8_192_rs_net_1), 
        .C(\mem_9_rs[1] ), .Y(\mem_9_[1]_net_1 ));
    CFG1 #( .INIT(2'h1) )  un1_data_out8_69_set_RNO (.A(
        un1_data_out8_69_net_1), .Y(un1_data_out8_69_i));
    SLE un1_data_out8_77_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_9__1_sqmuxa), .ALn(un1_data_out8_77_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_data_out8_77_set_net_1));
    CFG4 #( .INIT(16'hEAC0) )  \data_out_2_15_i_0_i_0[1]  (.A(
        \mem_10_[1]_net_1 ), .B(\mem_12_[1]_net_1 ), .C(
        \mem_12__2_i_0_0_a2[0] ), .D(\mem_10__2_i_0_0_a2[0] ), .Y(
        \data_out_2_15_i_0_i_0[1]_net_1 ));
    CFG1 #( .INIT(2'h1) )  un1_data_out8_77_set_RNO (.A(
        un1_data_out8_77_net_1), .Y(un1_data_out8_77_i));
    SLE \mem_14_[7]  (.D(CoreAPB3_0_APBmslave4_PWDATA[7]), .CLK(
        FCCC_0_GL1), .EN(mem_14__1_sqmuxa), .ALn(un1_data_out8_223_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_14_rs[7] ));
    CFG3 #( .INIT(8'hF8) )  \mem_2__RNI2U0J[3]  (.A(
        un1_data_out8_31_set_net_1), .B(un1_data_out8_163_rs_net_1), 
        .C(\mem_2_rs[3] ), .Y(\mem_2_[3]_net_1 ));
    CFG3 #( .INIT(8'hF2) )  un1_data_out8_242 (.A(\mem_12_[2]_net_1 ), 
        .B(\mem_12__2_i_0_0_a2[0] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_242_i));
    CFG1 #( .INIT(2'h1) )  un1_data_out8_3_set_RNO (.A(
        un1_data_out8_3_net_1), .Y(un1_data_out8_3_i));
    SLE \mem_6_[5]  (.D(CoreAPB3_0_APBmslave4_PWDATA[5]), .CLK(
        FCCC_0_GL1), .EN(mem_6__1_sqmuxa), .ALn(un1_data_out8_173_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_6_rs[5] ));
    SLE un1_data_out8_135_rs (.D(VCC_net_1), .CLK(
        un1_data_out8_55_net_1), .EN(VCC_net_1), .ALn(
        un1_data_out8_135_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(VCC_net_1), .Q(un1_data_out8_135_rs_net_1));
    SLE un1_data_out8_146_rs (.D(VCC_net_1), .CLK(
        un1_data_out8_83_net_1), .EN(VCC_net_1), .ALn(
        un1_data_out8_146_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(VCC_net_1), .Q(un1_data_out8_146_rs_net_1));
    CFG3 #( .INIT(8'hF2) )  un1_data_out8_137 (.A(\mem_4_[1]_net_1 ), 
        .B(\mem_4__2_i_0_0_a2[0] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_137_i));
    SLE \mem_15_[5]  (.D(CoreAPB3_0_APBmslave4_PWDATA[5]), .CLK(
        FCCC_0_GL1), .EN(mem_15__1_sqmuxa), .ALn(un1_data_out8_252_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_15_rs[5] ));
    SLE un1_data_out8_186_rs (.D(VCC_net_1), .CLK(
        un1_data_out8_70_net_1), .EN(VCC_net_1), .ALn(
        un1_data_out8_186_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(VCC_net_1), .Q(un1_data_out8_186_rs_net_1));
    SLE \mem_0_[7]  (.D(CoreAPB3_0_APBmslave4_PWDATA[7]), .CLK(
        FCCC_0_GL1), .EN(mem_0__1_sqmuxa), .ALn(un1_data_out8_151_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_0_rs[7] ));
    CFG3 #( .INIT(8'hF8) )  un1_data_out8_104_set_RNI2T9U (.A(
        un1_data_out8_104_set_net_1), .B(un1_data_out8_208_rs_net_1), 
        .C(\mem_13_rs[0] ), .Y(\mem_13_[0]_net_1 ));
    CFG4 #( .INIT(16'hECA0) )  \data_out_2_15_i_i_7[6]  (.A(
        \mem_8_[6]_net_1 ), .B(\mem_0_[6]_net_1 ), .C(
        mem_8__2_i_0_0_a2[2]), .D(mem_0__2_i_0_0_a2[0]), .Y(
        \data_out_2_15_i_i_7[6]_net_1 ));
    SLE \mem_0_[5]  (.D(CoreAPB3_0_APBmslave4_PWDATA[5]), .CLK(
        FCCC_0_GL1), .EN(mem_0__1_sqmuxa), .ALn(un1_data_out8_149_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_0_rs[5] ));
    SLE \mem_15_[1]  (.D(CoreAPB3_0_APBmslave4_PWDATA[1]), .CLK(
        FCCC_0_GL1), .EN(mem_15__1_sqmuxa), .ALn(un1_data_out8_248_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_15_rs[1] ));
    CFG1 #( .INIT(2'h1) )  un1_data_out8_39_set_RNO (.A(
        un1_data_out8_39_net_1), .Y(un1_data_out8_39_i));
    CFG2 #( .INIT(4'h8) )  mem_15__1_sqmuxa_0_a3_0_a3 (.A(
        mem_14__1_sqmuxa_0_a2_0_a3_0_a2_net_1), .B(
        \mem_15__2_i_0_0_a2[0] ), .Y(mem_15__1_sqmuxa));
    SLE un1_data_out8_238_rs (.D(VCC_net_1), .CLK(
        un1_data_out8_16_net_1), .EN(VCC_net_1), .ALn(
        un1_data_out8_238_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(VCC_net_1), .Q(un1_data_out8_238_rs_net_1));
    SLE un1_data_out8_209_rs (.D(VCC_net_1), .CLK(
        un1_data_out8_105_net_1), .EN(VCC_net_1), .ALn(
        un1_data_out8_209_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(VCC_net_1), .Q(un1_data_out8_209_rs_net_1));
    SLE un1_data_out8_1_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_7__1_sqmuxa), .ALn(un1_data_out8_1_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_data_out8_1_set_net_1));
    CFG3 #( .INIT(8'h02) )  un1_data_out8_9 (.A(\mem_1_[0]_net_1 ), .B(
        \mem_1__2_i_0_0_a2[0] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_9_net_1));
    SLE un1_data_out8_25_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_2__1_sqmuxa), .ALn(un1_data_out8_25_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_data_out8_25_set_net_1));
    SLE un1_data_out8_85_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_0__1_sqmuxa), .ALn(un1_data_out8_85_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_data_out8_85_set_net_1));
    CFG1 #( .INIT(2'h1) )  un1_data_out8_59_set_RNO (.A(
        un1_data_out8_59_net_1), .Y(un1_data_out8_59_i));
    SLE un1_data_out8_149_rs (.D(VCC_net_1), .CLK(
        un1_data_out8_85_net_1), .EN(VCC_net_1), .ALn(
        un1_data_out8_149_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(VCC_net_1), .Q(un1_data_out8_149_rs_net_1));
    SLE un1_data_out8_30_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_6__1_sqmuxa), .ALn(un1_data_out8_30_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_data_out8_30_set_net_1));
    CFG3 #( .INIT(8'h02) )  un1_data_out8_108 (.A(\mem_13_[4]_net_1 ), 
        .B(\mem_13__2_i_0_0_a2[0] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_108_net_1));
    SLE un1_data_out8_93_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_11__1_sqmuxa), .ALn(un1_data_out8_93_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_data_out8_93_set_net_1));
    CFG3 #( .INIT(8'h02) )  un1_data_out8_10 (.A(\mem_4_[7]_net_1 ), 
        .B(\mem_4__2_i_0_0_a2[0] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_10_net_1));
    SLE un1_data_out8_189_rs (.D(VCC_net_1), .CLK(
        un1_data_out8_14_net_1), .EN(VCC_net_1), .ALn(
        un1_data_out8_189_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(VCC_net_1), .Q(un1_data_out8_189_rs_net_1));
    CFG3 #( .INIT(8'h02) )  un1_data_out8_61 (.A(\mem_15_[4]_net_1 ), 
        .B(\mem_15__2_i_0_0_a2[0] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_61_net_1));
    SLE \data_out[6]  (.D(N_19), .CLK(FCCC_0_GL1), .EN(rd_enable), 
        .ALn(MSS_RESET_N_M2F_c), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(
        CoreAPB3_0_APBmslave5_PRDATA[6]));
    CFG1 #( .INIT(2'h1) )  un1_data_out8_49_set_RNO (.A(
        un1_data_out8_49_net_1), .Y(un1_data_out8_49_i));
    SLE un1_data_out8_193_rs (.D(VCC_net_1), .CLK(
        un1_data_out8_41_net_1), .EN(VCC_net_1), .ALn(
        un1_data_out8_193_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(VCC_net_1), .Q(un1_data_out8_193_rs_net_1));
    SLE \data_out[0]  (.D(N_11), .CLK(FCCC_0_GL1), .EN(rd_enable), 
        .ALn(MSS_RESET_N_M2F_c), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(
        CoreAPB3_0_APBmslave5_PRDATA[0]));
    SLE un1_data_out8_228_rs (.D(VCC_net_1), .CLK(
        un1_data_out8_91_net_1), .EN(VCC_net_1), .ALn(
        un1_data_out8_228_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(VCC_net_1), .Q(un1_data_out8_228_rs_net_1));
    CFG3 #( .INIT(8'hF8) )  un1_data_out8_211_rs_RNI2RC71 (.A(
        un1_data_out8_107_set_net_1), .B(un1_data_out8_211_rs_net_1), 
        .C(\mem_13_rs[3] ), .Y(\mem_13_[3]_net_1 ));
    CFG3 #( .INIT(8'hF2) )  un1_data_out8_177 (.A(\mem_6_[7]_net_1 ), 
        .B(\mem_6__2_i_0_0_a2[2] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_177_i));
    CFG1 #( .INIT(2'h1) )  un1_data_out8_76_set_RNO (.A(
        un1_data_out8_76_net_1), .Y(un1_data_out8_76_i));
    SLE un1_data_out8_153_rs (.D(VCC_net_1), .CLK(
        un1_data_out8_11_net_1), .EN(VCC_net_1), .ALn(
        un1_data_out8_153_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(VCC_net_1), .Q(un1_data_out8_153_rs_net_1));
    SLE un1_data_out8_94_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_11__1_sqmuxa), .ALn(un1_data_out8_94_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_data_out8_94_set_net_1));
    CFG1 #( .INIT(2'h1) )  un1_data_out8_14_set_RNO (.A(
        un1_data_out8_14_net_1), .Y(un1_data_out8_14_i));
    SLE un1_data_out8_75_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_9__1_sqmuxa), .ALn(un1_data_out8_75_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_data_out8_75_set_net_1));
    CFG3 #( .INIT(8'hF8) )  un1_data_out8_44_set_RNICP0N (.A(
        un1_data_out8_44_set_net_1), .B(un1_data_out8_158_rs_net_1), 
        .C(\mem_1_rs[6] ), .Y(\mem_1_[6]_net_1 ));
    CFG4 #( .INIT(16'hECA0) )  \data_out_2_15_i_0_i_7[0]  (.A(
        \mem_8_[0]_net_1 ), .B(\mem_0_[0]_net_1 ), .C(
        mem_8__2_i_0_0_a2[2]), .D(mem_0__2_i_0_0_a2[0]), .Y(
        \data_out_2_15_i_0_i_7[0]_net_1 ));
    CFG3 #( .INIT(8'h02) )  un1_data_out8_96 (.A(\mem_10_[3]_net_1 ), 
        .B(\mem_10__2_i_0_0_a2[0] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_96_net_1));
    CFG3 #( .INIT(8'hF8) )  un1_data_out8_65_set_RNI7LEV (.A(
        un1_data_out8_65_set_net_1), .B(un1_data_out8_140_rs_net_1), 
        .C(\mem_4_rs[4] ), .Y(\mem_4_[4]_net_1 ));
    SLE \mem_8_[1]  (.D(CoreAPB3_0_APBmslave4_PWDATA[1]), .CLK(
        FCCC_0_GL1), .EN(mem_8__1_sqmuxa), .ALn(un1_data_out8_237_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_8_rs[1] ));
    SLE \mem_1_[7]  (.D(CoreAPB3_0_APBmslave4_PWDATA[7]), .CLK(
        FCCC_0_GL1), .EN(mem_1__1_sqmuxa), .ALn(un1_data_out8_159_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_1_rs[7] ));
    SLE un1_data_out8_255_rs (.D(VCC_net_1), .CLK(
        un1_data_out8_61_net_1), .EN(VCC_net_1), .ALn(
        un1_data_out8_255_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(VCC_net_1), .Q(un1_data_out8_255_rs_net_1));
    SLE un1_data_out8_66_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_8__1_sqmuxa), .ALn(un1_data_out8_66_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_data_out8_66_set_net_1));
    SLE \mem_9_[7]  (.D(CoreAPB3_0_APBmslave4_PWDATA[7]), .CLK(
        FCCC_0_GL1), .EN(mem_9__1_sqmuxa), .ALn(un1_data_out8_204_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_9_rs[7] ));
    CFG3 #( .INIT(8'hF2) )  un1_data_out8_225 (.A(\mem_7_[3]_net_1 ), 
        .B(\mem_7__2_i_0_0_a2[1] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_225_i));
    CFG4 #( .INIT(16'hFFFE) )  \data_out_2_15_i_0_i_12[3]  (.A(
        \data_out_2_15_i_0_i_2[3]_net_1 ), .B(
        \data_out_2_15_i_0_i_1[3]_net_1 ), .C(
        \data_out_2_15_i_0_i_3[3]_net_1 ), .D(
        \data_out_2_15_i_0_i_0[3]_net_1 ), .Y(
        \data_out_2_15_i_0_i_12[3]_net_1 ));
    SLE un1_data_out8_5_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_8__1_sqmuxa), .ALn(un1_data_out8_5_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_data_out8_5_set_net_1));
    CFG4 #( .INIT(16'hFFFE) )  \data_out_2_15_i_0_i_12[7]  (.A(
        \data_out_2_15_i_0_i_2[7]_net_1 ), .B(
        \data_out_2_15_i_0_i_1[7]_net_1 ), .C(
        \data_out_2_15_i_0_i_3[7]_net_1 ), .D(
        \data_out_2_15_i_0_i_0[7]_net_1 ), .Y(
        \data_out_2_15_i_0_i_12[7]_net_1 ));
    SLE \mem_1_[5]  (.D(CoreAPB3_0_APBmslave4_PWDATA[5]), .CLK(
        FCCC_0_GL1), .EN(mem_1__1_sqmuxa), .ALn(un1_data_out8_157_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_1_rs[5] ));
    CFG1 #( .INIT(2'h1) )  un1_data_out8_84_set_RNO (.A(
        un1_data_out8_84_net_1), .Y(un1_data_out8_84_i));
    CFG3 #( .INIT(8'h02) )  un1_data_out8_82 (.A(\mem_0_[2]_net_1 ), 
        .B(mem_0__2_i_0_0_a2[0]), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_82_net_1));
    CFG3 #( .INIT(8'hF8) )  un1_data_out8_23_set_RNIRPRV (.A(
        un1_data_out8_23_set_net_1), .B(un1_data_out8_247_rs_net_1), 
        .C(\mem_12_rs[7] ), .Y(\mem_12_[7]_net_1 ));
    CFG3 #( .INIT(8'hF8) )  un1_data_out8_186_rs_RNIJQTS (.A(
        un1_data_out8_70_set_net_1), .B(un1_data_out8_186_rs_net_1), 
        .C(\mem_8_rs[6] ), .Y(\mem_8_[6]_net_1 ));
    SLE \mem_9_[5]  (.D(CoreAPB3_0_APBmslave4_PWDATA[5]), .CLK(
        FCCC_0_GL1), .EN(mem_9__1_sqmuxa), .ALn(un1_data_out8_200_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_9_rs[5] ));
    CFG4 #( .INIT(16'hEAC0) )  \data_out_2_15_i_i_3[6]  (.A(
        \mem_15_[6]_net_1 ), .B(\mem_7_[6]_net_1 ), .C(
        \mem_7__2_i_0_0_a2[1] ), .D(\mem_15__2_i_0_0_a2[0] ), .Y(
        \data_out_2_15_i_i_3[6]_net_1 ));
    SLE un1_data_out8_22_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_12__1_sqmuxa), .ALn(un1_data_out8_22_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_data_out8_22_set_net_1));
    SLE un1_data_out8_82_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_0__1_sqmuxa), .ALn(un1_data_out8_82_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_data_out8_82_set_net_1));
    SLE un1_data_out8_198_rs (.D(VCC_net_1), .CLK(
        un1_data_out8_76_net_1), .EN(VCC_net_1), .ALn(
        un1_data_out8_198_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(VCC_net_1), .Q(un1_data_out8_198_rs_net_1));
    CFG3 #( .INIT(8'h02) )  un1_data_out8_124 (.A(\mem_7_[0]_net_1 ), 
        .B(\mem_7__2_i_0_0_a2[1] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_124_net_1));
    SLE un1_data_out8_158_rs (.D(VCC_net_1), .CLK(
        un1_data_out8_44_net_1), .EN(VCC_net_1), .ALn(
        un1_data_out8_158_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(VCC_net_1), .Q(un1_data_out8_158_rs_net_1));
    CFG3 #( .INIT(8'hF2) )  un1_data_out8_255 (.A(\mem_15_[4]_net_1 ), 
        .B(\mem_15__2_i_0_0_a2[0] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_255_i));
    CFG3 #( .INIT(8'h02) )  un1_data_out8_51 (.A(\mem_3_[5]_net_1 ), 
        .B(\mem_3__2_i_0_0_a2[0] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_51_net_1));
    SLE un1_data_out8_177_rs (.D(VCC_net_1), .CLK(
        un1_data_out8_122_net_1), .EN(VCC_net_1), .ALn(
        un1_data_out8_177_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(VCC_net_1), .Q(un1_data_out8_177_rs_net_1));
    CFG3 #( .INIT(8'hF8) )  \mem_6__RNIGGAL[5]  (.A(
        un1_data_out8_38_set_net_1), .B(un1_data_out8_173_rs_net_1), 
        .C(\mem_6_rs[5] ), .Y(\mem_6_[5]_net_1 ));
    SLE un1_data_out8_143_rs (.D(VCC_net_1), .CLK(
        un1_data_out8_8_net_1), .EN(VCC_net_1), .ALn(
        un1_data_out8_143_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(VCC_net_1), .Q(un1_data_out8_143_rs_net_1));
    SLE un1_data_out8_234_rs (.D(VCC_net_1), .CLK(
        un1_data_out8_94_net_1), .EN(VCC_net_1), .ALn(
        un1_data_out8_234_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(VCC_net_1), .Q(un1_data_out8_234_rs_net_1));
    CFG1 #( .INIT(2'h1) )  un1_data_out8_17_set_RNO (.A(
        un1_data_out8_17_net_1), .Y(un1_data_out8_17_i));
    CFG3 #( .INIT(8'hF8) )  \mem_12__RNII1001[4]  (.A(
        un1_data_out8_20_set_net_1), .B(un1_data_out8_244_rs_net_1), 
        .C(\mem_12_rs[4] ), .Y(\mem_12_[4]_net_1 ));
    SLE \mem_12_[4]  (.D(CoreAPB3_0_APBmslave4_PWDATA[4]), .CLK(
        FCCC_0_GL1), .EN(mem_12__1_sqmuxa), .ALn(un1_data_out8_244_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_12_rs[4] ));
    SLE \mem_10_[3]  (.D(CoreAPB3_0_APBmslave4_PWDATA[3]), .CLK(
        FCCC_0_GL1), .EN(mem_10__1_sqmuxa), .ALn(un1_data_out8_172_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_10_rs[3] ));
    CFG3 #( .INIT(8'h02) )  un1_data_out8_85 (.A(\mem_0_[5]_net_1 ), 
        .B(mem_0__2_i_0_0_a2[0]), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_85_net_1));
    CFG1 #( .INIT(2'h1) )  un1_data_out8_114_set_RNO (.A(
        un1_data_out8_114_net_1), .Y(un1_data_out8_114_i));
    SLE un1_data_out8_183_rs (.D(VCC_net_1), .CLK(
        un1_data_out8_48_net_1), .EN(VCC_net_1), .ALn(
        un1_data_out8_183_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(VCC_net_1), .Q(un1_data_out8_183_rs_net_1));
    CFG4 #( .INIT(16'h0400) )  \WRITE_GEN.mem_10__2_i_0_0_a2[0]  (.A(
        CoreAPB3_0_APBmslave4_PADDR[2]), .B(
        CoreAPB3_0_APBmslave4_PADDR[5]), .C(
        CoreAPB3_0_APBmslave4_PADDR[4]), .D(
        CoreAPB3_0_APBmslave4_PADDR[3]), .Y(\mem_10__2_i_0_0_a2[0] ));
    CFG4 #( .INIT(16'hECA0) )  \data_out_2_15_i_0_i_7[3]  (.A(
        \mem_8_[3]_net_1 ), .B(\mem_0_[3]_net_1 ), .C(
        mem_8__2_i_0_0_a2[2]), .D(mem_0__2_i_0_0_a2[0]), .Y(
        \data_out_2_15_i_0_i_7[3]_net_1 ));
    CFG4 #( .INIT(16'hEAC0) )  \data_out_2_15_i_i_4[4]  (.A(
        \mem_4_[4]_net_1 ), .B(\mem_2_[4]_net_1 ), .C(
        \mem_2__2_i_0_0_a2[0] ), .D(\mem_4__2_i_0_0_a2[0] ), .Y(
        \data_out_2_15_i_i_4[4]_net_1 ));
    CFG3 #( .INIT(8'h02) )  un1_data_out8_72 (.A(\mem_9_[0]_net_1 ), 
        .B(\mem_9__2_i_0_0_a2[0] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_72_net_1));
    CFG3 #( .INIT(8'hF2) )  un1_data_out8_154 (.A(\mem_1_[2]_net_1 ), 
        .B(\mem_1__2_i_0_0_a2[0] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_154_i));
    SLE un1_data_out8_245_rs (.D(VCC_net_1), .CLK(
        un1_data_out8_21_net_1), .EN(VCC_net_1), .ALn(
        un1_data_out8_245_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(VCC_net_1), .Q(un1_data_out8_245_rs_net_1));
    CFG3 #( .INIT(8'hF2) )  un1_data_out8_161 (.A(\mem_2_[1]_net_1 ), 
        .B(\mem_2__2_i_0_0_a2[0] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_161_i));
    CFG3 #( .INIT(8'hF2) )  un1_data_out8_245 (.A(\mem_12_[5]_net_1 ), 
        .B(\mem_12__2_i_0_0_a2[0] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_245_i));
    SLE \mem_3_[3]  (.D(CoreAPB3_0_APBmslave4_PWDATA[3]), .CLK(
        FCCC_0_GL1), .EN(mem_3__1_sqmuxa), .ALn(un1_data_out8_131_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_3_rs[3] ));
    SLE un1_data_out8_72_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_9__1_sqmuxa), .ALn(un1_data_out8_72_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_data_out8_72_set_net_1));
    CFG3 #( .INIT(8'hF2) )  un1_data_out8_234 (.A(\mem_11_[6]_net_1 ), 
        .B(\mem_11__2_i_0_0_a2[2] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_234_i));
    CFG3 #( .INIT(8'h02) )  un1_data_out8_90 (.A(\mem_11_[2]_net_1 ), 
        .B(\mem_11__2_i_0_0_a2[2] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_90_net_1));
    CFG3 #( .INIT(8'hF8) )  un1_data_out8_191_rs_RNI8SLS (.A(
        un1_data_out8_43_set_net_1), .B(un1_data_out8_191_rs_net_1), 
        .C(\mem_5_rs[2] ), .Y(\mem_5_[2]_net_1 ));
    SLE un1_data_out8_224_rs (.D(VCC_net_1), .CLK(
        un1_data_out8_89_net_1), .EN(VCC_net_1), .ALn(
        un1_data_out8_224_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(VCC_net_1), .Q(un1_data_out8_224_rs_net_1));
    CFG1 #( .INIT(2'h1) )  un1_data_out8_87_set_RNO (.A(
        un1_data_out8_87_net_1), .Y(un1_data_out8_87_i));
    CFG3 #( .INIT(8'hF8) )  un1_data_out8_148_rs_RNIC3TN (.A(
        un1_data_out8_84_set_net_1), .B(un1_data_out8_148_rs_net_1), 
        .C(\mem_0_rs[4] ), .Y(\mem_0_[4]_net_1 ));
    SLE \mem_13_[2]  (.D(CoreAPB3_0_APBmslave4_PWDATA[2]), .CLK(
        FCCC_0_GL1), .EN(mem_13__1_sqmuxa), .ALn(un1_data_out8_210_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_13_rs[2] ));
    CFG3 #( .INIT(8'hF2) )  un1_data_out8_210 (.A(\mem_13_[2]_net_1 ), 
        .B(\mem_13__2_i_0_0_a2[0] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_210_i));
    CFG3 #( .INIT(8'h02) )  un1_data_out8_84 (.A(\mem_0_[4]_net_1 ), 
        .B(mem_0__2_i_0_0_a2[0]), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_84_net_1));
    SLE un1_data_out8_166_rs (.D(VCC_net_1), .CLK(
        un1_data_out8_37_net_1), .EN(VCC_net_1), .ALn(
        un1_data_out8_166_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(VCC_net_1), .Q(un1_data_out8_166_rs_net_1));
    CFG3 #( .INIT(8'hF2) )  un1_data_out8_192 (.A(\mem_9_[1]_net_1 ), 
        .B(\mem_9__2_i_0_0_a2[0] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_192_i));
    CFG4 #( .INIT(16'h8000) )  \WRITE_GEN.mem_15__2_i_0_0_a2[0]  (.A(
        CoreAPB3_0_APBmslave4_PADDR[2]), .B(
        CoreAPB3_0_APBmslave4_PADDR[5]), .C(
        CoreAPB3_0_APBmslave4_PADDR[4]), .D(
        CoreAPB3_0_APBmslave4_PADDR[3]), .Y(\mem_15__2_i_0_0_a2[0] ));
    SLE un1_data_out8_59_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_15__1_sqmuxa), .ALn(un1_data_out8_59_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_data_out8_59_set_net_1));
    CFG3 #( .INIT(8'hF2) )  un1_data_out8_144 (.A(\mem_0_[1]_net_1 ), 
        .B(mem_0__2_i_0_0_a2[0]), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_144_i));
    SLE un1_data_out8_98_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_10__1_sqmuxa), .ALn(un1_data_out8_98_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_data_out8_98_set_net_1));
    SLE \mem_12_[6]  (.D(CoreAPB3_0_APBmslave4_PWDATA[6]), .CLK(
        FCCC_0_GL1), .EN(mem_12__1_sqmuxa), .ALn(un1_data_out8_246_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_12_rs[6] ));
    CFG3 #( .INIT(8'h02) )  un1_data_out8_75 (.A(\mem_9_[3]_net_1 ), 
        .B(\mem_9__2_i_0_0_a2[0] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_75_net_1));
    CFG3 #( .INIT(8'hF8) )  un1_data_out8_48_set_RNIGQ08 (.A(
        un1_data_out8_48_set_net_1), .B(un1_data_out8_183_rs_net_1), 
        .C(\mem_7_rs[2] ), .Y(\mem_7_[2]_net_1 ));
    CFG4 #( .INIT(16'hFFFE) )  \data_out_2_15_i_0_i[7]  (.A(
        \data_out_2_15_i_0_i_4[7]_net_1 ), .B(
        \data_out_2_15_i_0_i_5[7]_net_1 ), .C(
        \data_out_2_15_i_0_i_12[7]_net_1 ), .D(
        \data_out_2_15_i_0_i_11[7]_net_1 ), .Y(N_5));
    SLE un1_data_out8_148_rs (.D(VCC_net_1), .CLK(
        un1_data_out8_84_net_1), .EN(VCC_net_1), .ALn(
        un1_data_out8_148_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(VCC_net_1), .Q(un1_data_out8_148_rs_net_1));
    CFG3 #( .INIT(8'hF2) )  un1_data_out8_166 (.A(\mem_2_[6]_net_1 ), 
        .B(\mem_2__2_i_0_0_a2[0] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_166_i));
    SLE un1_data_out8_188_rs (.D(VCC_net_1), .CLK(
        un1_data_out8_71_net_1), .EN(VCC_net_1), .ALn(
        un1_data_out8_188_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(VCC_net_1), .Q(un1_data_out8_188_rs_net_1));
    SLE \mem_11_[2]  (.D(CoreAPB3_0_APBmslave4_PWDATA[2]), .CLK(
        FCCC_0_GL1), .EN(mem_11__1_sqmuxa), .ALn(un1_data_out8_226_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_11_rs[2] ));
    CFG4 #( .INIT(16'hEAC0) )  \data_out_2_15_i_i_4[5]  (.A(
        \mem_4_[5]_net_1 ), .B(\mem_2_[5]_net_1 ), .C(
        \mem_2__2_i_0_0_a2[0] ), .D(\mem_4__2_i_0_0_a2[0] ), .Y(
        \data_out_2_15_i_i_4[5]_net_1 ));
    CFG4 #( .INIT(16'hEAC0) )  \data_out_2_15_i_i_4[2]  (.A(
        \mem_4_[2]_net_1 ), .B(\mem_2_[2]_net_1 ), .C(
        \mem_2__2_i_0_0_a2[0] ), .D(\mem_4__2_i_0_0_a2[0] ), .Y(
        \data_out_2_15_i_i_4[2]_net_1 ));
    SLE un1_data_out8_195_rs (.D(VCC_net_1), .CLK(
        un1_data_out8_47_net_1), .EN(VCC_net_1), .ALn(
        un1_data_out8_195_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(VCC_net_1), .Q(un1_data_out8_195_rs_net_1));
    CFG3 #( .INIT(8'hF2) )  un1_data_out8_221 (.A(\mem_14_[5]_net_1 ), 
        .B(\mem_14__2_i_0_0_a2[2] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_221_i));
    CFG3 #( .INIT(8'h02) )  un1_data_out8_74 (.A(\mem_9_[2]_net_1 ), 
        .B(\mem_9__2_i_0_0_a2[0] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_74_net_1));
    SLE \mem_7_[2]  (.D(CoreAPB3_0_APBmslave4_PWDATA[2]), .CLK(
        FCCC_0_GL1), .EN(mem_7__1_sqmuxa), .ALn(un1_data_out8_183_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_7_rs[2] ));
    SLE un1_data_out8_169_rs (.D(VCC_net_1), .CLK(
        un1_data_out8_34_net_1), .EN(VCC_net_1), .ALn(
        un1_data_out8_169_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(VCC_net_1), .Q(un1_data_out8_169_rs_net_1));
    CFG2 #( .INIT(4'h8) )  mem_10__1_sqmuxa_0_a3_0_a3 (.A(
        mem_14__1_sqmuxa_0_a2_0_a3_0_a2_net_1), .B(
        \mem_10__2_i_0_0_a2[0] ), .Y(mem_10__1_sqmuxa));
    SLE un1_data_out8_51_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_3__1_sqmuxa), .ALn(un1_data_out8_51_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_data_out8_51_set_net_1));
    SLE un1_data_out8_155_rs (.D(VCC_net_1), .CLK(
        un1_data_out8_15_net_1), .EN(VCC_net_1), .ALn(
        un1_data_out8_155_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(VCC_net_1), .Q(un1_data_out8_155_rs_net_1));
    CFG1 #( .INIT(2'h1) )  un1_data_out8_16_set_RNO (.A(
        un1_data_out8_16_net_1), .Y(un1_data_out8_16_i));
    SLE un1_data_out8_110_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_13__1_sqmuxa), .ALn(un1_data_out8_110_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_data_out8_110_set_net_1));
    SLE \mem_2_[2]  (.D(CoreAPB3_0_APBmslave4_PWDATA[2]), .CLK(
        FCCC_0_GL1), .EN(mem_2__1_sqmuxa), .ALn(un1_data_out8_162_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_2_rs[2] ));
    CFG3 #( .INIT(8'h02) )  un1_data_out8_101 (.A(\mem_10_[4]_net_1 ), 
        .B(\mem_10__2_i_0_0_a2[0] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_101_net_1));
    CFG1 #( .INIT(2'h1) )  un1_data_out8_73_set_RNO (.A(
        un1_data_out8_73_net_1), .Y(un1_data_out8_73_i));
    SLE un1_data_out8_120_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_6__1_sqmuxa), .ALn(un1_data_out8_120_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_data_out8_120_set_net_1));
    CFG3 #( .INIT(8'h02) )  un1_data_out8_6 (.A(\mem_4_[3]_net_1 ), .B(
        \mem_4__2_i_0_0_a2[0] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_6_net_1));
    CFG3 #( .INIT(8'h02) )  un1_data_out8_38 (.A(\mem_6_[5]_net_1 ), 
        .B(\mem_6__2_i_0_0_a2[2] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_38_net_1));
    CFG3 #( .INIT(8'hF8) )  \mem_6__RNIB1OQ[4]  (.A(
        un1_data_out8_36_set_net_1), .B(un1_data_out8_171_rs_net_1), 
        .C(\mem_6_rs[4] ), .Y(\mem_6_[4]_net_1 ));
    CFG4 #( .INIT(16'hECA0) )  \data_out_2_15_i_i_5[5]  (.A(
        \mem_6_[5]_net_1 ), .B(\mem_1_[5]_net_1 ), .C(
        \mem_6__2_i_0_0_a2[2] ), .D(\mem_1__2_i_0_0_a2[0] ), .Y(
        \data_out_2_15_i_i_5[5]_net_1 ));
    CFG1 #( .INIT(2'h1) )  un1_data_out8_103_set_RNO (.A(
        un1_data_out8_103_net_1), .Y(un1_data_out8_103_i));
    SLE un1_data_out8_100_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_10__1_sqmuxa), .ALn(un1_data_out8_100_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_data_out8_100_set_net_1));
    CFG3 #( .INIT(8'hF2) )  un1_data_out8_251 (.A(\mem_15_[0]_net_1 ), 
        .B(\mem_15__2_i_0_0_a2[0] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_251_i));
    SLE \mem_5_[7]  (.D(CoreAPB3_0_APBmslave4_PWDATA[7]), .CLK(
        FCCC_0_GL1), .EN(mem_5__1_sqmuxa), .ALn(un1_data_out8_201_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_5_rs[7] ));
    CFG4 #( .INIT(16'h0080) )  \WRITE_GEN.mem_13__2_i_0_0_a2[0]  (.A(
        CoreAPB3_0_APBmslave4_PADDR[2]), .B(
        CoreAPB3_0_APBmslave4_PADDR[5]), .C(
        CoreAPB3_0_APBmslave4_PADDR[4]), .D(
        CoreAPB3_0_APBmslave4_PADDR[3]), .Y(\mem_13__2_i_0_0_a2[0] ));
    SLE \mem_4_[2]  (.D(CoreAPB3_0_APBmslave4_PWDATA[2]), .CLK(
        FCCC_0_GL1), .EN(mem_4__1_sqmuxa), .ALn(un1_data_out8_138_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_4_rs[2] ));
    CFG1 #( .INIT(2'h1) )  un1_data_out8_86_set_RNO (.A(
        un1_data_out8_86_net_1), .Y(un1_data_out8_86_i));
    CFG3 #( .INIT(8'hF8) )  un1_data_out8_153_rs_RNIS90M (.A(
        un1_data_out8_11_set_net_1), .B(un1_data_out8_153_rs_net_1), 
        .C(\mem_1_rs[1] ), .Y(\mem_1_[1]_net_1 ));
    SLE \mem_8_[6]  (.D(CoreAPB3_0_APBmslave4_PWDATA[6]), .CLK(
        FCCC_0_GL1), .EN(mem_8__1_sqmuxa), .ALn(un1_data_out8_186_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_8_rs[6] ));
    CFG3 #( .INIT(8'hF2) )  un1_data_out8_185 (.A(\mem_4_[7]_net_1 ), 
        .B(\mem_4__2_i_0_0_a2[0] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_185_i));
    CFG3 #( .INIT(8'hF2) )  un1_data_out8_212 (.A(\mem_13_[4]_net_1 ), 
        .B(\mem_13__2_i_0_0_a2[0] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_212_i));
    SLE \mem_5_[5]  (.D(CoreAPB3_0_APBmslave4_PWDATA[5]), .CLK(
        FCCC_0_GL1), .EN(mem_5__1_sqmuxa), .ALn(un1_data_out8_197_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_5_rs[5] ));
    CFG3 #( .INIT(8'hF8) )  \mem_6__RNI4FVN[0]  (.A(
        un1_data_out8_28_set_net_1), .B(un1_data_out8_203_rs_net_1), 
        .C(\mem_6_rs[0] ), .Y(\mem_6_[0]_net_1 ));
    CFG1 #( .INIT(2'h1) )  un1_data_out8_105_set_RNO (.A(
        un1_data_out8_105_net_1), .Y(un1_data_out8_105_i));
    CFG3 #( .INIT(8'h02) )  un1_data_out8_106 (.A(\mem_13_[2]_net_1 ), 
        .B(\mem_13__2_i_0_0_a2[0] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_106_net_1));
    CFG3 #( .INIT(8'hF2) )  un1_data_out8_197 (.A(\mem_5_[5]_net_1 ), 
        .B(\mem_5__2_i_0_0_a2[0] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_197_i));
    CFG3 #( .INIT(8'hF2) )  un1_data_out8_241 (.A(\mem_8_[3]_net_1 ), 
        .B(mem_8__2_i_0_0_a2[2]), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_241_i));
    CFG3 #( .INIT(8'hF8) )  un1_data_out8_149_rs_RNIFB6T (.A(
        un1_data_out8_85_set_net_1), .B(un1_data_out8_149_rs_net_1), 
        .C(\mem_0_rs[5] ), .Y(\mem_0_[5]_net_1 ));
    CFG4 #( .INIT(16'h0001) )  \WRITE_GEN.mem_0__2_i_0_0_a2[0]  (.A(
        CoreAPB3_0_APBmslave4_PADDR[2]), .B(
        CoreAPB3_0_APBmslave4_PADDR[5]), .C(
        CoreAPB3_0_APBmslave4_PADDR[4]), .D(
        CoreAPB3_0_APBmslave4_PADDR[3]), .Y(mem_0__2_i_0_0_a2[0]));
    CFG3 #( .INIT(8'h02) )  un1_data_out8_33 (.A(\mem_2_[4]_net_1 ), 
        .B(\mem_2__2_i_0_0_a2[0] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_33_net_1));
    CFG1 #( .INIT(2'h1) )  un1_data_out8_107_set_RNO (.A(
        un1_data_out8_107_net_1), .Y(un1_data_out8_107_i));
    SLE un1_data_out8_145_rs (.D(VCC_net_1), .CLK(
        un1_data_out8_82_net_1), .EN(VCC_net_1), .ALn(
        un1_data_out8_145_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(VCC_net_1), .Q(un1_data_out8_145_rs_net_1));
    CFG4 #( .INIT(16'hECA0) )  \data_out_2_15_i_0_i_5[3]  (.A(
        \mem_6_[3]_net_1 ), .B(\mem_1_[3]_net_1 ), .C(
        \mem_6__2_i_0_0_a2[2] ), .D(\mem_1__2_i_0_0_a2[0] ), .Y(
        \data_out_2_15_i_0_i_5[3]_net_1 ));
    CFG3 #( .INIT(8'hF2) )  un1_data_out8_227 (.A(\mem_7_[4]_net_1 ), 
        .B(\mem_7__2_i_0_0_a2[1] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_227_i));
    SLE un1_data_out8_201_rs (.D(VCC_net_1), .CLK(
        un1_data_out8_26_net_1), .EN(VCC_net_1), .ALn(
        un1_data_out8_201_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(VCC_net_1), .Q(un1_data_out8_201_rs_net_1));
    CFG3 #( .INIT(8'h02) )  un1_data_out8_66 (.A(\mem_8_[3]_net_1 ), 
        .B(mem_8__2_i_0_0_a2[2]), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_66_net_1));
    CFG3 #( .INIT(8'hF8) )  un1_data_out8_75_set_RNINJ8Q (.A(
        un1_data_out8_75_set_net_1), .B(un1_data_out8_196_rs_net_1), 
        .C(\mem_9_rs[3] ), .Y(\mem_9_[3]_net_1 ));
    SLE un1_data_out8_185_rs (.D(VCC_net_1), .CLK(
        un1_data_out8_10_net_1), .EN(VCC_net_1), .ALn(
        un1_data_out8_185_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(VCC_net_1), .Q(un1_data_out8_185_rs_net_1));
    CFG3 #( .INIT(8'h02) )  un1_data_out8_120 (.A(\mem_6_[6]_net_1 ), 
        .B(\mem_6__2_i_0_0_a2[2] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_120_net_1));
    CFG4 #( .INIT(16'hFFF8) )  \data_out_2_15_i_0_i_11[7]  (.A(
        \mem_5__2_i_0_0_a2[0] ), .B(\mem_5_[7]_net_1 ), .C(
        \data_out_2_15_i_0_i_7[7]_net_1 ), .D(N_381), .Y(
        \data_out_2_15_i_0_i_11[7]_net_1 ));
    SLE un1_data_out8_26_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_5__1_sqmuxa), .ALn(un1_data_out8_26_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_data_out8_26_set_net_1));
    SLE un1_data_out8_86_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_0__1_sqmuxa), .ALn(un1_data_out8_86_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_data_out8_86_set_net_1));
    SLE un1_data_out8_69_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_8__1_sqmuxa), .ALn(un1_data_out8_69_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_data_out8_69_set_net_1));
    CFG3 #( .INIT(8'hF8) )  \mem_15__RNI16E11[1]  (.A(
        un1_data_out8_58_set_net_1), .B(un1_data_out8_248_rs_net_1), 
        .C(\mem_15_rs[1] ), .Y(\mem_15_[1]_net_1 ));
    CFG3 #( .INIT(8'hF2) )  un1_data_out8_135 (.A(\mem_3_[7]_net_1 ), 
        .B(\mem_3__2_i_0_0_a2[0] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_135_i));
    SLE un1_data_out8_233_rs (.D(VCC_net_1), .CLK(
        un1_data_out8_1_net_1), .EN(VCC_net_1), .ALn(
        un1_data_out8_233_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(VCC_net_1), .Q(un1_data_out8_233_rs_net_1));
    SLE un1_data_out8_163_rs (.D(VCC_net_1), .CLK(
        un1_data_out8_31_net_1), .EN(VCC_net_1), .ALn(
        un1_data_out8_163_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(VCC_net_1), .Q(un1_data_out8_163_rs_net_1));
    CFG3 #( .INIT(8'h02) )  un1_data_out8_5 (.A(\mem_8_[1]_net_1 ), .B(
        mem_8__2_i_0_0_a2[2]), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_5_net_1));
    CFG2 #( .INIT(4'h8) )  mem_2__1_sqmuxa_0_a3_0_a3 (.A(
        mem_14__1_sqmuxa_0_a2_0_a3_0_a2_net_1), .B(
        \mem_2__2_i_0_0_a2[0] ), .Y(mem_2__1_sqmuxa));
    SLE un1_data_out8_248_rs (.D(VCC_net_1), .CLK(
        un1_data_out8_58_net_1), .EN(VCC_net_1), .ALn(
        un1_data_out8_248_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(VCC_net_1), .Q(un1_data_out8_248_rs_net_1));
    CFG4 #( .INIT(16'hECA0) )  \data_out_2_15_i_0_i_7[1]  (.A(
        \mem_8_[1]_net_1 ), .B(\mem_0_[1]_net_1 ), .C(
        mem_8__2_i_0_0_a2[2]), .D(mem_0__2_i_0_0_a2[0]), .Y(
        \data_out_2_15_i_0_i_7[1]_net_1 ));
    CFG3 #( .INIT(8'hF2) )  un1_data_out8_150 (.A(\mem_0_[6]_net_1 ), 
        .B(mem_0__2_i_0_0_a2[0]), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_150_i));
    SLE un1_data_out8_112_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_14__1_sqmuxa), .ALn(un1_data_out8_112_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_data_out8_112_set_net_1));
    SLE \mem_7_[1]  (.D(CoreAPB3_0_APBmslave4_PWDATA[1]), .CLK(
        FCCC_0_GL1), .EN(mem_7__1_sqmuxa), .ALn(un1_data_out8_181_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_7_rs[1] ));
    SLE \mem_10_[0]  (.D(CoreAPB3_0_APBmslave4_PWDATA[0]), .CLK(
        FCCC_0_GL1), .EN(mem_10__1_sqmuxa), .ALn(un1_data_out8_206_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_10_rs[0] ));
    CFG3 #( .INIT(8'hF2) )  un1_data_out8_223 (.A(\mem_14_[7]_net_1 ), 
        .B(\mem_14__2_i_0_0_a2[2] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_223_i));
    SLE un1_data_out8_176_rs (.D(VCC_net_1), .CLK(
        un1_data_out8_102_net_1), .EN(VCC_net_1), .ALn(
        un1_data_out8_176_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(VCC_net_1), .Q(un1_data_out8_176_rs_net_1));
    SLE \mem_13_[7]  (.D(CoreAPB3_0_APBmslave4_PWDATA[7]), .CLK(
        FCCC_0_GL1), .EN(mem_13__1_sqmuxa), .ALn(un1_data_out8_215_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_13_rs[7] ));
    CFG1 #( .INIT(2'h1) )  un1_data_out8_60_set_RNO (.A(
        un1_data_out8_60_net_1), .Y(un1_data_out8_60_i));
    SLE un1_data_out8_61_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_15__1_sqmuxa), .ALn(un1_data_out8_61_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_data_out8_61_set_net_1));
    SLE un1_data_out8_223_rs (.D(VCC_net_1), .CLK(
        un1_data_out8_119_net_1), .EN(VCC_net_1), .ALn(
        un1_data_out8_223_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(VCC_net_1), .Q(un1_data_out8_223_rs_net_1));
    SLE \mem_14_[5]  (.D(CoreAPB3_0_APBmslave4_PWDATA[5]), .CLK(
        FCCC_0_GL1), .EN(mem_14__1_sqmuxa), .ALn(un1_data_out8_221_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_14_rs[5] ));
    SLE un1_data_out8_76_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_9__1_sqmuxa), .ALn(un1_data_out8_76_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_data_out8_76_set_net_1));
    SLE un1_data_out8_122_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_6__1_sqmuxa), .ALn(un1_data_out8_122_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_data_out8_122_set_net_1));
    SLE \mem_2_[1]  (.D(CoreAPB3_0_APBmslave4_PWDATA[1]), .CLK(
        FCCC_0_GL1), .EN(mem_2__1_sqmuxa), .ALn(un1_data_out8_161_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_2_rs[1] ));
    CFG3 #( .INIT(8'h02) )  un1_data_out8_37 (.A(\mem_2_[6]_net_1 ), 
        .B(\mem_2__2_i_0_0_a2[0] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_37_net_1));
    CFG3 #( .INIT(8'hF2) )  un1_data_out8_247 (.A(\mem_12_[7]_net_1 ), 
        .B(\mem_12__2_i_0_0_a2[0] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_247_i));
    SLE un1_data_out8_102_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_10__1_sqmuxa), .ALn(un1_data_out8_102_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_data_out8_102_set_net_1));
    CFG4 #( .INIT(16'h1000) )  \WRITE_GEN.mem_6__2_i_0_0_a2[2]  (.A(
        CoreAPB3_0_APBmslave4_PADDR[2]), .B(
        CoreAPB3_0_APBmslave4_PADDR[5]), .C(
        CoreAPB3_0_APBmslave4_PADDR[4]), .D(
        CoreAPB3_0_APBmslave4_PADDR[3]), .Y(\mem_6__2_i_0_0_a2[2] ));
    CFG1 #( .INIT(2'h1) )  un1_data_out8_68_set_RNO (.A(
        un1_data_out8_68_net_1), .Y(un1_data_out8_68_i));
    SLE un1_data_out8_53_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_3__1_sqmuxa), .ALn(un1_data_out8_53_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_data_out8_53_set_net_1));
    SLE \mem_3_[4]  (.D(CoreAPB3_0_APBmslave4_PWDATA[4]), .CLK(
        FCCC_0_GL1), .EN(mem_3__1_sqmuxa), .ALn(un1_data_out8_132_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_3_rs[4] ));
    CFG3 #( .INIT(8'hF2) )  un1_data_out8_140 (.A(\mem_4_[4]_net_1 ), 
        .B(\mem_4__2_i_0_0_a2[0] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_140_i));
    CFG1 #( .INIT(2'h1) )  un1_data_out8_108_set_RNO (.A(
        un1_data_out8_108_net_1), .Y(un1_data_out8_108_i));
    SLE un1_data_out8_254_rs (.D(VCC_net_1), .CLK(
        un1_data_out8_60_net_1), .EN(VCC_net_1), .ALn(
        un1_data_out8_254_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(VCC_net_1), .Q(un1_data_out8_254_rs_net_1));
    CFG3 #( .INIT(8'hF2) )  un1_data_out8_238 (.A(\mem_12_[0]_net_1 ), 
        .B(\mem_12__2_i_0_0_a2[0] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_238_i));
    SLE un1_data_out8_168_rs (.D(VCC_net_1), .CLK(
        un1_data_out8_98_net_1), .EN(VCC_net_1), .ALn(
        un1_data_out8_168_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(VCC_net_1), .Q(un1_data_out8_168_rs_net_1));
    SLE \mem_4_[1]  (.D(CoreAPB3_0_APBmslave4_PWDATA[1]), .CLK(
        FCCC_0_GL1), .EN(mem_4__1_sqmuxa), .ALn(un1_data_out8_137_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_4_rs[1] ));
    CFG3 #( .INIT(8'h02) )  un1_data_out8_60 (.A(\mem_15_[7]_net_1 ), 
        .B(\mem_15__2_i_0_0_a2[0] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_60_net_1));
    CFG4 #( .INIT(16'hECA0) )  \data_out_2_15_i_i_1[4]  (.A(
        \mem_14_[4]_net_1 ), .B(\mem_9_[4]_net_1 ), .C(
        \mem_14__2_i_0_0_a2[2] ), .D(\mem_9__2_i_0_0_a2[0] ), .Y(
        \data_out_2_15_i_i_1[4]_net_1 ));
    CFG3 #( .INIT(8'h02) )  un1_data_out8_56 (.A(\mem_15_[3]_net_1 ), 
        .B(\mem_15__2_i_0_0_a2[0] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_56_net_1));
    CFG3 #( .INIT(8'hF2) )  un1_data_out8_253 (.A(\mem_15_[6]_net_1 ), 
        .B(\mem_15__2_i_0_0_a2[0] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_253_i));
    CFG3 #( .INIT(8'hF2) )  un1_data_out8_175 (.A(\mem_6_[6]_net_1 ), 
        .B(\mem_6__2_i_0_0_a2[2] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_175_i));
    CFG3 #( .INIT(8'h02) )  un1_data_out8_123 (.A(\mem_3_[1]_net_1 ), 
        .B(\mem_3__2_i_0_0_a2[0] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_123_net_1));
    CFG1 #( .INIT(2'h1) )  un1_data_out8_9_set_RNO (.A(
        un1_data_out8_9_net_1), .Y(un1_data_out8_9_i));
    SLE \mem_11_[7]  (.D(CoreAPB3_0_APBmslave4_PWDATA[7]), .CLK(
        FCCC_0_GL1), .EN(mem_11__1_sqmuxa), .ALn(un1_data_out8_236_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_11_rs[7] ));
    SLE \mem_14_[1]  (.D(CoreAPB3_0_APBmslave4_PWDATA[1]), .CLK(
        FCCC_0_GL1), .EN(mem_14__1_sqmuxa), .ALn(un1_data_out8_217_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_14_rs[1] ));
    CFG3 #( .INIT(8'hF2) )  un1_data_out8_189 (.A(\mem_5_[1]_net_1 ), 
        .B(\mem_5__2_i_0_0_a2[0] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_189_i));
    CFG3 #( .INIT(8'hF8) )  un1_data_out8_68_set_RNIGNVU (.A(
        un1_data_out8_68_set_net_1), .B(un1_data_out8_142_rs_net_1), 
        .C(\mem_8_rs[4] ), .Y(\mem_8_[4]_net_1 ));
    CFG1 #( .INIT(2'h1) )  un1_data_out8_24_set_RNO (.A(
        un1_data_out8_24_net_1), .Y(un1_data_out8_24_i));
    SLE un1_data_out8_132_rs (.D(VCC_net_1), .CLK(
        un1_data_out8_49_net_1), .EN(VCC_net_1), .ALn(
        un1_data_out8_132_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(VCC_net_1), .Q(un1_data_out8_132_rs_net_1));
    SLE un1_data_out8_179_rs (.D(VCC_net_1), .CLK(
        un1_data_out8_124_net_1), .EN(VCC_net_1), .ALn(
        un1_data_out8_179_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(VCC_net_1), .Q(un1_data_out8_179_rs_net_1));
    CFG4 #( .INIT(16'hECA0) )  \data_out_2_15_i_0_i_1[1]  (.A(
        \mem_14_[1]_net_1 ), .B(\mem_9_[1]_net_1 ), .C(
        \mem_14__2_i_0_0_a2[2] ), .D(\mem_9__2_i_0_0_a2[0] ), .Y(
        \data_out_2_15_i_0_i_1[1]_net_1 ));
    CFG4 #( .INIT(16'hEAC0) )  \data_out_2_15_i_0_i_0[7]  (.A(
        \mem_10_[7]_net_1 ), .B(\mem_12_[7]_net_1 ), .C(
        \mem_12__2_i_0_0_a2[0] ), .D(\mem_10__2_i_0_0_a2[0] ), .Y(
        \data_out_2_15_i_0_i_0[7]_net_1 ));
    SLE un1_data_out8_54_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_7__1_sqmuxa), .ALn(un1_data_out8_54_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_data_out8_54_set_net_1));
    CFG3 #( .INIT(8'hF8) )  un1_data_out8_200_rs_RNIDCL01 (.A(
        un1_data_out8_77_set_net_1), .B(un1_data_out8_200_rs_net_1), 
        .C(\mem_9_rs[5] ), .Y(\mem_9_[5]_net_1 ));
    CFG1 #( .INIT(2'h1) )  un1_data_out8_30_set_RNO (.A(
        un1_data_out8_30_net_1), .Y(un1_data_out8_30_i));
    CFG1 #( .INIT(2'h1) )  un1_data_out8_13_set_RNO (.A(
        un1_data_out8_13_net_1), .Y(un1_data_out8_13_i));
    CFG3 #( .INIT(8'hF8) )  un1_data_out8_26_set_RNI647P (.A(
        un1_data_out8_26_set_net_1), .B(un1_data_out8_201_rs_net_1), 
        .C(\mem_5_rs[7] ), .Y(\mem_5_[7]_net_1 ));
    CFG4 #( .INIT(16'hEAC0) )  \data_out_2_15_i_i_3[4]  (.A(
        \mem_15_[4]_net_1 ), .B(\mem_7_[4]_net_1 ), .C(
        \mem_7__2_i_0_0_a2[1] ), .D(\mem_15__2_i_0_0_a2[0] ), .Y(
        \data_out_2_15_i_i_3[4]_net_1 ));
    CFG3 #( .INIT(8'hF2) )  un1_data_out8_243 (.A(\mem_12_[3]_net_1 ), 
        .B(\mem_12__2_i_0_0_a2[0] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_243_i));
    CFG1 #( .INIT(2'h1) )  un1_data_out8_1_set_RNO (.A(
        un1_data_out8_1_net_1), .Y(un1_data_out8_1_i));
    CFG1 #( .INIT(2'h1) )  un1_data_out8_50_set_RNO (.A(
        un1_data_out8_50_net_1), .Y(un1_data_out8_50_i));
    CFG3 #( .INIT(8'hF8) )  un1_data_out8_209_rs_RNI55JJ (.A(
        un1_data_out8_105_set_net_1), .B(un1_data_out8_209_rs_net_1), 
        .C(\mem_13_rs[1] ), .Y(\mem_13_[1]_net_1 ));
    SLE un1_data_out8_202_rs (.D(VCC_net_1), .CLK(
        un1_data_out8_78_net_1), .EN(VCC_net_1), .ALn(
        un1_data_out8_202_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(VCC_net_1), .Q(un1_data_out8_202_rs_net_1));
    SLE un1_data_out8_237_rs (.D(VCC_net_1), .CLK(
        un1_data_out8_5_net_1), .EN(VCC_net_1), .ALn(
        un1_data_out8_237_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(VCC_net_1), .Q(un1_data_out8_237_rs_net_1));
    CFG3 #( .INIT(8'hF8) )  \mem_6__RNI0RUI[1]  (.A(
        un1_data_out8_30_set_net_1), .B(un1_data_out8_205_rs_net_1), 
        .C(\mem_6_rs[1] ), .Y(\mem_6_[1]_net_1 ));
    SLE un1_data_out8_215_rs (.D(VCC_net_1), .CLK(
        un1_data_out8_111_net_1), .EN(VCC_net_1), .ALn(
        un1_data_out8_215_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(VCC_net_1), .Q(un1_data_out8_215_rs_net_1));
    CFG3 #( .INIT(8'hF2) )  un1_data_out8_153 (.A(\mem_1_[1]_net_1 ), 
        .B(\mem_1__2_i_0_0_a2[0] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_153_i));
    CFG1 #( .INIT(2'h1) )  un1_data_out8_38_set_RNO (.A(
        un1_data_out8_38_net_1), .Y(un1_data_out8_38_i));
    SLE \mem_6_[3]  (.D(CoreAPB3_0_APBmslave4_PWDATA[3]), .CLK(
        FCCC_0_GL1), .EN(mem_6__1_sqmuxa), .ALn(un1_data_out8_169_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_6_rs[3] ));
    CFG3 #( .INIT(8'hF8) )  \mem_6__RNIRB1M[6]  (.A(
        un1_data_out8_120_set_net_1), .B(un1_data_out8_175_rs_net_1), 
        .C(\mem_6_rs[6] ), .Y(\mem_6_[6]_net_1 ));
    CFG1 #( .INIT(2'h1) )  un1_data_out8_58_set_RNO (.A(
        un1_data_out8_58_net_1), .Y(un1_data_out8_58_i));
    CFG1 #( .INIT(2'h1) )  un1_data_out8_40_set_RNO (.A(
        un1_data_out8_40_net_1), .Y(un1_data_out8_40_i));
    CFG3 #( .INIT(8'hF8) )  \mem_6__RNI5AHT[2]  (.A(
        un1_data_out8_32_set_net_1), .B(un1_data_out8_207_rs_net_1), 
        .C(\mem_6_rs[2] ), .Y(\mem_6_[2]_net_1 ));
    CFG1 #( .INIT(2'h1) )  un1_data_out8_83_set_RNO (.A(
        un1_data_out8_83_net_1), .Y(un1_data_out8_83_i));
    CFG3 #( .INIT(8'hF2) )  un1_data_out8_139 (.A(\mem_4_[3]_net_1 ), 
        .B(\mem_4__2_i_0_0_a2[0] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_139_i));
    CFG1 #( .INIT(2'h1) )  un1_data_out8_122_set_RNO (.A(
        un1_data_out8_122_net_1), .Y(un1_data_out8_122_i));
    SLE un1_data_out8_227_rs (.D(VCC_net_1), .CLK(
        un1_data_out8_52_net_1), .EN(VCC_net_1), .ALn(
        un1_data_out8_227_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(VCC_net_1), .Q(un1_data_out8_227_rs_net_1));
    SLE un1_data_out8_244_rs (.D(VCC_net_1), .CLK(
        un1_data_out8_20_net_1), .EN(VCC_net_1), .ALn(
        un1_data_out8_244_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(VCC_net_1), .Q(un1_data_out8_244_rs_net_1));
    CFG2 #( .INIT(4'h8) )  mem_9__1_sqmuxa_0_a3_0_a3 (.A(
        mem_14__1_sqmuxa_0_a2_0_a3_0_a2_net_1), .B(
        \mem_9__2_i_0_0_a2[0] ), .Y(mem_9__1_sqmuxa));
    CFG3 #( .INIT(8'hF2) )  un1_data_out8_143 (.A(\mem_4_[6]_net_1 ), 
        .B(\mem_4__2_i_0_0_a2[0] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_143_i));
    CFG1 #( .INIT(2'h1) )  un1_data_out8_48_set_RNO (.A(
        un1_data_out8_48_net_1), .Y(un1_data_out8_48_i));
    CFG3 #( .INIT(8'hF2) )  un1_data_out8_215 (.A(\mem_13_[7]_net_1 ), 
        .B(\mem_13__2_i_0_0_a2[0] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_215_i));
    SLE \mem_3_[0]  (.D(CoreAPB3_0_APBmslave4_PWDATA[0]), .CLK(
        FCCC_0_GL1), .EN(mem_3__1_sqmuxa), .ALn(un1_data_out8_128_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_3_rs[0] ));
    CFG1 #( .INIT(2'h1) )  un1_data_out8_27_set_RNO (.A(
        un1_data_out8_27_net_1), .Y(un1_data_out8_27_i));
    CFG3 #( .INIT(8'hF8) )  \mem_6__RNIFCUM[3]  (.A(
        un1_data_out8_34_set_net_1), .B(un1_data_out8_169_rs_net_1), 
        .C(\mem_6_rs[3] ), .Y(\mem_6_[3]_net_1 ));
    SLE \mem_0_[3]  (.D(CoreAPB3_0_APBmslave4_PWDATA[3]), .CLK(
        FCCC_0_GL1), .EN(mem_0__1_sqmuxa), .ALn(un1_data_out8_146_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_0_rs[3] ));
    SLE un1_data_out8_119_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_14__1_sqmuxa), .ALn(un1_data_out8_119_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_data_out8_119_set_net_1));
    CFG3 #( .INIT(8'h02) )  un1_data_out8_50 (.A(\mem_7_[3]_net_1 ), 
        .B(\mem_7__2_i_0_0_a2[1] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_50_net_1));
    CFG3 #( .INIT(8'hF2) )  un1_data_out8_229 (.A(\mem_7_[5]_net_1 ), 
        .B(\mem_7__2_i_0_0_a2[1] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_229_i));
    CFG3 #( .INIT(8'hF8) )  un1_data_out8_249_rs_RNI4ENM (.A(
        un1_data_out8_59_set_net_1), .B(un1_data_out8_249_rs_net_1), 
        .C(\mem_15_rs[2] ), .Y(\mem_15_[2]_net_1 ));
    CFG3 #( .INIT(8'h02) )  un1_data_out8_81 (.A(\mem_0_[1]_net_1 ), 
        .B(mem_0__2_i_0_0_a2[0]), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_81_net_1));
    CFG4 #( .INIT(16'hEAC0) )  \data_out_2_15_i_i_2[4]  (.A(
        \mem_13_[4]_net_1 ), .B(\mem_11_[4]_net_1 ), .C(
        \mem_11__2_i_0_0_a2[2] ), .D(\mem_13__2_i_0_0_a2[0] ), .Y(
        \data_out_2_15_i_i_2[4]_net_1 ));
    CFG3 #( .INIT(8'h02) )  un1_data_out8_22 (.A(\mem_12_[6]_net_1 ), 
        .B(\mem_12__2_i_0_0_a2[0] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_22_net_1));
    CFG3 #( .INIT(8'hF2) )  un1_data_out8_188 (.A(\mem_8_[7]_net_1 ), 
        .B(mem_8__2_i_0_0_a2[2]), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_188_i));
    CFG3 #( .INIT(8'h02) )  un1_data_out8_114 (.A(\mem_14_[2]_net_1 ), 
        .B(\mem_14__2_i_0_0_a2[2] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_114_net_1));
    CFG3 #( .INIT(8'h02) )  un1_data_out8_18 (.A(\mem_12_[2]_net_1 ), 
        .B(\mem_12__2_i_0_0_a2[0] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_18_net_1));
    CFG3 #( .INIT(8'hF8) )  un1_data_out8_76_set_RNIRUK01 (.A(
        un1_data_out8_76_set_net_1), .B(un1_data_out8_198_rs_net_1), 
        .C(\mem_9_rs[4] ), .Y(\mem_9_[4]_net_1 ));
    SLE un1_data_out8_165_rs (.D(VCC_net_1), .CLK(
        un1_data_out8_35_net_1), .EN(VCC_net_1), .ALn(
        un1_data_out8_165_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(VCC_net_1), .Q(un1_data_out8_165_rs_net_1));
    SLE un1_data_out8_109_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_13__1_sqmuxa), .ALn(un1_data_out8_109_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_data_out8_109_set_net_1));
    CFG3 #( .INIT(8'hF8) )  un1_data_out8_190_rs_RNIBI3N (.A(
        un1_data_out8_72_set_net_1), .B(un1_data_out8_190_rs_net_1), 
        .C(\mem_9_rs[0] ), .Y(\mem_9_[0]_net_1 ));
    CFG4 #( .INIT(16'hEAC0) )  \data_out_2_15_i_i_2[6]  (.A(
        \mem_13_[6]_net_1 ), .B(\mem_11_[6]_net_1 ), .C(
        \mem_11__2_i_0_0_a2[2] ), .D(\mem_13__2_i_0_0_a2[0] ), .Y(
        \data_out_2_15_i_i_2[6]_net_1 ));
    CFG1 #( .INIT(2'h1) )  un1_data_out8_94_set_RNO (.A(
        un1_data_out8_94_net_1), .Y(un1_data_out8_94_i));
    SLE \mem_15_[4]  (.D(CoreAPB3_0_APBmslave4_PWDATA[4]), .CLK(
        FCCC_0_GL1), .EN(mem_15__1_sqmuxa), .ALn(un1_data_out8_255_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_15_rs[4] ));
    CFG3 #( .INIT(8'hF8) )  un1_data_out8_146_rs_RNI8OGH (.A(
        un1_data_out8_83_set_net_1), .B(un1_data_out8_146_rs_net_1), 
        .C(\mem_0_rs[3] ), .Y(\mem_0_[3]_net_1 ));
    SLE un1_data_out8_63_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_15__1_sqmuxa), .ALn(un1_data_out8_63_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_data_out8_63_set_net_1));
    CFG3 #( .INIT(8'h02) )  un1_data_out8_42 (.A(\mem_1_[5]_net_1 ), 
        .B(\mem_1__2_i_0_0_a2[0] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_42_net_1));
    SLE un1_data_out8_173_rs (.D(VCC_net_1), .CLK(
        un1_data_out8_38_net_1), .EN(VCC_net_1), .ALn(
        un1_data_out8_173_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(VCC_net_1), .Q(un1_data_out8_173_rs_net_1));
    CFG3 #( .INIT(8'hF8) )  un1_data_out8_224_rs_RNIRK1N (.A(
        un1_data_out8_89_set_net_1), .B(un1_data_out8_224_rs_net_1), 
        .C(\mem_11_rs[1] ), .Y(\mem_11_[1]_net_1 ));
    CFG1 #( .INIT(2'h1) )  un1_data_out8_62_set_RNO (.A(
        un1_data_out8_62_net_1), .Y(un1_data_out8_62_i));
    CFG3 #( .INIT(8'hF2) )  un1_data_out8_200 (.A(\mem_9_[5]_net_1 ), 
        .B(\mem_9__2_i_0_0_a2[0] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_200_i));
    CFG3 #( .INIT(8'hF2) )  un1_data_out8_179 (.A(\mem_7_[0]_net_1 ), 
        .B(\mem_7__2_i_0_0_a2[1] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_179_i));
    CFG1 #( .INIT(2'h1) )  un1_data_out8_75_set_RNO (.A(
        un1_data_out8_75_net_1), .Y(un1_data_out8_75_i));
    SLE \mem_12_[3]  (.D(CoreAPB3_0_APBmslave4_PWDATA[3]), .CLK(
        FCCC_0_GL1), .EN(mem_12__1_sqmuxa), .ALn(un1_data_out8_243_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_12_rs[3] ));
    CFG2 #( .INIT(4'h8) )  mem_11__1_sqmuxa_0_a2_0_a3_0_a3 (.A(
        mem_14__1_sqmuxa_0_a2_0_a3_0_a2_net_1), .B(
        \mem_11__2_i_0_0_a2[2] ), .Y(mem_11__1_sqmuxa));
    SLE un1_data_out8_3_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_7__1_sqmuxa), .ALn(un1_data_out8_3_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_data_out8_3_set_net_1));
    CFG3 #( .INIT(8'h02) )  un1_data_out8_71 (.A(\mem_8_[7]_net_1 ), 
        .B(mem_8__2_i_0_0_a2[2]), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_71_net_1));
    SLE un1_data_out8_6_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_4__1_sqmuxa), .ALn(un1_data_out8_6_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_data_out8_6_set_net_1));
    CFG3 #( .INIT(8'h02) )  un1_data_out8_25 (.A(\mem_2_[0]_net_1 ), 
        .B(\mem_2__2_i_0_0_a2[0] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_25_net_1));
    SLE un1_data_out8_58_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_15__1_sqmuxa), .ALn(un1_data_out8_58_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_data_out8_58_set_net_1));
    CFG3 #( .INIT(8'hF8) )  \mem_2__RNIVS5M[0]  (.A(
        un1_data_out8_25_set_net_1), .B(un1_data_out8_160_rs_net_1), 
        .C(\mem_2_rs[0] ), .Y(\mem_2_[0]_net_1 ));
    CFG1 #( .INIT(2'h1) )  un1_data_out8_111_set_RNO (.A(
        un1_data_out8_111_net_1), .Y(un1_data_out8_111_i));
    CFG3 #( .INIT(8'hF8) )  un1_data_out8_127_set_RNIKSKH (.A(
        un1_data_out8_127_set_net_1), .B(un1_data_out8_131_rs_net_1), 
        .C(\mem_3_rs[3] ), .Y(\mem_3_[3]_net_1 ));
    CFG3 #( .INIT(8'hF2) )  un1_data_out8_138 (.A(\mem_4_[2]_net_1 ), 
        .B(\mem_4__2_i_0_0_a2[0] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_138_i));
    CFG3 #( .INIT(8'h02) )  un1_data_out8_13 (.A(\mem_1_[2]_net_1 ), 
        .B(\mem_1__2_i_0_0_a2[0] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_13_net_1));
    SLE un1_data_out8_47_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_5__1_sqmuxa), .ALn(un1_data_out8_47_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_data_out8_47_set_net_1));
    SLE \mem_7_[6]  (.D(CoreAPB3_0_APBmslave4_PWDATA[6]), .CLK(
        FCCC_0_GL1), .EN(mem_7__1_sqmuxa), .ALn(un1_data_out8_231_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_7_rs[6] ));
    SLE un1_data_out8_90_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_11__1_sqmuxa), .ALn(un1_data_out8_90_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_data_out8_90_set_net_1));
    SLE un1_data_out8_29_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_2__1_sqmuxa), .ALn(un1_data_out8_29_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_data_out8_29_set_net_1));
    SLE un1_data_out8_89_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_11__1_sqmuxa), .ALn(un1_data_out8_89_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_data_out8_89_set_net_1));
    SLE un1_data_out8_64_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_8__1_sqmuxa), .ALn(un1_data_out8_64_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_data_out8_64_set_net_1));
    CFG2 #( .INIT(4'h8) )  \data_out_2_15_i_i_a3_8[5]  (.A(
        \mem_3__2_i_0_0_a2[0] ), .B(\mem_3_[5]_net_1 ), .Y(
        \data_out_2_15_i_i_a3_8[5]_net_1 ));
    CFG3 #( .INIT(8'hF2) )  un1_data_out8_249 (.A(\mem_15_[2]_net_1 ), 
        .B(\mem_15__2_i_0_0_a2[0] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_249_i));
    SLE \mem_15_[6]  (.D(CoreAPB3_0_APBmslave4_PWDATA[6]), .CLK(
        FCCC_0_GL1), .EN(mem_15__1_sqmuxa), .ALn(un1_data_out8_253_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_15_rs[6] ));
    CFG3 #( .INIT(8'h02) )  un1_data_out8_45 (.A(\mem_5_[5]_net_1 ), 
        .B(\mem_5__2_i_0_0_a2[0] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_45_net_1));
    CFG1 #( .INIT(2'h1) )  un1_data_out8_71_set_RNO (.A(
        un1_data_out8_71_net_1), .Y(un1_data_out8_71_i));
    CFG3 #( .INIT(8'hF8) )  un1_data_out8_215_rs_RNI5OUS (.A(
        un1_data_out8_111_set_net_1), .B(un1_data_out8_215_rs_net_1), 
        .C(\mem_13_rs[7] ), .Y(\mem_13_[7]_net_1 ));
    SLE \mem_2_[6]  (.D(CoreAPB3_0_APBmslave4_PWDATA[6]), .CLK(
        FCCC_0_GL1), .EN(mem_2__1_sqmuxa), .ALn(un1_data_out8_166_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_2_rs[6] ));
    CFG3 #( .INIT(8'h02) )  un1_data_out8_24 (.A(\mem_5_[6]_net_1 ), 
        .B(\mem_5__2_i_0_0_a2[0] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_24_net_1));
    CFG1 #( .INIT(2'h1) )  un1_data_out8_26_set_RNO (.A(
        un1_data_out8_26_net_1), .Y(un1_data_out8_26_i));
    SLE \mem_1_[3]  (.D(CoreAPB3_0_APBmslave4_PWDATA[3]), .CLK(
        FCCC_0_GL1), .EN(mem_1__1_sqmuxa), .ALn(un1_data_out8_155_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_1_rs[3] ));
    SLE \mem_9_[3]  (.D(CoreAPB3_0_APBmslave4_PWDATA[3]), .CLK(
        FCCC_0_GL1), .EN(mem_9__1_sqmuxa), .ALn(un1_data_out8_196_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_9_rs[3] ));
    CFG4 #( .INIT(16'hFFFE) )  \data_out_2_15_i_0_i_12[1]  (.A(
        \data_out_2_15_i_0_i_2[1]_net_1 ), .B(
        \data_out_2_15_i_0_i_1[1]_net_1 ), .C(
        \data_out_2_15_i_0_i_3[1]_net_1 ), .D(
        \data_out_2_15_i_0_i_0[1]_net_1 ), .Y(
        \data_out_2_15_i_0_i_12[1]_net_1 ));
    CFG1 #( .INIT(2'h1) )  un1_data_out8_97_set_RNO (.A(
        un1_data_out8_97_net_1), .Y(un1_data_out8_97_i));
    CFG3 #( .INIT(8'hF8) )  \mem_7__RNIHHAP[5]  (.A(
        un1_data_out8_54_set_net_1), .B(un1_data_out8_229_rs_net_1), 
        .C(\mem_7_rs[5] ), .Y(\mem_7_[5]_net_1 ));
    CFG3 #( .INIT(8'hF8) )  un1_data_out8_138_rs_RNIL15L (.A(
        un1_data_out8_4_set_net_1), .B(un1_data_out8_138_rs_net_1), .C(
        \mem_4_rs[2] ), .Y(\mem_4_[2]_net_1 ));
    CFG1 #( .INIT(2'h1) )  un1_data_out8_32_set_RNO (.A(
        un1_data_out8_32_net_1), .Y(un1_data_out8_32_i));
    SLE un1_data_out8_178_rs (.D(VCC_net_1), .CLK(
        un1_data_out8_103_net_1), .EN(VCC_net_1), .ALn(
        un1_data_out8_178_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(VCC_net_1), .Q(un1_data_out8_178_rs_net_1));
    CFG3 #( .INIT(8'h80) )  mem_14__1_sqmuxa_0_a2_0_a3_0_a2 (.A(
        CoreAPB3_0_APBmslave4_PENABLE), .B(PRDATA_0_iv_0_0_a2_1[3]), 
        .C(CoreAPB3_0_APBmslave4_PWRITE), .Y(
        mem_14__1_sqmuxa_0_a2_0_a3_0_a2_net_1));
    SLE \mem_4_[6]  (.D(CoreAPB3_0_APBmslave4_PWDATA[6]), .CLK(
        FCCC_0_GL1), .EN(mem_4__1_sqmuxa), .ALn(un1_data_out8_143_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_4_rs[6] ));
    SLE un1_data_out8_253_rs (.D(VCC_net_1), .CLK(
        un1_data_out8_63_net_1), .EN(VCC_net_1), .ALn(
        un1_data_out8_253_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(VCC_net_1), .Q(un1_data_out8_253_rs_net_1));
    CFG1 #( .INIT(2'h1) )  un1_data_out8_116_set_RNO (.A(
        un1_data_out8_116_net_1), .Y(un1_data_out8_116_i));
    CFG3 #( .INIT(8'h02) )  un1_data_out8_44 (.A(\mem_1_[6]_net_1 ), 
        .B(\mem_1__2_i_0_0_a2[0] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_44_net_1));
    CFG1 #( .INIT(2'h1) )  un1_data_out8_52_set_RNO (.A(
        un1_data_out8_52_net_1), .Y(un1_data_out8_52_i));
    SLE un1_data_out8_21_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_12__1_sqmuxa), .ALn(un1_data_out8_21_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_data_out8_21_set_net_1));
    SLE un1_data_out8_81_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_0__1_sqmuxa), .ALn(un1_data_out8_81_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_data_out8_81_set_net_1));
    SLE un1_data_out8_79_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_9__1_sqmuxa), .ALn(un1_data_out8_79_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_data_out8_79_set_net_1));
    CFG3 #( .INIT(8'hF2) )  un1_data_out8_211 (.A(\mem_13_[3]_net_1 ), 
        .B(\mem_13__2_i_0_0_a2[0] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_211_i));
    CFG3 #( .INIT(8'h02) )  un1_data_out8_39 (.A(\mem_2_[7]_net_1 ), 
        .B(\mem_2__2_i_0_0_a2[0] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_39_net_1));
    SLE \data_out[7]  (.D(N_5), .CLK(FCCC_0_GL1), .EN(rd_enable), .ALn(
        MSS_RESET_N_M2F_c), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(
        CoreAPB3_0_APBmslave5_PRDATA[7]));
    CFG3 #( .INIT(8'hF8) )  un1_data_out8_56_set_RNIQBFK (.A(
        un1_data_out8_56_set_net_1), .B(un1_data_out8_250_rs_net_1), 
        .C(\mem_15_rs[3] ), .Y(\mem_15_[3]_net_1 ));
    CFG1 #( .INIT(2'h1) )  un1_data_out8_42_set_RNO (.A(
        un1_data_out8_42_net_1), .Y(un1_data_out8_42_i));
    CFG3 #( .INIT(8'hF2) )  un1_data_out8_178 (.A(\mem_10_[6]_net_1 ), 
        .B(\mem_10__2_i_0_0_a2[0] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_178_i));
    CFG3 #( .INIT(8'h02) )  un1_data_out8_17 (.A(\mem_12_[1]_net_1 ), 
        .B(\mem_12__2_i_0_0_a2[0] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_17_net_1));
    SLE un1_data_out8_17_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_12__1_sqmuxa), .ALn(un1_data_out8_17_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_data_out8_17_set_net_1));
    CFG4 #( .INIT(16'hFFF8) )  \data_out_2_15_i_0_i_11[0]  (.A(
        \mem_5__2_i_0_0_a2[0] ), .B(\mem_5_[0]_net_1 ), .C(
        \data_out_2_15_i_0_i_7[0]_net_1 ), .D(N_641), .Y(
        \data_out_2_15_i_0_i_11[0]_net_1 ));
    CFG3 #( .INIT(8'h02) )  un1_data_out8_98 (.A(\mem_10_[1]_net_1 ), 
        .B(\mem_10__2_i_0_0_a2[0] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_98_net_1));
    SLE un1_data_out8_218_rs (.D(VCC_net_1), .CLK(
        un1_data_out8_114_net_1), .EN(VCC_net_1), .ALn(
        un1_data_out8_218_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(VCC_net_1), .Q(un1_data_out8_218_rs_net_1));
    CFG3 #( .INIT(8'hF2) )  un1_data_out8_202 (.A(\mem_9_[6]_net_1 ), 
        .B(\mem_9__2_i_0_0_a2[0] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_202_i));
    CFG3 #( .INIT(8'hF2) )  un1_data_out8_195 (.A(\mem_5_[4]_net_1 ), 
        .B(\mem_5__2_i_0_0_a2[0] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_195_i));
    CFG3 #( .INIT(8'hF2) )  un1_data_out8_226 (.A(\mem_11_[2]_net_1 ), 
        .B(\mem_11__2_i_0_0_a2[2] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_226_i));
    SLE un1_data_out8_111_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_13__1_sqmuxa), .ALn(un1_data_out8_111_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_data_out8_111_set_net_1));
    CFG1 #( .INIT(2'h1) )  un1_data_out8_110_set_RNO (.A(
        un1_data_out8_110_net_1), .Y(un1_data_out8_110_i));
    SLE un1_data_out8_71_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_8__1_sqmuxa), .ALn(un1_data_out8_71_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_data_out8_71_set_net_1));
    SLE un1_data_out8_192_rs (.D(VCC_net_1), .CLK(
        un1_data_out8_73_net_1), .EN(VCC_net_1), .ALn(
        un1_data_out8_192_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(VCC_net_1), .Q(un1_data_out8_192_rs_net_1));
    SLE un1_data_out8_121_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_3__1_sqmuxa), .ALn(un1_data_out8_121_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_data_out8_121_set_net_1));
    SLE un1_data_out8_45_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_5__1_sqmuxa), .ALn(un1_data_out8_45_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_data_out8_45_set_net_1));
    SLE un1_data_out8_243_rs (.D(VCC_net_1), .CLK(
        un1_data_out8_19_net_1), .EN(VCC_net_1), .ALn(
        un1_data_out8_243_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(VCC_net_1), .Q(un1_data_out8_243_rs_net_1));
    CFG4 #( .INIT(16'h0040) )  \WRITE_GEN.mem_12__2_i_0_0_a2[0]  (.A(
        CoreAPB3_0_APBmslave4_PADDR[2]), .B(
        CoreAPB3_0_APBmslave4_PADDR[5]), .C(
        CoreAPB3_0_APBmslave4_PADDR[4]), .D(
        CoreAPB3_0_APBmslave4_PADDR[3]), .Y(\mem_12__2_i_0_0_a2[0] ));
    SLE un1_data_out8_152_rs (.D(VCC_net_1), .CLK(
        un1_data_out8_9_net_1), .EN(VCC_net_1), .ALn(
        un1_data_out8_152_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(VCC_net_1), .Q(un1_data_out8_152_rs_net_1));
    SLE un1_data_out8_101_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_10__1_sqmuxa), .ALn(un1_data_out8_101_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_data_out8_101_set_net_1));
    SLE \mem_6_[4]  (.D(CoreAPB3_0_APBmslave4_PWDATA[4]), .CLK(
        FCCC_0_GL1), .EN(mem_6__1_sqmuxa), .ALn(un1_data_out8_171_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_6_rs[4] ));
    CFG1 #( .INIT(2'h1) )  un1_data_out8_79_set_RNO (.A(
        un1_data_out8_79_net_1), .Y(un1_data_out8_79_i));
    CFG1 #( .INIT(2'h1) )  un1_data_out8_96_set_RNO (.A(
        un1_data_out8_96_net_1), .Y(un1_data_out8_96_i));
    SLE un1_data_out8_68_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_8__1_sqmuxa), .ALn(un1_data_out8_68_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_data_out8_68_set_net_1));
    CFG1 #( .INIT(2'h1) )  un1_data_out8_7_set_RNO (.A(
        un1_data_out8_7_net_1), .Y(un1_data_out8_7_i));
    CFG3 #( .INIT(8'h02) )  un1_data_out8_93 (.A(\mem_11_[5]_net_1 ), 
        .B(\mem_11__2_i_0_0_a2[2] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_93_net_1));
    CFG4 #( .INIT(16'hECA0) )  \data_out_2_15_i_i_7[5]  (.A(
        \mem_8_[5]_net_1 ), .B(\mem_0_[5]_net_1 ), .C(
        mem_8__2_i_0_0_a2[2]), .D(mem_0__2_i_0_0_a2[0]), .Y(
        \data_out_2_15_i_i_7[5]_net_1 ));
    SLE un1_data_out8_175_rs (.D(VCC_net_1), .CLK(
        un1_data_out8_120_net_1), .EN(VCC_net_1), .ALn(
        un1_data_out8_175_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(VCC_net_1), .Q(un1_data_out8_175_rs_net_1));
    CFG3 #( .INIT(8'hF2) )  un1_data_out8_217 (.A(\mem_14_[1]_net_1 ), 
        .B(\mem_14__2_i_0_0_a2[2] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_217_i));
    CFG3 #( .INIT(8'h02) )  un1_data_out8_8 (.A(\mem_4_[6]_net_1 ), .B(
        \mem_4__2_i_0_0_a2[0] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_8_net_1));
    CFG1 #( .INIT(2'h1) )  un1_data_out8_124_set_RNO (.A(
        un1_data_out8_124_net_1), .Y(un1_data_out8_124_i));
    SLE \data_out[2]  (.D(N_13), .CLK(FCCC_0_GL1), .EN(rd_enable), 
        .ALn(MSS_RESET_N_M2F_c), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(
        CoreAPB3_0_APBmslave5_PRDATA[2]));
    CFG3 #( .INIT(8'h02) )  un1_data_out8_110 (.A(\mem_13_[6]_net_1 ), 
        .B(\mem_13__2_i_0_0_a2[0] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_110_net_1));
    SLE \mem_0_[4]  (.D(CoreAPB3_0_APBmslave4_PWDATA[4]), .CLK(
        FCCC_0_GL1), .EN(mem_0__1_sqmuxa), .ALn(un1_data_out8_148_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_0_rs[4] ));
    CFG3 #( .INIT(8'hF2) )  un1_data_out8_181 (.A(\mem_7_[1]_net_1 ), 
        .B(\mem_7__2_i_0_0_a2[1] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_181_i));
    CFG1 #( .INIT(2'h1) )  un1_data_out8_15_set_RNO (.A(
        un1_data_out8_15_net_1), .Y(un1_data_out8_15_i));
    CFG3 #( .INIT(8'hF8) )  \mem_3__RNI429V[5]  (.A(
        un1_data_out8_51_set_net_1), .B(un1_data_out8_133_rs_net_1), 
        .C(\mem_3_rs[5] ), .Y(\mem_3_[5]_net_1 ));
    SLE un1_data_out8_239_rs (.D(VCC_net_1), .CLK(
        un1_data_out8_64_net_1), .EN(VCC_net_1), .ALn(
        un1_data_out8_239_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(VCC_net_1), .Q(un1_data_out8_239_rs_net_1));
    VCC VCC (.Y(VCC_net_1));
    CFG3 #( .INIT(8'hF2) )  un1_data_out8_246 (.A(\mem_12_[6]_net_1 ), 
        .B(\mem_12__2_i_0_0_a2[0] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_246_i));
    CFG4 #( .INIT(16'hEAC0) )  \data_out_2_15_i_i_0[2]  (.A(
        \mem_10_[2]_net_1 ), .B(\mem_12_[2]_net_1 ), .C(
        \mem_12__2_i_0_0_a2[0] ), .D(\mem_10__2_i_0_0_a2[0] ), .Y(
        \data_out_2_15_i_i_0[2]_net_1 ));
    CFG4 #( .INIT(16'hECA0) )  \data_out_2_15_i_0_i_1[0]  (.A(
        \mem_14_[0]_net_1 ), .B(\mem_9_[0]_net_1 ), .C(
        \mem_14__2_i_0_0_a2[2] ), .D(\mem_9__2_i_0_0_a2[0] ), .Y(
        \data_out_2_15_i_0_i_1[0]_net_1 ));
    CFG4 #( .INIT(16'hECA0) )  \data_out_2_15_i_0_i_5[0]  (.A(
        \mem_1_[0]_net_1 ), .B(\mem_2_[0]_net_1 ), .C(
        \mem_1__2_i_0_0_a2[0] ), .D(\mem_2__2_i_0_0_a2[0] ), .Y(
        \data_out_2_15_i_0_i_5[0]_net_1 ));
    SLE un1_data_out8_200_rs (.D(VCC_net_1), .CLK(
        un1_data_out8_77_net_1), .EN(VCC_net_1), .ALn(
        un1_data_out8_200_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(VCC_net_1), .Q(un1_data_out8_200_rs_net_1));
    CFG3 #( .INIT(8'hF8) )  un1_data_out8_177_rs_RNI0RJG (.A(
        un1_data_out8_122_set_net_1), .B(un1_data_out8_177_rs_net_1), 
        .C(\mem_6_rs[7] ), .Y(\mem_6_[7]_net_1 ));
    SLE un1_data_out8_15_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_1__1_sqmuxa), .ALn(un1_data_out8_15_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_data_out8_15_set_net_1));
    SLE un1_data_out8_142_rs (.D(VCC_net_1), .CLK(
        un1_data_out8_68_net_1), .EN(VCC_net_1), .ALn(
        un1_data_out8_142_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(VCC_net_1), .Q(un1_data_out8_142_rs_net_1));
    CFG1 #( .INIT(2'h1) )  un1_data_out8_85_set_RNO (.A(
        un1_data_out8_85_net_1), .Y(un1_data_out8_85_i));
    CFG3 #( .INIT(8'hF8) )  \mem_7__RNIMSVP[7]  (.A(
        un1_data_out8_1_set_net_1), .B(un1_data_out8_233_rs_net_1), .C(
        \mem_7_rs[7] ), .Y(\mem_7_[7]_net_1 ));
    CFG1 #( .INIT(2'h1) )  un1_data_out8_11_set_RNO (.A(
        un1_data_out8_11_net_1), .Y(un1_data_out8_11_i));
    SLE un1_data_out8_229_rs (.D(VCC_net_1), .CLK(
        un1_data_out8_54_net_1), .EN(VCC_net_1), .ALn(
        un1_data_out8_229_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(VCC_net_1), .Q(un1_data_out8_229_rs_net_1));
    CFG3 #( .INIT(8'h02) )  un1_data_out8_7 (.A(\mem_8_[0]_net_1 ), .B(
        mem_8__2_i_0_0_a2[2]), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_7_net_1));
    CFG3 #( .INIT(8'hF2) )  un1_data_out8_213 (.A(\mem_13_[5]_net_1 ), 
        .B(\mem_13__2_i_0_0_a2[0] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_213_i));
    SLE un1_data_out8_182_rs (.D(VCC_net_1), .CLK(
        un1_data_out8_88_net_1), .EN(VCC_net_1), .ALn(
        un1_data_out8_182_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(VCC_net_1), .Q(un1_data_out8_182_rs_net_1));
    SLE \mem_12_[0]  (.D(CoreAPB3_0_APBmslave4_PWDATA[0]), .CLK(
        FCCC_0_GL1), .EN(mem_12__1_sqmuxa), .ALn(un1_data_out8_238_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_12_rs[0] ));
    SLE un1_data_out8_42_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_1__1_sqmuxa), .ALn(un1_data_out8_42_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_data_out8_42_set_net_1));
    SLE un1_data_out8_214_rs (.D(VCC_net_1), .CLK(
        un1_data_out8_110_net_1), .EN(VCC_net_1), .ALn(
        un1_data_out8_214_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(VCC_net_1), .Q(un1_data_out8_214_rs_net_1));
    SLE \mem_5_[3]  (.D(CoreAPB3_0_APBmslave4_PWDATA[3]), .CLK(
        FCCC_0_GL1), .EN(mem_5__1_sqmuxa), .ALn(un1_data_out8_193_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_5_rs[3] ));
    CFG3 #( .INIT(8'h02) )  un1_data_out8_97 (.A(\mem_10_[0]_net_1 ), 
        .B(\mem_10__2_i_0_0_a2[0] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_97_net_1));
    SLE un1_data_out8_23_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_12__1_sqmuxa), .ALn(un1_data_out8_23_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_data_out8_23_set_net_1));
    CFG3 #( .INIT(8'hF2) )  un1_data_out8_186 (.A(\mem_8_[6]_net_1 ), 
        .B(mem_8__2_i_0_0_a2[2]), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_186_i));
    CFG3 #( .INIT(8'h02) )  un1_data_out8_86 (.A(\mem_0_[6]_net_1 ), 
        .B(mem_0__2_i_0_0_a2[0]), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_86_net_1));
    SLE un1_data_out8_83_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_0__1_sqmuxa), .ALn(un1_data_out8_83_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_data_out8_83_set_net_1));
    CFG3 #( .INIT(8'hF2) )  un1_data_out8_131 (.A(\mem_3_[3]_net_1 ), 
        .B(\mem_3__2_i_0_0_a2[0] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_131_i));
    CFG4 #( .INIT(16'h4000) )  \WRITE_GEN.mem_14__2_i_0_0_a2[2]  (.A(
        CoreAPB3_0_APBmslave4_PADDR[2]), .B(
        CoreAPB3_0_APBmslave4_PADDR[5]), .C(
        CoreAPB3_0_APBmslave4_PADDR[4]), .D(
        CoreAPB3_0_APBmslave4_PADDR[3]), .Y(\mem_14__2_i_0_0_a2[2] ));
    SLE \mem_6_[0]  (.D(CoreAPB3_0_APBmslave4_PWDATA[0]), .CLK(
        FCCC_0_GL1), .EN(mem_6__1_sqmuxa), .ALn(un1_data_out8_203_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_6_rs[0] ));
    CFG1 #( .INIT(2'h1) )  un1_data_out8_23_set_RNO (.A(
        un1_data_out8_23_net_1), .Y(un1_data_out8_23_i));
    SLE un1_data_out8_247_rs (.D(VCC_net_1), .CLK(
        un1_data_out8_23_net_1), .EN(VCC_net_1), .ALn(
        un1_data_out8_247_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(VCC_net_1), .Q(un1_data_out8_247_rs_net_1));
    CFG3 #( .INIT(8'hF2) )  un1_data_out8_164 (.A(\mem_2_[4]_net_1 ), 
        .B(\mem_2__2_i_0_0_a2[0] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_164_i));
    SLE un1_data_out8_118_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_14__1_sqmuxa), .ALn(un1_data_out8_118_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_data_out8_118_set_net_1));
    CFG3 #( .INIT(8'hF2) )  un1_data_out8_199 (.A(\mem_5_[6]_net_1 ), 
        .B(\mem_5__2_i_0_0_a2[0] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_199_i));
    SLE \mem_13_[5]  (.D(CoreAPB3_0_APBmslave4_PWDATA[5]), .CLK(
        FCCC_0_GL1), .EN(mem_13__1_sqmuxa), .ALn(un1_data_out8_213_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_13_rs[5] ));
    CFG1 #( .INIT(2'h1) )  un1_data_out8_81_set_RNO (.A(
        un1_data_out8_81_net_1), .Y(un1_data_out8_81_i));
    CFG3 #( .INIT(8'hF8) )  un1_data_out8_63_set_RNIUGGL (.A(
        un1_data_out8_63_set_net_1), .B(un1_data_out8_253_rs_net_1), 
        .C(\mem_15_rs[6] ), .Y(\mem_15_[6]_net_1 ));
    CFG3 #( .INIT(8'hF8) )  un1_data_out8_151_rs_RNIC10H (.A(
        un1_data_out8_87_set_net_1), .B(un1_data_out8_151_rs_net_1), 
        .C(\mem_0_rs[7] ), .Y(\mem_0_[7]_net_1 ));
    CFG3 #( .INIT(8'h02) )  un1_data_out8_113 (.A(\mem_14_[1]_net_1 ), 
        .B(\mem_14__2_i_0_0_a2[2] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_113_net_1));
    SLE un1_data_out8_108_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_13__1_sqmuxa), .ALn(un1_data_out8_108_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_data_out8_108_set_net_1));
    SLE un1_data_out8_24_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_5__1_sqmuxa), .ALn(un1_data_out8_24_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_data_out8_24_set_net_1));
    SLE un1_data_out8_84_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_0__1_sqmuxa), .ALn(un1_data_out8_84_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_data_out8_84_set_net_1));
    SLE \mem_0_[0]  (.D(CoreAPB3_0_APBmslave4_PWDATA[0]), .CLK(
        FCCC_0_GL1), .EN(mem_0__1_sqmuxa), .ALn(un1_data_out8_147_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_0_rs[0] ));
    CFG3 #( .INIT(8'hF8) )  un1_data_out8_179_rs_RNIU5CF (.A(
        un1_data_out8_124_set_net_1), .B(un1_data_out8_179_rs_net_1), 
        .C(\mem_7_rs[0] ), .Y(\mem_7_[0]_net_1 ));
    SLE \mem_1_[4]  (.D(CoreAPB3_0_APBmslave4_PWDATA[4]), .CLK(
        FCCC_0_GL1), .EN(mem_1__1_sqmuxa), .ALn(un1_data_out8_156_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_1_rs[4] ));
    CFG4 #( .INIT(16'hECA0) )  \data_out_2_15_i_0_i_5[1]  (.A(
        \mem_6_[1]_net_1 ), .B(\mem_1_[1]_net_1 ), .C(
        \mem_6__2_i_0_0_a2[2] ), .D(\mem_1__2_i_0_0_a2[0] ), .Y(
        \data_out_2_15_i_0_i_5[1]_net_1 ));
    CFG3 #( .INIT(8'hF2) )  un1_data_out8_136 (.A(\mem_4_[0]_net_1 ), 
        .B(\mem_4__2_i_0_0_a2[0] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_136_i));
    SLE un1_data_out8_117_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_14__1_sqmuxa), .ALn(un1_data_out8_117_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_data_out8_117_set_net_1));
    CFG2 #( .INIT(4'h8) )  \data_out_2_15_i_i_a3_8[4]  (.A(
        \mem_3__2_i_0_0_a2[0] ), .B(\mem_3_[4]_net_1 ), .Y(
        \data_out_2_15_i_i_a3_8[4]_net_1 ));
    SLE \mem_9_[4]  (.D(CoreAPB3_0_APBmslave4_PWDATA[4]), .CLK(
        FCCC_0_GL1), .EN(mem_9__1_sqmuxa), .ALn(un1_data_out8_198_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_9_rs[4] ));
    CFG3 #( .INIT(8'h02) )  un1_data_out8_76 (.A(\mem_9_[4]_net_1 ), 
        .B(\mem_9__2_i_0_0_a2[0] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_76_net_1));
    SLE un1_data_out8_73_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_9__1_sqmuxa), .ALn(un1_data_out8_73_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_data_out8_73_set_net_1));
    CFG4 #( .INIT(16'hFFFE) )  \data_out_2_15_i_0_i[3]  (.A(
        \data_out_2_15_i_0_i_4[3]_net_1 ), .B(
        \data_out_2_15_i_0_i_5[3]_net_1 ), .C(
        \data_out_2_15_i_0_i_12[3]_net_1 ), .D(
        \data_out_2_15_i_0_i_11[3]_net_1 ), .Y(N_7));
    SLE \mem_13_[1]  (.D(CoreAPB3_0_APBmslave4_PWDATA[1]), .CLK(
        FCCC_0_GL1), .EN(mem_13__1_sqmuxa), .ALn(un1_data_out8_209_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_13_rs[1] ));
    SLE \mem_11_[5]  (.D(CoreAPB3_0_APBmslave4_PWDATA[5]), .CLK(
        FCCC_0_GL1), .EN(mem_11__1_sqmuxa), .ALn(un1_data_out8_232_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_11_rs[5] ));
    SLE un1_data_out8_127_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_3__1_sqmuxa), .ALn(un1_data_out8_127_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_data_out8_127_set_net_1));
    CFG4 #( .INIT(16'hEAC0) )  \data_out_2_15_i_i_2[5]  (.A(
        \mem_13_[5]_net_1 ), .B(\mem_11_[5]_net_1 ), .C(
        \mem_11__2_i_0_0_a2[2] ), .D(\mem_13__2_i_0_0_a2[0] ), .Y(
        \data_out_2_15_i_i_2[5]_net_1 ));
    CFG3 #( .INIT(8'hF8) )  un1_data_out8_90_set_RNIMSQD (.A(
        un1_data_out8_90_set_net_1), .B(un1_data_out8_226_rs_net_1), 
        .C(\mem_11_rs[2] ), .Y(\mem_11_[2]_net_1 ));
    CFG2 #( .INIT(4'h8) )  \data_out_2_15_i_0_i_a3_8[1]  (.A(
        \mem_3__2_i_0_0_a2[0] ), .B(\mem_3_[1]_net_1 ), .Y(N_413));
    SLE un1_data_out8_107_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_13__1_sqmuxa), .ALn(un1_data_out8_107_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_data_out8_107_set_net_1));
    CFG3 #( .INIT(8'hF2) )  un1_data_out8_205 (.A(\mem_6_[1]_net_1 ), 
        .B(\mem_6__2_i_0_0_a2[2] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_205_i));
    SLE un1_data_out8_12_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_5__1_sqmuxa), .ALn(un1_data_out8_12_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_data_out8_12_set_net_1));
    CFG3 #( .INIT(8'hF2) )  un1_data_out8_171 (.A(\mem_6_[4]_net_1 ), 
        .B(\mem_6__2_i_0_0_a2[2] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_171_i));
    CFG2 #( .INIT(4'h8) )  mem_13__1_sqmuxa_0_a3_0_a3 (.A(
        mem_14__1_sqmuxa_0_a2_0_a3_0_a2_net_1), .B(
        \mem_13__2_i_0_0_a2[0] ), .Y(mem_13__1_sqmuxa));
    SLE un1_data_out8_74_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_9__1_sqmuxa), .ALn(un1_data_out8_74_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_data_out8_74_set_net_1));
    CFG3 #( .INIT(8'h02) )  un1_data_out8_80 (.A(\mem_0_[0]_net_1 ), 
        .B(mem_0__2_i_0_0_a2[0]), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_80_net_1));
    SLE \mem_11_[1]  (.D(CoreAPB3_0_APBmslave4_PWDATA[1]), .CLK(
        FCCC_0_GL1), .EN(mem_11__1_sqmuxa), .ALn(un1_data_out8_224_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_11_rs[1] ));
    CFG1 #( .INIT(2'h1) )  un1_data_out8_19_set_RNO (.A(
        un1_data_out8_19_net_1), .Y(un1_data_out8_19_i));
    CFG3 #( .INIT(8'hF8) )  \mem_2__RNI39LF[1]  (.A(
        un1_data_out8_27_set_net_1), .B(un1_data_out8_161_rs_net_1), 
        .C(\mem_2_rs[1] ), .Y(\mem_2_[1]_net_1 ));
    CFG3 #( .INIT(8'h02) )  un1_data_out8_104 (.A(\mem_13_[0]_net_1 ), 
        .B(\mem_13__2_i_0_0_a2[0] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_104_net_1));
    CFG4 #( .INIT(16'hECA0) )  \data_out_2_15_i_0_i_5[7]  (.A(
        \mem_6_[7]_net_1 ), .B(\mem_1_[7]_net_1 ), .C(
        \mem_6__2_i_0_0_a2[2] ), .D(\mem_1__2_i_0_0_a2[0] ), .Y(
        \data_out_2_15_i_0_i_5[7]_net_1 ));
    CFG3 #( .INIT(8'hF2) )  un1_data_out8_198 (.A(\mem_9_[4]_net_1 ), 
        .B(\mem_9__2_i_0_0_a2[0] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_198_i));
    CFG4 #( .INIT(16'hFFFE) )  \data_out_2_15_i_i[5]  (.A(
        \data_out_2_15_i_i_4[5]_net_1 ), .B(
        \data_out_2_15_i_i_5[5]_net_1 ), .C(
        \data_out_2_15_i_i_12[5]_net_1 ), .D(
        \data_out_2_15_i_i_11[5]_net_1 ), .Y(N_17));
    CFG3 #( .INIT(8'h02) )  un1_data_out8_19 (.A(\mem_12_[3]_net_1 ), 
        .B(\mem_12__2_i_0_0_a2[0] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_19_net_1));
    CFG1 #( .INIT(2'h1) )  un1_data_out8_93_set_RNO (.A(
        un1_data_out8_93_net_1), .Y(un1_data_out8_93_i));
    CFG3 #( .INIT(8'h02) )  un1_data_out8_68 (.A(\mem_8_[4]_net_1 ), 
        .B(mem_8__2_i_0_0_a2[2]), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_68_net_1));
    CFG3 #( .INIT(8'hF2) )  un1_data_out8_219 (.A(\mem_14_[3]_net_1 ), 
        .B(\mem_14__2_i_0_0_a2[2] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_219_i));
    CFG3 #( .INIT(8'hF2) )  un1_data_out8_176 (.A(\mem_10_[5]_net_1 ), 
        .B(\mem_10__2_i_0_0_a2[0] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_176_i));
    CFG1 #( .INIT(2'h1) )  un1_data_out8_89_set_RNO (.A(
        un1_data_out8_89_net_1), .Y(un1_data_out8_89_i));
    CFG3 #( .INIT(8'h02) )  un1_data_out8_21 (.A(\mem_12_[5]_net_1 ), 
        .B(\mem_12__2_i_0_0_a2[0] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_21_net_1));
    CFG4 #( .INIT(16'hFFFE) )  \data_out_2_15_i_0_i_12[0]  (.A(
        \data_out_2_15_i_0_i_2[0]_net_1 ), .B(
        \data_out_2_15_i_0_i_1[0]_net_1 ), .C(
        \data_out_2_15_i_0_i_3[0]_net_1 ), .D(
        \data_out_2_15_i_0_i_0[0]_net_1 ), .Y(
        \data_out_2_15_i_0_i_12[0]_net_1 ));
    SLE \mem_1_[0]  (.D(CoreAPB3_0_APBmslave4_PWDATA[0]), .CLK(
        FCCC_0_GL1), .EN(mem_1__1_sqmuxa), .ALn(un1_data_out8_152_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_1_rs[0] ));
    CFG4 #( .INIT(16'hECA0) )  \data_out_2_15_i_i_7[4]  (.A(
        \mem_8_[4]_net_1 ), .B(\mem_0_[4]_net_1 ), .C(
        mem_8__2_i_0_0_a2[2]), .D(mem_0__2_i_0_0_a2[0]), .Y(
        \data_out_2_15_i_i_7[4]_net_1 ));
    CFG4 #( .INIT(16'hFFFE) )  \data_out_2_15_i_i_12[4]  (.A(
        \data_out_2_15_i_i_2[4]_net_1 ), .B(
        \data_out_2_15_i_i_1[4]_net_1 ), .C(
        \data_out_2_15_i_i_3[4]_net_1 ), .D(
        \data_out_2_15_i_i_0[4]_net_1 ), .Y(
        \data_out_2_15_i_i_12[4]_net_1 ));
    CFG3 #( .INIT(8'h02) )  un1_data_out8_70 (.A(\mem_8_[6]_net_1 ), 
        .B(mem_8__2_i_0_0_a2[2]), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_70_net_1));
    CFG4 #( .INIT(16'h0200) )  \WRITE_GEN.mem_3__2_i_0_0_a2[0]  (.A(
        CoreAPB3_0_APBmslave4_PADDR[2]), .B(
        CoreAPB3_0_APBmslave4_PADDR[5]), .C(
        CoreAPB3_0_APBmslave4_PADDR[4]), .D(
        CoreAPB3_0_APBmslave4_PADDR[3]), .Y(\mem_3__2_i_0_0_a2[0] ));
    SLE \mem_9_[0]  (.D(CoreAPB3_0_APBmslave4_PWDATA[0]), .CLK(
        FCCC_0_GL1), .EN(mem_9__1_sqmuxa), .ALn(un1_data_out8_190_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_9_rs[0] ));
    SLE un1_data_out8_130_rs (.D(VCC_net_1), .CLK(
        un1_data_out8_125_net_1), .EN(VCC_net_1), .ALn(
        un1_data_out8_130_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(VCC_net_1), .Q(un1_data_out8_130_rs_net_1));
    SLE \mem_15_[3]  (.D(CoreAPB3_0_APBmslave4_PWDATA[3]), .CLK(
        FCCC_0_GL1), .EN(mem_15__1_sqmuxa), .ALn(un1_data_out8_250_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_15_rs[3] ));
    SLE \mem_14_[4]  (.D(CoreAPB3_0_APBmslave4_PWDATA[4]), .CLK(
        FCCC_0_GL1), .EN(mem_14__1_sqmuxa), .ALn(un1_data_out8_220_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_14_rs[4] ));
    SLE un1_data_out8_50_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_7__1_sqmuxa), .ALn(un1_data_out8_50_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_data_out8_50_set_net_1));
    CFG3 #( .INIT(8'h02) )  un1_data_out8_41 (.A(\mem_5_[3]_net_1 ), 
        .B(\mem_5__2_i_0_0_a2[0] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_41_net_1));
    CFG3 #( .INIT(8'h02) )  un1_data_out8_122 (.A(\mem_6_[7]_net_1 ), 
        .B(\mem_6__2_i_0_0_a2[2] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_122_net_1));
    SLE un1_data_out8_28_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_6__1_sqmuxa), .ALn(un1_data_out8_28_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_data_out8_28_set_net_1));
    SLE un1_data_out8_88_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_11__1_sqmuxa), .ALn(un1_data_out8_88_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_data_out8_88_set_net_1));
    CFG3 #( .INIT(8'h02) )  un1_data_out8_63 (.A(\mem_15_[6]_net_1 ), 
        .B(\mem_15__2_i_0_0_a2[0] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_63_net_1));
    CFG4 #( .INIT(16'hFFF8) )  \data_out_2_15_i_0_i_11[1]  (.A(
        \mem_5__2_i_0_0_a2[0] ), .B(\mem_5_[1]_net_1 ), .C(
        \data_out_2_15_i_0_i_7[1]_net_1 ), .D(N_413), .Y(
        \data_out_2_15_i_0_i_11[1]_net_1 ));
    SLE un1_data_out8_206_rs (.D(VCC_net_1), .CLK(
        un1_data_out8_97_net_1), .EN(VCC_net_1), .ALn(
        un1_data_out8_206_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(VCC_net_1), .Q(un1_data_out8_206_rs_net_1));
    SLE \mem_10_[2]  (.D(CoreAPB3_0_APBmslave4_PWDATA[2]), .CLK(
        FCCC_0_GL1), .EN(mem_10__1_sqmuxa), .ALn(un1_data_out8_170_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_10_rs[2] ));
    CFG4 #( .INIT(16'h0100) )  \WRITE_GEN.mem_2__2_i_0_0_a2[0]  (.A(
        CoreAPB3_0_APBmslave4_PADDR[2]), .B(
        CoreAPB3_0_APBmslave4_PADDR[5]), .C(
        CoreAPB3_0_APBmslave4_PADDR[4]), .D(
        CoreAPB3_0_APBmslave4_PADDR[3]), .Y(\mem_2__2_i_0_0_a2[0] ));
    CFG3 #( .INIT(8'hF8) )  un1_data_out8_194_rs_RNIJ8S31 (.A(
        un1_data_out8_74_set_net_1), .B(un1_data_out8_194_rs_net_1), 
        .C(\mem_9_rs[2] ), .Y(\mem_9_[2]_net_1 ));
    CFG4 #( .INIT(16'hEAC0) )  \data_out_2_15_i_0_i_3[7]  (.A(
        \mem_15_[7]_net_1 ), .B(\mem_7_[7]_net_1 ), .C(
        \mem_7__2_i_0_0_a2[1] ), .D(\mem_15__2_i_0_0_a2[0] ), .Y(
        \data_out_2_15_i_0_i_3[7]_net_1 ));
    CFG3 #( .INIT(8'hF8) )  \mem_10__RNIAAIG[6]  (.A(
        un1_data_out8_103_set_net_1), .B(un1_data_out8_178_rs_net_1), 
        .C(\mem_10_rs[6] ), .Y(\mem_10_[6]_net_1 ));
    SLE un1_data_out8_162_rs (.D(VCC_net_1), .CLK(
        un1_data_out8_29_net_1), .EN(VCC_net_1), .ALn(
        un1_data_out8_162_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(VCC_net_1), .Q(un1_data_out8_162_rs_net_1));
    CFG3 #( .INIT(8'hF8) )  un1_data_out8_144_rs_RNI28UM (.A(
        un1_data_out8_81_set_net_1), .B(un1_data_out8_144_rs_net_1), 
        .C(\mem_0_rs[1] ), .Y(\mem_0_[1]_net_1 ));
    SLE \mem_3_[2]  (.D(CoreAPB3_0_APBmslave4_PWDATA[2]), .CLK(
        FCCC_0_GL1), .EN(mem_3__1_sqmuxa), .ALn(un1_data_out8_130_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_3_rs[2] ));
    CFG4 #( .INIT(16'hEAC0) )  \data_out_2_15_i_0_i_3[3]  (.A(
        \mem_15_[3]_net_1 ), .B(\mem_7_[3]_net_1 ), .C(
        \mem_7__2_i_0_0_a2[1] ), .D(\mem_15__2_i_0_0_a2[0] ), .Y(
        \data_out_2_15_i_0_i_3[3]_net_1 ));
    SLE un1_data_out8_116_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_14__1_sqmuxa), .ALn(un1_data_out8_116_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_data_out8_116_set_net_1));
    SLE un1_data_out8_213_rs (.D(VCC_net_1), .CLK(
        un1_data_out8_109_net_1), .EN(VCC_net_1), .ALn(
        un1_data_out8_213_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(VCC_net_1), .Q(un1_data_out8_213_rs_net_1));
    CFG3 #( .INIT(8'hF2) )  un1_data_out8_152 (.A(\mem_1_[0]_net_1 ), 
        .B(\mem_1__2_i_0_0_a2[0] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_152_i));
    SLE \mem_14_[6]  (.D(CoreAPB3_0_APBmslave4_PWDATA[6]), .CLK(
        FCCC_0_GL1), .EN(mem_14__1_sqmuxa), .ALn(un1_data_out8_222_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_14_rs[6] ));
    CFG2 #( .INIT(4'h8) )  mem_1__1_sqmuxa_0_a3_0_a3 (.A(
        mem_14__1_sqmuxa_0_a2_0_a3_0_a2_net_1), .B(
        \mem_1__2_i_0_0_a2[0] ), .Y(mem_1__1_sqmuxa));
    CFG3 #( .INIT(8'h02) )  un1_data_out8_58 (.A(\mem_15_[1]_net_1 ), 
        .B(\mem_15__2_i_0_0_a2[0] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_58_net_1));
    CFG1 #( .INIT(2'h1) )  un1_data_out8_2_set_RNO (.A(
        un1_data_out8_2_net_1), .Y(un1_data_out8_2_i));
    CFG3 #( .INIT(8'hF2) )  un1_data_out8_201 (.A(\mem_5_[7]_net_1 ), 
        .B(\mem_5__2_i_0_0_a2[0] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_201_i));
    SLE un1_data_out8_126_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_7__1_sqmuxa), .ALn(un1_data_out8_126_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_data_out8_126_set_net_1));
    SLE un1_data_out8_46_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_1__1_sqmuxa), .ALn(un1_data_out8_46_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_data_out8_46_set_net_1));
    SLE un1_data_out8_78_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_9__1_sqmuxa), .ALn(un1_data_out8_78_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_data_out8_78_set_net_1));
    SLE un1_data_out8_37_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_2__1_sqmuxa), .ALn(un1_data_out8_37_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_data_out8_37_set_net_1));
    CFG3 #( .INIT(8'hF8) )  \mem_2__RNIIEUO[7]  (.A(
        un1_data_out8_39_set_net_1), .B(un1_data_out8_167_rs_net_1), 
        .C(\mem_2_rs[7] ), .Y(\mem_2_[7]_net_1 ));
    CFG3 #( .INIT(8'hF2) )  un1_data_out8_160 (.A(\mem_2_[0]_net_1 ), 
        .B(\mem_2__2_i_0_0_a2[0] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_160_i));
    SLE un1_data_out8_106_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_13__1_sqmuxa), .ALn(un1_data_out8_106_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_data_out8_106_set_net_1));
    CFG4 #( .INIT(16'hFFFE) )  \data_out_2_15_i_0_i[0]  (.A(
        \data_out_2_15_i_0_i_4[0]_net_1 ), .B(
        \data_out_2_15_i_0_i_5[0]_net_1 ), .C(
        \data_out_2_15_i_0_i_12[0]_net_1 ), .D(
        \data_out_2_15_i_0_i_11[0]_net_1 ), .Y(N_11));
    SLE \mem_8_[7]  (.D(CoreAPB3_0_APBmslave4_PWDATA[7]), .CLK(
        FCCC_0_GL1), .EN(mem_8__1_sqmuxa), .ALn(un1_data_out8_188_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_8_rs[7] ));
    CFG3 #( .INIT(8'hF8) )  un1_data_out8_45_set_RNIJPKR (.A(
        un1_data_out8_45_set_net_1), .B(un1_data_out8_197_rs_net_1), 
        .C(\mem_5_rs[5] ), .Y(\mem_5_[5]_net_1 ));
    SLE \mem_5_[4]  (.D(CoreAPB3_0_APBmslave4_PWDATA[4]), .CLK(
        FCCC_0_GL1), .EN(mem_5__1_sqmuxa), .ALn(un1_data_out8_195_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_5_rs[4] ));
    CFG3 #( .INIT(8'hF2) )  un1_data_out8_142 (.A(\mem_8_[4]_net_1 ), 
        .B(mem_8__2_i_0_0_a2[2]), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_142_i));
    CFG3 #( .INIT(8'h02) )  un1_data_out8_67 (.A(\mem_4_[5]_net_1 ), 
        .B(\mem_4__2_i_0_0_a2[0] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_67_net_1));
    SLE \data_out[1]  (.D(N_9), .CLK(FCCC_0_GL1), .EN(rd_enable), .ALn(
        MSS_RESET_N_M2F_c), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(GND_net_1), .Q(
        CoreAPB3_0_APBmslave5_PRDATA[1]));
    SLE \mem_8_[5]  (.D(CoreAPB3_0_APBmslave4_PWDATA[5]), .CLK(
        FCCC_0_GL1), .EN(mem_8__1_sqmuxa), .ALn(un1_data_out8_184_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_8_rs[5] ));
    CFG3 #( .INIT(8'h02) )  un1_data_out8_99 (.A(\mem_10_[2]_net_1 ), 
        .B(\mem_10__2_i_0_0_a2[0] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_99_net_1));
    CFG3 #( .INIT(8'hF8) )  un1_data_out8_71_set_RNIN5AJ (.A(
        un1_data_out8_71_set_net_1), .B(un1_data_out8_188_rs_net_1), 
        .C(\mem_8_rs[7] ), .Y(\mem_8_[7]_net_1 ));
    CFG3 #( .INIT(8'h02) )  un1_data_out8_53 (.A(\mem_3_[6]_net_1 ), 
        .B(\mem_3__2_i_0_0_a2[0] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_53_net_1));
    SLE un1_data_out8_231_rs (.D(VCC_net_1), .CLK(
        un1_data_out8_3_net_1), .EN(VCC_net_1), .ALn(
        un1_data_out8_231_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(VCC_net_1), .Q(un1_data_out8_231_rs_net_1));
    CFG3 #( .INIT(8'hF8) )  un1_data_out8_24_set_RNIJI051 (.A(
        un1_data_out8_24_set_net_1), .B(un1_data_out8_199_rs_net_1), 
        .C(\mem_5_rs[6] ), .Y(\mem_5_[6]_net_1 ));
    CFG4 #( .INIT(16'hEAC0) )  \data_out_2_15_i_0_i_3[1]  (.A(
        \mem_15_[1]_net_1 ), .B(\mem_7_[1]_net_1 ), .C(
        \mem_7__2_i_0_0_a2[1] ), .D(\mem_15__2_i_0_0_a2[0] ), .Y(
        \data_out_2_15_i_0_i_3[1]_net_1 ));
    CFG3 #( .INIT(8'hF8) )  \mem_15__RNIR8701[5]  (.A(
        un1_data_out8_62_set_net_1), .B(un1_data_out8_252_rs_net_1), 
        .C(\mem_15_rs[5] ), .Y(\mem_15_[5]_net_1 ));
    CFG4 #( .INIT(16'hFFFE) )  \data_out_2_15_i_i[2]  (.A(
        \data_out_2_15_i_i_4[2]_net_1 ), .B(
        \data_out_2_15_i_i_5[2]_net_1 ), .C(
        \data_out_2_15_i_i_12[2]_net_1 ), .D(
        \data_out_2_15_i_i_11[2]_net_1 ), .Y(N_13));
    CFG3 #( .INIT(8'h02) )  un1_data_out8_127 (.A(\mem_3_[3]_net_1 ), 
        .B(\mem_3__2_i_0_0_a2[0] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_127_net_1));
    CFG1 #( .INIT(2'h1) )  un1_data_out8_8_set_RNO (.A(
        un1_data_out8_8_net_1), .Y(un1_data_out8_8_i));
    CFG1 #( .INIT(2'h1) )  un1_data_out8_109_set_RNO (.A(
        un1_data_out8_109_net_1), .Y(un1_data_out8_109_i));
    CFG3 #( .INIT(8'hF2) )  un1_data_out8_216 (.A(\mem_14_[0]_net_1 ), 
        .B(\mem_14__2_i_0_0_a2[2] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_216_i));
    CFG3 #( .INIT(8'hF8) )  un1_data_out8_15_set_RNI42VO (.A(
        un1_data_out8_15_set_net_1), .B(un1_data_out8_155_rs_net_1), 
        .C(\mem_1_rs[3] ), .Y(\mem_1_[3]_net_1 ));
    CFG2 #( .INIT(4'h8) )  \data_out_2_15_i_0_i_a3_8[0]  (.A(
        \mem_3__2_i_0_0_a2[0] ), .B(\mem_3_[0]_net_1 ), .Y(N_641));
    CFG4 #( .INIT(16'hEAC0) )  \data_out_2_15_i_0_i_4[7]  (.A(
        \mem_4_[7]_net_1 ), .B(\mem_2_[7]_net_1 ), .C(
        \mem_2__2_i_0_0_a2[0] ), .D(\mem_4__2_i_0_0_a2[0] ), .Y(
        \data_out_2_15_i_0_i_4[7]_net_1 ));
    SLE un1_data_out8_221_rs (.D(VCC_net_1), .CLK(
        un1_data_out8_117_net_1), .EN(VCC_net_1), .ALn(
        un1_data_out8_221_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(VCC_net_1), .Q(un1_data_out8_221_rs_net_1));
    SLE un1_data_out8_16_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_12__1_sqmuxa), .ALn(un1_data_out8_16_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_data_out8_16_set_net_1));
    SLE un1_data_out8_60_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_15__1_sqmuxa), .ALn(un1_data_out8_60_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_data_out8_60_set_net_1));
    CFG3 #( .INIT(8'hF2) )  un1_data_out8_230 (.A(\mem_11_[4]_net_1 ), 
        .B(\mem_11__2_i_0_0_a2[2] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_230_i));
    SLE un1_data_out8_249_rs (.D(VCC_net_1), .CLK(
        un1_data_out8_59_net_1), .EN(VCC_net_1), .ALn(
        un1_data_out8_249_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(VCC_net_1), .Q(un1_data_out8_249_rs_net_1));
    CFG3 #( .INIT(8'h02) )  un1_data_out8 (.A(\mem_4_[0]_net_1 ), .B(
        \mem_4__2_i_0_0_a2[0] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_net_1));
    CFG3 #( .INIT(8'hF8) )  \mem_10__RNI2KPJ[4]  (.A(
        un1_data_out8_101_set_net_1), .B(un1_data_out8_174_rs_net_1), 
        .C(\mem_10_rs[4] ), .Y(\mem_10_[4]_net_1 ));
    CFG3 #( .INIT(8'hF2) )  un1_data_out8_207 (.A(\mem_6_[2]_net_1 ), 
        .B(\mem_6__2_i_0_0_a2[2] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_207_i));
    CFG1 #( .INIT(2'h1) )  un1_data_out8_25_set_RNO (.A(
        un1_data_out8_25_net_1), .Y(un1_data_out8_25_i));
    SLE un1_data_out8_217_rs (.D(VCC_net_1), .CLK(
        un1_data_out8_113_net_1), .EN(VCC_net_1), .ALn(
        un1_data_out8_217_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(VCC_net_1), .Q(un1_data_out8_217_rs_net_1));
    CFG3 #( .INIT(8'hF8) )  un1_data_out8_255_rs_RNISCAF (.A(
        un1_data_out8_61_set_net_1), .B(un1_data_out8_255_rs_net_1), 
        .C(\mem_15_rs[4] ), .Y(\mem_15_[4]_net_1 ));
    CFG3 #( .INIT(8'hF2) )  un1_data_out8_163 (.A(\mem_2_[3]_net_1 ), 
        .B(\mem_2__2_i_0_0_a2[0] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_163_i));
    CFG3 #( .INIT(8'hF8) )  un1_data_out8_109_set_RNI8BV11 (.A(
        un1_data_out8_109_set_net_1), .B(un1_data_out8_213_rs_net_1), 
        .C(\mem_13_rs[5] ), .Y(\mem_13_[5]_net_1 ));
    CFG3 #( .INIT(8'h02) )  un1_data_out8_100 (.A(\mem_10_[7]_net_1 ), 
        .B(\mem_10__2_i_0_0_a2[0] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_100_net_1));
    CFG3 #( .INIT(8'hF8) )  \mem_14__RNIAK9M[3]  (.A(
        un1_data_out8_115_set_net_1), .B(un1_data_out8_219_rs_net_1), 
        .C(\mem_14_rs[3] ), .Y(\mem_14_[3]_net_1 ));
    CFG3 #( .INIT(8'hF8) )  \mem_10__RNISK1P[3]  (.A(
        un1_data_out8_96_set_net_1), .B(un1_data_out8_172_rs_net_1), 
        .C(\mem_10_rs[3] ), .Y(\mem_10_[3]_net_1 ));
    CFG3 #( .INIT(8'hF2) )  un1_data_out8_157 (.A(\mem_1_[5]_net_1 ), 
        .B(\mem_1__2_i_0_0_a2[0] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_157_i));
    CFG4 #( .INIT(16'h0002) )  \WRITE_GEN.mem_1__2_i_0_0_a2[0]  (.A(
        CoreAPB3_0_APBmslave4_PADDR[2]), .B(
        CoreAPB3_0_APBmslave4_PADDR[5]), .C(
        CoreAPB3_0_APBmslave4_PADDR[4]), .D(
        CoreAPB3_0_APBmslave4_PADDR[3]), .Y(\mem_1__2_i_0_0_a2[0] ));
    SLE \mem_5_[0]  (.D(CoreAPB3_0_APBmslave4_PWDATA[0]), .CLK(
        FCCC_0_GL1), .EN(mem_5__1_sqmuxa), .ALn(un1_data_out8_187_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_5_rs[0] ));
    CFG3 #( .INIT(8'hF2) )  un1_data_out8_191 (.A(\mem_5_[2]_net_1 ), 
        .B(\mem_5__2_i_0_0_a2[0] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_191_i));
    CFG3 #( .INIT(8'hF8) )  un1_data_out8_176_rs_RNI6V5A (.A(
        un1_data_out8_102_set_net_1), .B(un1_data_out8_176_rs_net_1), 
        .C(\mem_10_rs[5] ), .Y(\mem_10_[5]_net_1 ));
    CFG3 #( .INIT(8'hF8) )  un1_data_out8_225_rs_RNI7J5K (.A(
        un1_data_out8_50_set_net_1), .B(un1_data_out8_225_rs_net_1), 
        .C(\mem_7_rs[3] ), .Y(\mem_7_[3]_net_1 ));
    CFG3 #( .INIT(8'h02) )  un1_data_out8_57 (.A(\mem_15_[0]_net_1 ), 
        .B(\mem_15__2_i_0_0_a2[0] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_57_net_1));
    SLE \mem_3_[1]  (.D(CoreAPB3_0_APBmslave4_PWDATA[1]), .CLK(
        FCCC_0_GL1), .EN(mem_3__1_sqmuxa), .ALn(un1_data_out8_129_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_3_rs[1] ));
    CFG1 #( .INIT(2'h1) )  un1_data_out8_70_set_RNO (.A(
        un1_data_out8_70_net_1), .Y(un1_data_out8_70_i));
    CFG1 #( .INIT(2'h1) )  un1_data_out8_6_set_RNO (.A(
        un1_data_out8_6_net_1), .Y(un1_data_out8_6_i));
    SLE un1_data_out8_35_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_2__1_sqmuxa), .ALn(un1_data_out8_35_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_data_out8_35_set_net_1));
    CFG1 #( .INIT(2'h1) )  un1_data_out8_21_set_RNO (.A(
        un1_data_out8_21_net_1), .Y(un1_data_out8_21_i));
    CFG3 #( .INIT(8'h02) )  un1_data_out8_2 (.A(\mem_4_[1]_net_1 ), .B(
        \mem_4__2_i_0_0_a2[0] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_2_net_1));
    CFG3 #( .INIT(8'hF2) )  un1_data_out8_147 (.A(\mem_0_[0]_net_1 ), 
        .B(mem_0__2_i_0_0_a2[0]), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_147_i));
    CFG1 #( .INIT(2'h1) )  un1_data_out8_121_set_RNO (.A(
        un1_data_out8_121_net_1), .Y(un1_data_out8_121_i));
    CFG1 #( .INIT(2'h1) )  un1_data_out8_78_set_RNO (.A(
        un1_data_out8_78_net_1), .Y(un1_data_out8_78_i));
    CFG3 #( .INIT(8'hF2) )  un1_data_out8_203 (.A(\mem_6_[0]_net_1 ), 
        .B(\mem_6__2_i_0_0_a2[2] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_203_i));
    CFG3 #( .INIT(8'hF8) )  \mem_11__RNI1QVM[7]  (.A(
        un1_data_out8_95_set_net_1), .B(un1_data_out8_236_rs_net_1), 
        .C(\mem_11_rs[7] ), .Y(\mem_11_[7]_net_1 ));
    SLE \mem_10_[7]  (.D(CoreAPB3_0_APBmslave4_PWDATA[7]), .CLK(
        FCCC_0_GL1), .EN(mem_10__1_sqmuxa), .ALn(un1_data_out8_180_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_10_rs[7] ));
    CFG3 #( .INIT(8'h02) )  un1_data_out8_4 (.A(\mem_4_[2]_net_1 ), .B(
        \mem_4__2_i_0_0_a2[0] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_4_net_1));
    CFG3 #( .INIT(8'hF2) )  un1_data_out8_196 (.A(\mem_9_[3]_net_1 ), 
        .B(\mem_9__2_i_0_0_a2[0] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_196_i));
    SLE \mem_15_[0]  (.D(CoreAPB3_0_APBmslave4_PWDATA[0]), .CLK(
        FCCC_0_GL1), .EN(mem_15__1_sqmuxa), .ALn(un1_data_out8_251_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_15_rs[0] ));
    SLE un1_data_out8_172_rs (.D(VCC_net_1), .CLK(
        un1_data_out8_96_net_1), .EN(VCC_net_1), .ALn(
        un1_data_out8_172_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(VCC_net_1), .Q(un1_data_out8_172_rs_net_1));
    SLE un1_data_out8_232_rs (.D(VCC_net_1), .CLK(
        un1_data_out8_93_net_1), .EN(VCC_net_1), .ALn(
        un1_data_out8_232_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(VCC_net_1), .Q(un1_data_out8_232_rs_net_1));
    SLE un1_data_out8_190_rs (.D(VCC_net_1), .CLK(
        un1_data_out8_72_net_1), .EN(VCC_net_1), .ALn(
        un1_data_out8_190_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(VCC_net_1), .Q(un1_data_out8_190_rs_net_1));
    CFG3 #( .INIT(8'h02) )  un1_data_out8_103 (.A(\mem_10_[6]_net_1 ), 
        .B(\mem_10__2_i_0_0_a2[0] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_103_net_1));
    CFG4 #( .INIT(16'hFFF8) )  \data_out_2_15_i_i_11[6]  (.A(
        \mem_5__2_i_0_0_a2[0] ), .B(\mem_5_[6]_net_1 ), .C(
        \data_out_2_15_i_i_7[6]_net_1 ), .D(
        \data_out_2_15_i_i_a3_8[6]_net_1 ), .Y(
        \data_out_2_15_i_i_11[6]_net_1 ));
    CFG1 #( .INIT(2'h1) )  un1_data_out8_126_set_RNO (.A(
        un1_data_out8_126_net_1), .Y(un1_data_out8_126_i));
    CFG3 #( .INIT(8'hF2) )  un1_data_out8_232 (.A(\mem_11_[5]_net_1 ), 
        .B(\mem_11__2_i_0_0_a2[2] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_232_i));
    CFG1 #( .INIT(2'h1) )  un1_data_out8_95_set_RNO (.A(
        un1_data_out8_95_net_1), .Y(un1_data_out8_95_i));
    CFG3 #( .INIT(8'h02) )  un1_data_out8_26 (.A(\mem_5_[7]_net_1 ), 
        .B(\mem_5__2_i_0_0_a2[0] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_26_net_1));
    SLE un1_data_out8_150_rs (.D(VCC_net_1), .CLK(
        un1_data_out8_86_net_1), .EN(VCC_net_1), .ALn(
        un1_data_out8_150_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(VCC_net_1), .Q(un1_data_out8_150_rs_net_1));
    SLE un1_data_out8_222_rs (.D(VCC_net_1), .CLK(
        un1_data_out8_118_net_1), .EN(VCC_net_1), .ALn(
        un1_data_out8_222_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(VCC_net_1), .Q(un1_data_out8_222_rs_net_1));
    SLE un1_data_out8_32_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_6__1_sqmuxa), .ALn(un1_data_out8_32_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_data_out8_32_set_net_1));
    CFG3 #( .INIT(8'hF8) )  un1_data_out8_49_set_RNI9PCL (.A(
        un1_data_out8_49_set_net_1), .B(un1_data_out8_132_rs_net_1), 
        .C(\mem_3_rs[4] ), .Y(\mem_3_[4]_net_1 ));
    CFG3 #( .INIT(8'hF8) )  un1_data_out8_67_set_RNIB1UO (.A(
        un1_data_out8_67_set_net_1), .B(un1_data_out8_141_rs_net_1), 
        .C(\mem_4_rs[5] ), .Y(\mem_4_[5]_net_1 ));
    CFG3 #( .INIT(8'hF8) )  un1_data_out8_52_set_RNIC2OE (.A(
        un1_data_out8_52_set_net_1), .B(un1_data_out8_227_rs_net_1), 
        .C(\mem_7_rs[4] ), .Y(\mem_7_[4]_net_1 ));
    CFG3 #( .INIT(8'h02) )  un1_data_out8_46 (.A(\mem_1_[7]_net_1 ), 
        .B(\mem_1__2_i_0_0_a2[0] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_46_net_1));
    CFG4 #( .INIT(16'h0004) )  \WRITE_GEN.mem_8__2_i_0_0_a2[2]  (.A(
        CoreAPB3_0_APBmslave4_PADDR[2]), .B(
        CoreAPB3_0_APBmslave4_PADDR[5]), .C(
        CoreAPB3_0_APBmslave4_PADDR[4]), .D(
        CoreAPB3_0_APBmslave4_PADDR[3]), .Y(mem_8__2_i_0_0_a2[2]));
    CFG1 #( .INIT(2'h1) )  un1_data_out8_91_set_RNO (.A(
        un1_data_out8_91_net_1), .Y(un1_data_out8_91_i));
    CFG1 #( .INIT(2'h1) )  un1_data_out8_29_set_RNO (.A(
        un1_data_out8_29_net_1), .Y(un1_data_out8_29_i));
    CFG2 #( .INIT(4'h8) )  mem_0__1_sqmuxa_0_a3_0_a3 (.A(
        mem_14__1_sqmuxa_0_a2_0_a3_0_a2_net_1), .B(
        mem_0__2_i_0_0_a2[0]), .Y(mem_0__1_sqmuxa));
    SLE un1_data_out8_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_4__1_sqmuxa), .ALn(un1_data_out8_i), .ADn(GND_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_data_out8_set_net_1));
    SLE un1_data_out8_49_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_3__1_sqmuxa), .ALn(un1_data_out8_49_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_data_out8_49_set_net_1));
    CFG4 #( .INIT(16'hECA0) )  \data_out_2_15_i_i_7[2]  (.A(
        \mem_8_[2]_net_1 ), .B(\mem_0_[2]_net_1 ), .C(
        mem_8__2_i_0_0_a2[2]), .D(mem_0__2_i_0_0_a2[0]), .Y(
        \data_out_2_15_i_i_7[2]_net_1 ));
    CFG1 #( .INIT(2'h1) )  un1_data_out8_120_set_RNO (.A(
        un1_data_out8_120_net_1), .Y(un1_data_out8_120_i));
    CFG1 #( .INIT(2'h1) )  un1_data_out8_102_set_RNO (.A(
        un1_data_out8_102_net_1), .Y(un1_data_out8_102_i));
    CFG3 #( .INIT(8'hF2) )  un1_data_out8_224 (.A(\mem_11_[1]_net_1 ), 
        .B(\mem_11__2_i_0_0_a2[2] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_224_i));
    SLE un1_data_out8_140_rs (.D(VCC_net_1), .CLK(
        un1_data_out8_65_net_1), .EN(VCC_net_1), .ALn(
        un1_data_out8_140_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(VCC_net_1), .Q(un1_data_out8_140_rs_net_1));
    CFG3 #( .INIT(8'h02) )  un1_data_out8_69 (.A(\mem_8_[5]_net_1 ), 
        .B(mem_8__2_i_0_0_a2[2]), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_69_net_1));
    CFG3 #( .INIT(8'hF2) )  un1_data_out8_209 (.A(\mem_13_[1]_net_1 ), 
        .B(\mem_13__2_i_0_0_a2[0] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_209_i));
    SLE \mem_6_[2]  (.D(CoreAPB3_0_APBmslave4_PWDATA[2]), .CLK(
        FCCC_0_GL1), .EN(mem_6__1_sqmuxa), .ALn(un1_data_out8_207_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_6_rs[2] ));
    SLE un1_data_out8_180_rs (.D(VCC_net_1), .CLK(
        un1_data_out8_100_net_1), .EN(VCC_net_1), .ALn(
        un1_data_out8_180_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(VCC_net_1), .Q(un1_data_out8_180_rs_net_1));
    CFG3 #( .INIT(8'hF8) )  un1_data_out8_79_set_RNIL2ET (.A(
        un1_data_out8_79_set_net_1), .B(un1_data_out8_204_rs_net_1), 
        .C(\mem_9_rs[7] ), .Y(\mem_9_[7]_net_1 ));
    CFG3 #( .INIT(8'h02) )  un1_data_out8_20 (.A(\mem_12_[4]_net_1 ), 
        .B(\mem_12__2_i_0_0_a2[0] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_20_net_1));
    CFG1 #( .INIT(2'h1) )  un1_data_out8_72_set_RNO (.A(
        un1_data_out8_72_net_1), .Y(un1_data_out8_72_i));
    SLE un1_data_out8_41_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_5__1_sqmuxa), .ALn(un1_data_out8_41_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_data_out8_41_set_net_1));
    CFG3 #( .INIT(8'hF8) )  un1_data_out8_143_rs_RNIPAKK (.A(
        un1_data_out8_8_set_net_1), .B(un1_data_out8_143_rs_net_1), .C(
        \mem_4_rs[6] ), .Y(\mem_4_[6]_net_1 ));
    CFG3 #( .INIT(8'hF8) )  un1_data_out8_154_rs_RNI0MFV (.A(
        un1_data_out8_13_set_net_1), .B(un1_data_out8_154_rs_net_1), 
        .C(\mem_1_rs[2] ), .Y(\mem_1_[2]_net_1 ));
    CFG3 #( .INIT(8'hF8) )  \mem_11__RNISSFV[0]  (.A(
        un1_data_out8_88_set_net_1), .B(un1_data_out8_182_rs_net_1), 
        .C(\mem_11_rs[0] ), .Y(\mem_11_[0]_net_1 ));
    CFG3 #( .INIT(8'hF2) )  un1_data_out8_254 (.A(\mem_15_[7]_net_1 ), 
        .B(\mem_15__2_i_0_0_a2[0] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_254_i));
    CFG3 #( .INIT(8'hF8) )  un1_data_out8_set_RNIU3D21 (.A(
        un1_data_out8_set_net_1), .B(un1_data_out8_136_rs_net_1), .C(
        \mem_4_rs[0] ), .Y(\mem_4_[0]_net_1 ));
    SLE \mem_7_[7]  (.D(CoreAPB3_0_APBmslave4_PWDATA[7]), .CLK(
        FCCC_0_GL1), .EN(mem_7__1_sqmuxa), .ALn(un1_data_out8_233_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_7_rs[7] ));
    SLE un1_data_out8_114_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_14__1_sqmuxa), .ALn(un1_data_out8_114_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_data_out8_114_set_net_1));
    CFG2 #( .INIT(4'h8) )  \data_out_2_15_i_i_a3_8[2]  (.A(
        \mem_3__2_i_0_0_a2[0] ), .B(\mem_3_[2]_net_1 ), .Y(
        \data_out_2_15_i_i_a3_8[2]_net_1 ));
    CFG1 #( .INIT(2'h1) )  un1_data_out8_10_set_RNO (.A(
        un1_data_out8_10_net_1), .Y(un1_data_out8_10_i));
    CFG3 #( .INIT(8'h02) )  un1_data_out8_40 (.A(\mem_1_[4]_net_1 ), 
        .B(\mem_1__2_i_0_0_a2[0] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_40_net_1));
    SLE un1_data_out8_251_rs (.D(VCC_net_1), .CLK(
        un1_data_out8_57_net_1), .EN(VCC_net_1), .ALn(
        un1_data_out8_251_i), .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(
        GND_net_1), .LAT(VCC_net_1), .Q(un1_data_out8_251_rs_net_1));
    SLE \mem_0_[2]  (.D(CoreAPB3_0_APBmslave4_PWDATA[2]), .CLK(
        FCCC_0_GL1), .EN(mem_0__1_sqmuxa), .ALn(un1_data_out8_145_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_0_rs[2] ));
    SLE un1_data_out8_124_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_7__1_sqmuxa), .ALn(un1_data_out8_124_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_data_out8_124_set_net_1));
    CFG1 #( .INIT(2'h1) )  un1_data_out8_113_set_RNO (.A(
        un1_data_out8_113_net_1), .Y(un1_data_out8_113_i));
    SLE \mem_3_[6]  (.D(CoreAPB3_0_APBmslave4_PWDATA[6]), .CLK(
        FCCC_0_GL1), .EN(mem_3__1_sqmuxa), .ALn(un1_data_out8_134_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_3_rs[6] ));
    SLE \mem_2_[7]  (.D(CoreAPB3_0_APBmslave4_PWDATA[7]), .CLK(
        FCCC_0_GL1), .EN(mem_2__1_sqmuxa), .ALn(un1_data_out8_167_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_2_rs[7] ));
    CFG4 #( .INIT(16'hECA0) )  \data_out_2_15_i_i_1[5]  (.A(
        \mem_14_[5]_net_1 ), .B(\mem_9_[5]_net_1 ), .C(
        \mem_14__2_i_0_0_a2[2] ), .D(\mem_9__2_i_0_0_a2[0] ), .Y(
        \data_out_2_15_i_i_1[5]_net_1 ));
    SLE \mem_7_[5]  (.D(CoreAPB3_0_APBmslave4_PWDATA[5]), .CLK(
        FCCC_0_GL1), .EN(mem_7__1_sqmuxa), .ALn(un1_data_out8_229_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_7_rs[5] ));
    CFG4 #( .INIT(16'h2000) )  \WRITE_GEN.mem_7__2_i_0_0_a2[1]  (.A(
        CoreAPB3_0_APBmslave4_PADDR[2]), .B(
        CoreAPB3_0_APBmslave4_PADDR[5]), .C(
        CoreAPB3_0_APBmslave4_PADDR[4]), .D(
        CoreAPB3_0_APBmslave4_PADDR[3]), .Y(\mem_7__2_i_0_0_a2[1] ));
    SLE un1_data_out8_19_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_12__1_sqmuxa), .ALn(un1_data_out8_19_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_data_out8_19_set_net_1));
    SLE un1_data_out8_104_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_13__1_sqmuxa), .ALn(un1_data_out8_104_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_data_out8_104_set_net_1));
    SLE un1_data_out8_20_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_12__1_sqmuxa), .ALn(un1_data_out8_20_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_data_out8_20_set_net_1));
    CFG1 #( .INIT(2'h1) )  un1_data_out8_18_set_RNO (.A(
        un1_data_out8_18_net_1), .Y(un1_data_out8_18_i));
    SLE un1_data_out8_80_set (.D(GND_net_1), .CLK(FCCC_0_GL1), .EN(
        mem_0__1_sqmuxa), .ALn(un1_data_out8_80_i), .ADn(GND_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        un1_data_out8_80_set_net_1));
    CFG3 #( .INIT(8'hF2) )  un1_data_out8_244 (.A(\mem_12_[4]_net_1 ), 
        .B(\mem_12__2_i_0_0_a2[0] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_244_i));
    SLE \mem_2_[5]  (.D(CoreAPB3_0_APBmslave4_PWDATA[5]), .CLK(
        FCCC_0_GL1), .EN(mem_2__1_sqmuxa), .ALn(un1_data_out8_165_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_2_rs[5] ));
    CFG1 #( .INIT(2'h1) )  un1_data_out8_80_set_RNO (.A(
        un1_data_out8_80_net_1), .Y(un1_data_out8_80_i));
    SLE \mem_4_[7]  (.D(CoreAPB3_0_APBmslave4_PWDATA[7]), .CLK(
        FCCC_0_GL1), .EN(mem_4__1_sqmuxa), .ALn(un1_data_out8_185_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_4_rs[7] ));
    CFG1 #( .INIT(2'h1) )  un1_data_out8_99_set_RNO (.A(
        un1_data_out8_99_net_1), .Y(un1_data_out8_99_i));
    CFG1 #( .INIT(2'h1) )  un1_data_out8_115_set_RNO (.A(
        un1_data_out8_115_net_1), .Y(un1_data_out8_115_i));
    SLE \mem_14_[3]  (.D(CoreAPB3_0_APBmslave4_PWDATA[3]), .CLK(
        FCCC_0_GL1), .EN(mem_14__1_sqmuxa), .ALn(un1_data_out8_219_i), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\mem_14_rs[3] ));
    CFG3 #( .INIT(8'h02) )  un1_data_out8_112 (.A(\mem_14_[0]_net_1 ), 
        .B(\mem_14__2_i_0_0_a2[2] ), .C(MSS_RESET_N_M2F_c), .Y(
        un1_data_out8_112_net_1));
    
endmodule


module reg_apb_wrp(
       PRDATA_0_iv_0_0_a2_1,
       CoreAPB3_0_APBmslave5_PRDATA,
       CoreAPB3_0_APBmslave4_PWDATA,
       CoreAPB3_0_APBmslave4_PADDR,
       mem_8__2_i_0_0_a2,
       mem_0__2_i_0_0_a2,
       CoreAPB3_0_APBmslave4_PWRITE,
       MSS_RESET_N_M2F_c,
       FCCC_0_GL1,
       CoreAPB3_0_APBmslave4_PENABLE
    );
input  [3:3] PRDATA_0_iv_0_0_a2_1;
output [7:0] CoreAPB3_0_APBmslave5_PRDATA;
input  [7:0] CoreAPB3_0_APBmslave4_PWDATA;
input  [5:2] CoreAPB3_0_APBmslave4_PADDR;
output [2:2] mem_8__2_i_0_0_a2;
output [0:0] mem_0__2_i_0_0_a2;
input  CoreAPB3_0_APBmslave4_PWRITE;
input  MSS_RESET_N_M2F_c;
input  FCCC_0_GL1;
input  CoreAPB3_0_APBmslave4_PENABLE;

    wire rd_enable, GND_net_1, VCC_net_1;
    
    reg16x8 reg16x8_0 (.CoreAPB3_0_APBmslave5_PRDATA({
        CoreAPB3_0_APBmslave5_PRDATA[7], 
        CoreAPB3_0_APBmslave5_PRDATA[6], 
        CoreAPB3_0_APBmslave5_PRDATA[5], 
        CoreAPB3_0_APBmslave5_PRDATA[4], 
        CoreAPB3_0_APBmslave5_PRDATA[3], 
        CoreAPB3_0_APBmslave5_PRDATA[2], 
        CoreAPB3_0_APBmslave5_PRDATA[1], 
        CoreAPB3_0_APBmslave5_PRDATA[0]}), 
        .CoreAPB3_0_APBmslave4_PWDATA({CoreAPB3_0_APBmslave4_PWDATA[7], 
        CoreAPB3_0_APBmslave4_PWDATA[6], 
        CoreAPB3_0_APBmslave4_PWDATA[5], 
        CoreAPB3_0_APBmslave4_PWDATA[4], 
        CoreAPB3_0_APBmslave4_PWDATA[3], 
        CoreAPB3_0_APBmslave4_PWDATA[2], 
        CoreAPB3_0_APBmslave4_PWDATA[1], 
        CoreAPB3_0_APBmslave4_PWDATA[0]}), 
        .CoreAPB3_0_APBmslave4_PADDR({CoreAPB3_0_APBmslave4_PADDR[5], 
        CoreAPB3_0_APBmslave4_PADDR[4], CoreAPB3_0_APBmslave4_PADDR[3], 
        CoreAPB3_0_APBmslave4_PADDR[2]}), .mem_8__2_i_0_0_a2({
        mem_8__2_i_0_0_a2[2]}), .mem_0__2_i_0_0_a2({
        mem_0__2_i_0_0_a2[0]}), .PRDATA_0_iv_0_0_a2_1({
        PRDATA_0_iv_0_0_a2_1[3]}), .MSS_RESET_N_M2F_c(
        MSS_RESET_N_M2F_c), .FCCC_0_GL1(FCCC_0_GL1), .rd_enable(
        rd_enable), .CoreAPB3_0_APBmslave4_PENABLE(
        CoreAPB3_0_APBmslave4_PENABLE), .CoreAPB3_0_APBmslave4_PWRITE(
        CoreAPB3_0_APBmslave4_PWRITE));
    VCC VCC (.Y(VCC_net_1));
    CFG2 #( .INIT(4'h2) )  rd_enable_0_a3_0_a3 (.A(
        PRDATA_0_iv_0_0_a2_1[3]), .B(CoreAPB3_0_APBmslave4_PWRITE), .Y(
        rd_enable));
    GND GND (.Y(GND_net_1));
    
endmodule


module CoreGPIO_Z3(
       GPIO_OUT_1_c,
       CoreAPB3_0_APBmslave4_PWDATA,
       mem_8__2_i_0_0_a2,
       PRDATA_0_iv_0_0_a2_2_4,
       MSS_RESET_N_M2F_c,
       FCCC_0_GL1,
       CoreAPB3_0_APBmslave4_PWRITE,
       CoreAPB3_0_APBmslave4_PENABLE
    );
output [7:0] GPIO_OUT_1_c;
input  [7:0] CoreAPB3_0_APBmslave4_PWDATA;
input  [2:2] mem_8__2_i_0_0_a2;
input  [3:3] PRDATA_0_iv_0_0_a2_2_4;
input  MSS_RESET_N_M2F_c;
input  FCCC_0_GL1;
input  CoreAPB3_0_APBmslave4_PWRITE;
input  CoreAPB3_0_APBmslave4_PENABLE;

    wire VCC_net_1, GPOUT_reg35, GND_net_1;
    
    SLE \xhdl1.GEN_BITS[4].APB_8.GPOUT_reg[4]  (.D(
        CoreAPB3_0_APBmslave4_PWDATA[4]), .CLK(FCCC_0_GL1), .EN(
        GPOUT_reg35), .ALn(MSS_RESET_N_M2F_c), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        GPIO_OUT_1_c[4]));
    SLE \xhdl1.GEN_BITS[1].APB_8.GPOUT_reg[1]  (.D(
        CoreAPB3_0_APBmslave4_PWDATA[1]), .CLK(FCCC_0_GL1), .EN(
        GPOUT_reg35), .ALn(MSS_RESET_N_M2F_c), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        GPIO_OUT_1_c[1]));
    SLE \xhdl1.GEN_BITS[5].APB_8.GPOUT_reg[5]  (.D(
        CoreAPB3_0_APBmslave4_PWDATA[5]), .CLK(FCCC_0_GL1), .EN(
        GPOUT_reg35), .ALn(MSS_RESET_N_M2F_c), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        GPIO_OUT_1_c[5]));
    GND GND (.Y(GND_net_1));
    VCC VCC (.Y(VCC_net_1));
    SLE \xhdl1.GEN_BITS[3].APB_8.GPOUT_reg[3]  (.D(
        CoreAPB3_0_APBmslave4_PWDATA[3]), .CLK(FCCC_0_GL1), .EN(
        GPOUT_reg35), .ALn(MSS_RESET_N_M2F_c), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        GPIO_OUT_1_c[3]));
    SLE \xhdl1.GEN_BITS[2].APB_8.GPOUT_reg[2]  (.D(
        CoreAPB3_0_APBmslave4_PWDATA[2]), .CLK(FCCC_0_GL1), .EN(
        GPOUT_reg35), .ALn(MSS_RESET_N_M2F_c), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        GPIO_OUT_1_c[2]));
    SLE \xhdl1.GEN_BITS[7].APB_8.GPOUT_reg[7]  (.D(
        CoreAPB3_0_APBmslave4_PWDATA[7]), .CLK(FCCC_0_GL1), .EN(
        GPOUT_reg35), .ALn(MSS_RESET_N_M2F_c), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        GPIO_OUT_1_c[7]));
    CFG4 #( .INIT(16'h8000) )  
        \xhdl1.GEN_BITS[0].APB_8.GPOUT_reg35_0_a3_0_a3  (.A(
        mem_8__2_i_0_0_a2[2]), .B(PRDATA_0_iv_0_0_a2_2_4[3]), .C(
        CoreAPB3_0_APBmslave4_PWRITE), .D(
        CoreAPB3_0_APBmslave4_PENABLE), .Y(GPOUT_reg35));
    SLE \xhdl1.GEN_BITS[6].APB_8.GPOUT_reg[6]  (.D(
        CoreAPB3_0_APBmslave4_PWDATA[6]), .CLK(FCCC_0_GL1), .EN(
        GPOUT_reg35), .ALn(MSS_RESET_N_M2F_c), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        GPIO_OUT_1_c[6]));
    SLE \xhdl1.GEN_BITS[0].APB_8.GPOUT_reg[0]  (.D(
        CoreAPB3_0_APBmslave4_PWDATA[0]), .CLK(FCCC_0_GL1), .EN(
        GPOUT_reg35), .ALn(MSS_RESET_N_M2F_c), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        GPIO_OUT_1_c[0]));
    
endmodule


module hello_regs_COREAPBLSRAM_0_lsram_512to35328x32_512s_32s(
       lsram_width32_PRDATA,
       CoreAPB3_0_APBmslave4_PADDR,
       CoreAPB3_0_APBmslave4_PWDATA,
       FCCC_0_GL1,
       MSS_RESET_N_M2F_c,
       wen
    );
output [31:0] lsram_width32_PRDATA;
input  [8:0] CoreAPB3_0_APBmslave4_PADDR;
input  [31:0] CoreAPB3_0_APBmslave4_PWDATA;
input  FCCC_0_GL1;
input  MSS_RESET_N_M2F_c;
input  wen;

    wire VCC_net_1, GND_net_1;
    
    RAM1K18 block0 (.A_DOUT({nc0, lsram_width32_PRDATA[15], 
        lsram_width32_PRDATA[14], lsram_width32_PRDATA[13], 
        lsram_width32_PRDATA[12], lsram_width32_PRDATA[11], 
        lsram_width32_PRDATA[10], lsram_width32_PRDATA[9], 
        lsram_width32_PRDATA[8], nc1, lsram_width32_PRDATA[7], 
        lsram_width32_PRDATA[6], lsram_width32_PRDATA[5], 
        lsram_width32_PRDATA[4], lsram_width32_PRDATA[3], 
        lsram_width32_PRDATA[2], lsram_width32_PRDATA[1], 
        lsram_width32_PRDATA[0]}), .B_DOUT({nc2, 
        lsram_width32_PRDATA[31], lsram_width32_PRDATA[30], 
        lsram_width32_PRDATA[29], lsram_width32_PRDATA[28], 
        lsram_width32_PRDATA[27], lsram_width32_PRDATA[26], 
        lsram_width32_PRDATA[25], lsram_width32_PRDATA[24], nc3, 
        lsram_width32_PRDATA[23], lsram_width32_PRDATA[22], 
        lsram_width32_PRDATA[21], lsram_width32_PRDATA[20], 
        lsram_width32_PRDATA[19], lsram_width32_PRDATA[18], 
        lsram_width32_PRDATA[17], lsram_width32_PRDATA[16]}), .BUSY(), 
        .A_CLK(FCCC_0_GL1), .A_DOUT_CLK(VCC_net_1), .A_ARST_N(
        MSS_RESET_N_M2F_c), .A_DOUT_EN(VCC_net_1), .A_BLK({VCC_net_1, 
        VCC_net_1, VCC_net_1}), .A_DOUT_ARST_N(VCC_net_1), 
        .A_DOUT_SRST_N(VCC_net_1), .A_DIN({GND_net_1, 
        CoreAPB3_0_APBmslave4_PWDATA[15], 
        CoreAPB3_0_APBmslave4_PWDATA[14], 
        CoreAPB3_0_APBmslave4_PWDATA[13], 
        CoreAPB3_0_APBmslave4_PWDATA[12], 
        CoreAPB3_0_APBmslave4_PWDATA[11], 
        CoreAPB3_0_APBmslave4_PWDATA[10], 
        CoreAPB3_0_APBmslave4_PWDATA[9], 
        CoreAPB3_0_APBmslave4_PWDATA[8], GND_net_1, 
        CoreAPB3_0_APBmslave4_PWDATA[7], 
        CoreAPB3_0_APBmslave4_PWDATA[6], 
        CoreAPB3_0_APBmslave4_PWDATA[5], 
        CoreAPB3_0_APBmslave4_PWDATA[4], 
        CoreAPB3_0_APBmslave4_PWDATA[3], 
        CoreAPB3_0_APBmslave4_PWDATA[2], 
        CoreAPB3_0_APBmslave4_PWDATA[1], 
        CoreAPB3_0_APBmslave4_PWDATA[0]}), .A_ADDR({
        CoreAPB3_0_APBmslave4_PADDR[8], CoreAPB3_0_APBmslave4_PADDR[7], 
        CoreAPB3_0_APBmslave4_PADDR[6], CoreAPB3_0_APBmslave4_PADDR[5], 
        CoreAPB3_0_APBmslave4_PADDR[4], CoreAPB3_0_APBmslave4_PADDR[3], 
        CoreAPB3_0_APBmslave4_PADDR[2], CoreAPB3_0_APBmslave4_PADDR[1], 
        CoreAPB3_0_APBmslave4_PADDR[0], GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1}), .A_WEN({wen, wen}), .B_CLK(
        FCCC_0_GL1), .B_DOUT_CLK(VCC_net_1), .B_ARST_N(
        MSS_RESET_N_M2F_c), .B_DOUT_EN(VCC_net_1), .B_BLK({VCC_net_1, 
        VCC_net_1, VCC_net_1}), .B_DOUT_ARST_N(VCC_net_1), 
        .B_DOUT_SRST_N(VCC_net_1), .B_DIN({GND_net_1, 
        CoreAPB3_0_APBmslave4_PWDATA[31], 
        CoreAPB3_0_APBmslave4_PWDATA[30], 
        CoreAPB3_0_APBmslave4_PWDATA[29], 
        CoreAPB3_0_APBmslave4_PWDATA[28], 
        CoreAPB3_0_APBmslave4_PWDATA[27], 
        CoreAPB3_0_APBmslave4_PWDATA[26], 
        CoreAPB3_0_APBmslave4_PWDATA[25], 
        CoreAPB3_0_APBmslave4_PWDATA[24], GND_net_1, 
        CoreAPB3_0_APBmslave4_PWDATA[23], 
        CoreAPB3_0_APBmslave4_PWDATA[22], 
        CoreAPB3_0_APBmslave4_PWDATA[21], 
        CoreAPB3_0_APBmslave4_PWDATA[20], 
        CoreAPB3_0_APBmslave4_PWDATA[19], 
        CoreAPB3_0_APBmslave4_PWDATA[18], 
        CoreAPB3_0_APBmslave4_PWDATA[17], 
        CoreAPB3_0_APBmslave4_PWDATA[16]}), .B_ADDR({
        CoreAPB3_0_APBmslave4_PADDR[8], CoreAPB3_0_APBmslave4_PADDR[7], 
        CoreAPB3_0_APBmslave4_PADDR[6], CoreAPB3_0_APBmslave4_PADDR[5], 
        CoreAPB3_0_APBmslave4_PADDR[4], CoreAPB3_0_APBmslave4_PADDR[3], 
        CoreAPB3_0_APBmslave4_PADDR[2], CoreAPB3_0_APBmslave4_PADDR[1], 
        CoreAPB3_0_APBmslave4_PADDR[0], GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1}), .B_WEN({wen, wen}), .A_EN(
        VCC_net_1), .A_DOUT_LAT(VCC_net_1), .A_WIDTH({VCC_net_1, 
        GND_net_1, VCC_net_1}), .A_WMODE(GND_net_1), .B_EN(VCC_net_1), 
        .B_DOUT_LAT(VCC_net_1), .B_WIDTH({VCC_net_1, GND_net_1, 
        VCC_net_1}), .B_WMODE(GND_net_1), .SII_LOCK(GND_net_1));
    VCC VCC (.Y(VCC_net_1));
    GND GND (.Y(GND_net_1));
    
endmodule


module hello_regs_COREAPBLSRAM_0_COREAPBLSRAM_Z2(
       PRDATA_reg,
       lsram_width32_PRDATA,
       hello_regs_MSS_0_FIC_0_APB_MASTER_PADDR,
       CoreAPB3_0_APBmslave4_PADDR,
       CoreAPB3_0_APBmslave4_PWDATA,
       MSS_RESET_N_M2F_c,
       FCCC_0_GL1,
       PRDATA4,
       CoreAPB3_0_APBmslave4_PREADY,
       CoreAPB3_0_APBmslave4_PWRITE,
       CoreAPB3_0_APBmslave4_PENABLE,
       N_928,
       hello_regs_MSS_0_FIC_0_APB_MASTER_PSELx
    );
output [31:0] PRDATA_reg;
output [31:0] lsram_width32_PRDATA;
input  [27:24] hello_regs_MSS_0_FIC_0_APB_MASTER_PADDR;
input  [8:0] CoreAPB3_0_APBmslave4_PADDR;
input  [31:0] CoreAPB3_0_APBmslave4_PWDATA;
input  MSS_RESET_N_M2F_c;
input  FCCC_0_GL1;
output PRDATA4;
output CoreAPB3_0_APBmslave4_PREADY;
input  CoreAPB3_0_APBmslave4_PWRITE;
input  CoreAPB3_0_APBmslave4_PENABLE;
output N_928;
input  hello_regs_MSS_0_FIC_0_APB_MASTER_PSELx;

    wire VCC_net_1, GND_net_1, PREADY_reg6_i_0, 
        PREADY_reg6_0_a3_0_a3_0_net_1, wen;
    
    SLE \PRDATA_reg[13]  (.D(lsram_width32_PRDATA[13]), .CLK(
        FCCC_0_GL1), .EN(PRDATA4), .ALn(MSS_RESET_N_M2F_c), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(PRDATA_reg[13]));
    hello_regs_COREAPBLSRAM_0_lsram_512to35328x32_512s_32s 
        \genblk1.genblk1.lsram_512to35328x32_block0  (
        .lsram_width32_PRDATA({lsram_width32_PRDATA[31], 
        lsram_width32_PRDATA[30], lsram_width32_PRDATA[29], 
        lsram_width32_PRDATA[28], lsram_width32_PRDATA[27], 
        lsram_width32_PRDATA[26], lsram_width32_PRDATA[25], 
        lsram_width32_PRDATA[24], lsram_width32_PRDATA[23], 
        lsram_width32_PRDATA[22], lsram_width32_PRDATA[21], 
        lsram_width32_PRDATA[20], lsram_width32_PRDATA[19], 
        lsram_width32_PRDATA[18], lsram_width32_PRDATA[17], 
        lsram_width32_PRDATA[16], lsram_width32_PRDATA[15], 
        lsram_width32_PRDATA[14], lsram_width32_PRDATA[13], 
        lsram_width32_PRDATA[12], lsram_width32_PRDATA[11], 
        lsram_width32_PRDATA[10], lsram_width32_PRDATA[9], 
        lsram_width32_PRDATA[8], lsram_width32_PRDATA[7], 
        lsram_width32_PRDATA[6], lsram_width32_PRDATA[5], 
        lsram_width32_PRDATA[4], lsram_width32_PRDATA[3], 
        lsram_width32_PRDATA[2], lsram_width32_PRDATA[1], 
        lsram_width32_PRDATA[0]}), .CoreAPB3_0_APBmslave4_PADDR({
        CoreAPB3_0_APBmslave4_PADDR[8], CoreAPB3_0_APBmslave4_PADDR[7], 
        CoreAPB3_0_APBmslave4_PADDR[6], CoreAPB3_0_APBmslave4_PADDR[5], 
        CoreAPB3_0_APBmslave4_PADDR[4], CoreAPB3_0_APBmslave4_PADDR[3], 
        CoreAPB3_0_APBmslave4_PADDR[2], CoreAPB3_0_APBmslave4_PADDR[1], 
        CoreAPB3_0_APBmslave4_PADDR[0]}), 
        .CoreAPB3_0_APBmslave4_PWDATA({
        CoreAPB3_0_APBmslave4_PWDATA[31], 
        CoreAPB3_0_APBmslave4_PWDATA[30], 
        CoreAPB3_0_APBmslave4_PWDATA[29], 
        CoreAPB3_0_APBmslave4_PWDATA[28], 
        CoreAPB3_0_APBmslave4_PWDATA[27], 
        CoreAPB3_0_APBmslave4_PWDATA[26], 
        CoreAPB3_0_APBmslave4_PWDATA[25], 
        CoreAPB3_0_APBmslave4_PWDATA[24], 
        CoreAPB3_0_APBmslave4_PWDATA[23], 
        CoreAPB3_0_APBmslave4_PWDATA[22], 
        CoreAPB3_0_APBmslave4_PWDATA[21], 
        CoreAPB3_0_APBmslave4_PWDATA[20], 
        CoreAPB3_0_APBmslave4_PWDATA[19], 
        CoreAPB3_0_APBmslave4_PWDATA[18], 
        CoreAPB3_0_APBmslave4_PWDATA[17], 
        CoreAPB3_0_APBmslave4_PWDATA[16], 
        CoreAPB3_0_APBmslave4_PWDATA[15], 
        CoreAPB3_0_APBmslave4_PWDATA[14], 
        CoreAPB3_0_APBmslave4_PWDATA[13], 
        CoreAPB3_0_APBmslave4_PWDATA[12], 
        CoreAPB3_0_APBmslave4_PWDATA[11], 
        CoreAPB3_0_APBmslave4_PWDATA[10], 
        CoreAPB3_0_APBmslave4_PWDATA[9], 
        CoreAPB3_0_APBmslave4_PWDATA[8], 
        CoreAPB3_0_APBmslave4_PWDATA[7], 
        CoreAPB3_0_APBmslave4_PWDATA[6], 
        CoreAPB3_0_APBmslave4_PWDATA[5], 
        CoreAPB3_0_APBmslave4_PWDATA[4], 
        CoreAPB3_0_APBmslave4_PWDATA[3], 
        CoreAPB3_0_APBmslave4_PWDATA[2], 
        CoreAPB3_0_APBmslave4_PWDATA[1], 
        CoreAPB3_0_APBmslave4_PWDATA[0]}), .FCCC_0_GL1(FCCC_0_GL1), 
        .MSS_RESET_N_M2F_c(MSS_RESET_N_M2F_c), .wen(wen));
    SLE \PRDATA_reg[26]  (.D(lsram_width32_PRDATA[26]), .CLK(
        FCCC_0_GL1), .EN(PRDATA4), .ALn(MSS_RESET_N_M2F_c), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(PRDATA_reg[26]));
    SLE \PRDATA_reg[6]  (.D(lsram_width32_PRDATA[6]), .CLK(FCCC_0_GL1), 
        .EN(PRDATA4), .ALn(MSS_RESET_N_M2F_c), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(PRDATA_reg[6]));
    SLE \PRDATA_reg[14]  (.D(lsram_width32_PRDATA[14]), .CLK(
        FCCC_0_GL1), .EN(PRDATA4), .ALn(MSS_RESET_N_M2F_c), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(PRDATA_reg[14]));
    CFG4 #( .INIT(16'h0004) )  PREADY_reg6_0_a3_0_a2_0 (.A(
        hello_regs_MSS_0_FIC_0_APB_MASTER_PADDR[25]), .B(
        hello_regs_MSS_0_FIC_0_APB_MASTER_PSELx), .C(
        hello_regs_MSS_0_FIC_0_APB_MASTER_PADDR[27]), .D(
        hello_regs_MSS_0_FIC_0_APB_MASTER_PADDR[24]), .Y(N_928));
    SLE \PRDATA_reg[17]  (.D(lsram_width32_PRDATA[17]), .CLK(
        FCCC_0_GL1), .EN(PRDATA4), .ALn(MSS_RESET_N_M2F_c), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(PRDATA_reg[17]));
    SLE \PRDATA_reg[15]  (.D(lsram_width32_PRDATA[15]), .CLK(
        FCCC_0_GL1), .EN(PRDATA4), .ALn(MSS_RESET_N_M2F_c), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(PRDATA_reg[15]));
    VCC VCC (.Y(VCC_net_1));
    SLE \PRDATA_reg[9]  (.D(lsram_width32_PRDATA[9]), .CLK(FCCC_0_GL1), 
        .EN(PRDATA4), .ALn(MSS_RESET_N_M2F_c), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(PRDATA_reg[9]));
    CFG2 #( .INIT(4'h4) )  PREADY_reg6_0_a3_0_a3_0 (.A(
        CoreAPB3_0_APBmslave4_PWRITE), .B(CoreAPB3_0_APBmslave4_PREADY)
        , .Y(PREADY_reg6_0_a3_0_a3_0_net_1));
    SLE \PRDATA_reg[10]  (.D(lsram_width32_PRDATA[10]), .CLK(
        FCCC_0_GL1), .EN(PRDATA4), .ALn(MSS_RESET_N_M2F_c), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(PRDATA_reg[10]));
    SLE \PRDATA_reg[23]  (.D(lsram_width32_PRDATA[23]), .CLK(
        FCCC_0_GL1), .EN(PRDATA4), .ALn(MSS_RESET_N_M2F_c), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(PRDATA_reg[23]));
    SLE \PRDATA_reg[4]  (.D(lsram_width32_PRDATA[4]), .CLK(FCCC_0_GL1), 
        .EN(PRDATA4), .ALn(MSS_RESET_N_M2F_c), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(PRDATA_reg[4]));
    GND GND (.Y(GND_net_1));
    SLE \PRDATA_reg[24]  (.D(lsram_width32_PRDATA[24]), .CLK(
        FCCC_0_GL1), .EN(PRDATA4), .ALn(MSS_RESET_N_M2F_c), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(PRDATA_reg[24]));
    SLE \PRDATA_reg[27]  (.D(lsram_width32_PRDATA[27]), .CLK(
        FCCC_0_GL1), .EN(PRDATA4), .ALn(MSS_RESET_N_M2F_c), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(PRDATA_reg[27]));
    SLE \PRDATA_reg[19]  (.D(lsram_width32_PRDATA[19]), .CLK(
        FCCC_0_GL1), .EN(PRDATA4), .ALn(MSS_RESET_N_M2F_c), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(PRDATA_reg[19]));
    SLE \PRDATA_reg[2]  (.D(lsram_width32_PRDATA[2]), .CLK(FCCC_0_GL1), 
        .EN(PRDATA4), .ALn(MSS_RESET_N_M2F_c), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(PRDATA_reg[2]));
    SLE \PRDATA_reg[25]  (.D(lsram_width32_PRDATA[25]), .CLK(
        FCCC_0_GL1), .EN(PRDATA4), .ALn(MSS_RESET_N_M2F_c), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(PRDATA_reg[25]));
    SLE \PRDATA_reg[3]  (.D(lsram_width32_PRDATA[3]), .CLK(FCCC_0_GL1), 
        .EN(PRDATA4), .ALn(MSS_RESET_N_M2F_c), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(PRDATA_reg[3]));
    SLE \PRDATA_reg[11]  (.D(lsram_width32_PRDATA[11]), .CLK(
        FCCC_0_GL1), .EN(PRDATA4), .ALn(MSS_RESET_N_M2F_c), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(PRDATA_reg[11]));
    SLE \PRDATA_reg[18]  (.D(lsram_width32_PRDATA[18]), .CLK(
        FCCC_0_GL1), .EN(PRDATA4), .ALn(MSS_RESET_N_M2F_c), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(PRDATA_reg[18]));
    SLE \PRDATA_reg[20]  (.D(lsram_width32_PRDATA[20]), .CLK(
        FCCC_0_GL1), .EN(PRDATA4), .ALn(MSS_RESET_N_M2F_c), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(PRDATA_reg[20]));
    SLE \PRDATA_reg[30]  (.D(lsram_width32_PRDATA[30]), .CLK(
        FCCC_0_GL1), .EN(PRDATA4), .ALn(MSS_RESET_N_M2F_c), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(PRDATA_reg[30]));
    SLE \PRDATA_reg[12]  (.D(lsram_width32_PRDATA[12]), .CLK(
        FCCC_0_GL1), .EN(PRDATA4), .ALn(MSS_RESET_N_M2F_c), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(PRDATA_reg[12]));
    CFG4 #( .INIT(16'hBFFF) )  PREADY_reg6_i (.A(
        CoreAPB3_0_APBmslave4_PENABLE), .B(
        hello_regs_MSS_0_FIC_0_APB_MASTER_PADDR[26]), .C(
        PREADY_reg6_0_a3_0_a3_0_net_1), .D(N_928), .Y(PREADY_reg6_i_0));
    SLE \PRDATA_reg[5]  (.D(lsram_width32_PRDATA[5]), .CLK(FCCC_0_GL1), 
        .EN(PRDATA4), .ALn(MSS_RESET_N_M2F_c), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(PRDATA_reg[5]));
    SLE \PRDATA_reg[1]  (.D(lsram_width32_PRDATA[1]), .CLK(FCCC_0_GL1), 
        .EN(PRDATA4), .ALn(MSS_RESET_N_M2F_c), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(PRDATA_reg[1]));
    SLE \PRDATA_reg[16]  (.D(lsram_width32_PRDATA[16]), .CLK(
        FCCC_0_GL1), .EN(PRDATA4), .ALn(MSS_RESET_N_M2F_c), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(PRDATA_reg[16]));
    SLE \PRDATA_reg[8]  (.D(lsram_width32_PRDATA[8]), .CLK(FCCC_0_GL1), 
        .EN(PRDATA4), .ALn(MSS_RESET_N_M2F_c), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(PRDATA_reg[8]));
    SLE \PRDATA_reg[29]  (.D(lsram_width32_PRDATA[29]), .CLK(
        FCCC_0_GL1), .EN(PRDATA4), .ALn(MSS_RESET_N_M2F_c), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(PRDATA_reg[29]));
    SLE \PRDATA_reg[0]  (.D(lsram_width32_PRDATA[0]), .CLK(FCCC_0_GL1), 
        .EN(PRDATA4), .ALn(MSS_RESET_N_M2F_c), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(PRDATA_reg[0]));
    SLE \PRDATA_reg[21]  (.D(lsram_width32_PRDATA[21]), .CLK(
        FCCC_0_GL1), .EN(PRDATA4), .ALn(MSS_RESET_N_M2F_c), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(PRDATA_reg[21]));
    SLE \PRDATA_reg[31]  (.D(lsram_width32_PRDATA[31]), .CLK(
        FCCC_0_GL1), .EN(PRDATA4), .ALn(MSS_RESET_N_M2F_c), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(PRDATA_reg[31]));
    SLE \PRDATA_reg[7]  (.D(lsram_width32_PRDATA[7]), .CLK(FCCC_0_GL1), 
        .EN(PRDATA4), .ALn(MSS_RESET_N_M2F_c), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(PRDATA_reg[7]));
    CFG4 #( .INIT(16'h8000) )  wen_0_a3_0_a3 (.A(
        CoreAPB3_0_APBmslave4_PWRITE), .B(
        CoreAPB3_0_APBmslave4_PENABLE), .C(
        hello_regs_MSS_0_FIC_0_APB_MASTER_PADDR[26]), .D(N_928), .Y(
        wen));
    SLE PREADY_reg (.D(PREADY_reg6_i_0), .CLK(FCCC_0_GL1), .EN(
        VCC_net_1), .ALn(MSS_RESET_N_M2F_c), .ADn(GND_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        CoreAPB3_0_APBmslave4_PREADY));
    SLE \PRDATA_reg[28]  (.D(lsram_width32_PRDATA[28]), .CLK(
        FCCC_0_GL1), .EN(PRDATA4), .ALn(MSS_RESET_N_M2F_c), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(PRDATA_reg[28]));
    CFG4 #( .INIT(16'h4000) )  PRDATA4_0_a2_0_a2 (.A(
        CoreAPB3_0_APBmslave4_PWRITE), .B(
        CoreAPB3_0_APBmslave4_PENABLE), .C(
        hello_regs_MSS_0_FIC_0_APB_MASTER_PADDR[26]), .D(N_928), .Y(
        PRDATA4));
    SLE \PRDATA_reg[22]  (.D(lsram_width32_PRDATA[22]), .CLK(
        FCCC_0_GL1), .EN(PRDATA4), .ALn(MSS_RESET_N_M2F_c), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(PRDATA_reg[22]));
    
endmodule


module hello_regs(
       GPIO_IN,
       GPIO_OUT_1,
       MMUART_0_RXD,
       MMUART_0_TXD,
       MSS_RESET_N_M2F
    );
input  [7:0] GPIO_IN;
output [7:0] GPIO_OUT_1;
input  MMUART_0_RXD;
output MMUART_0_TXD;
output MSS_RESET_N_M2F;

    wire GND_net_1, FCCC_0_GL1, \CoreAPB3_0_APBmslave4_PADDR[0] , 
        \CoreAPB3_0_APBmslave4_PADDR[1] , 
        \CoreAPB3_0_APBmslave4_PADDR[2] , 
        \CoreAPB3_0_APBmslave4_PADDR[3] , 
        \CoreAPB3_0_APBmslave4_PADDR[4] , 
        \CoreAPB3_0_APBmslave4_PADDR[5] , 
        \CoreAPB3_0_APBmslave4_PADDR[6] , 
        \CoreAPB3_0_APBmslave4_PADDR[7] , 
        \CoreAPB3_0_APBmslave4_PADDR[8] , 
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PADDR[9] , 
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PADDR[10] , 
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PADDR[11] , 
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PADDR[12] , 
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PADDR[13] , 
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PADDR[14] , 
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PADDR[15] , 
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PADDR[16] , 
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PADDR[17] , 
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PADDR[18] , 
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PADDR[19] , 
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PADDR[20] , 
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PADDR[21] , 
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PADDR[22] , 
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PADDR[23] , 
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PADDR[24] , 
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PADDR[25] , 
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PADDR[26] , 
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PADDR[27] , 
        CoreAPB3_0_APBmslave4_PWRITE, CoreAPB3_0_APBmslave4_PENABLE, 
        hello_regs_MSS_0_FIC_0_APB_MASTER_PSELx, 
        \CoreAPB3_0_APBmslave4_PWDATA[0] , 
        \CoreAPB3_0_APBmslave4_PWDATA[1] , 
        \CoreAPB3_0_APBmslave4_PWDATA[2] , 
        \CoreAPB3_0_APBmslave4_PWDATA[3] , 
        \CoreAPB3_0_APBmslave4_PWDATA[4] , 
        \CoreAPB3_0_APBmslave4_PWDATA[5] , 
        \CoreAPB3_0_APBmslave4_PWDATA[6] , 
        \CoreAPB3_0_APBmslave4_PWDATA[7] , 
        \CoreAPB3_0_APBmslave4_PWDATA[8] , 
        \CoreAPB3_0_APBmslave4_PWDATA[9] , 
        \CoreAPB3_0_APBmslave4_PWDATA[10] , 
        \CoreAPB3_0_APBmslave4_PWDATA[11] , 
        \CoreAPB3_0_APBmslave4_PWDATA[12] , 
        \CoreAPB3_0_APBmslave4_PWDATA[13] , 
        \CoreAPB3_0_APBmslave4_PWDATA[14] , 
        \CoreAPB3_0_APBmslave4_PWDATA[15] , 
        \CoreAPB3_0_APBmslave4_PWDATA[16] , 
        \CoreAPB3_0_APBmslave4_PWDATA[17] , 
        \CoreAPB3_0_APBmslave4_PWDATA[18] , 
        \CoreAPB3_0_APBmslave4_PWDATA[19] , 
        \CoreAPB3_0_APBmslave4_PWDATA[20] , 
        \CoreAPB3_0_APBmslave4_PWDATA[21] , 
        \CoreAPB3_0_APBmslave4_PWDATA[22] , 
        \CoreAPB3_0_APBmslave4_PWDATA[23] , 
        \CoreAPB3_0_APBmslave4_PWDATA[24] , 
        \CoreAPB3_0_APBmslave4_PWDATA[25] , 
        \CoreAPB3_0_APBmslave4_PWDATA[26] , 
        \CoreAPB3_0_APBmslave4_PWDATA[27] , 
        \CoreAPB3_0_APBmslave4_PWDATA[28] , 
        \CoreAPB3_0_APBmslave4_PWDATA[29] , 
        \CoreAPB3_0_APBmslave4_PWDATA[30] , 
        \CoreAPB3_0_APBmslave4_PWDATA[31] , 
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[0] , 
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[1] , 
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[2] , 
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[3] , 
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[4] , 
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[5] , 
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[6] , 
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[7] , 
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[8] , 
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[9] , 
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[10] , 
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[11] , 
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[12] , 
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[13] , 
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[14] , 
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[15] , 
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[16] , 
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[17] , 
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[18] , 
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[19] , 
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[20] , 
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[21] , 
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[22] , 
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[23] , 
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[24] , 
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[25] , 
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[26] , 
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[27] , 
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[28] , 
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[29] , 
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[30] , 
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[31] , 
        \CoreAPB3_0_APBmslave5_PRDATA[0] , 
        \CoreAPB3_0_APBmslave5_PRDATA[1] , 
        \CoreAPB3_0_APBmslave5_PRDATA[2] , 
        \CoreAPB3_0_APBmslave5_PRDATA[3] , 
        \CoreAPB3_0_APBmslave5_PRDATA[4] , 
        \CoreAPB3_0_APBmslave5_PRDATA[5] , 
        \CoreAPB3_0_APBmslave5_PRDATA[6] , 
        \CoreAPB3_0_APBmslave5_PRDATA[7] , 
        CoreAPB3_0_APBmslave4_PREADY, 
        OSC_0_RCOSC_25_50MHZ_CCC_OUT_RCOSC_25_50MHZ_CCC, FCCC_0_LOCK, 
        VCC_net_1, \COREAPBLSRAM_0.lsram_width32_PRDATA[0] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[1] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[2] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[3] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[4] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[5] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[6] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[7] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[8] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[9] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[10] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[11] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[12] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[13] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[14] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[15] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[16] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[17] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[18] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[19] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[20] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[21] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[22] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[23] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[24] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[25] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[26] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[27] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[28] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[29] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[30] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[31] , 
        \COREAPBLSRAM_0.PRDATA4 , \COREAPBLSRAM_0.PRDATA_reg[0] , 
        \COREAPBLSRAM_0.PRDATA_reg[1] , \COREAPBLSRAM_0.PRDATA_reg[2] , 
        \COREAPBLSRAM_0.PRDATA_reg[3] , \COREAPBLSRAM_0.PRDATA_reg[4] , 
        \COREAPBLSRAM_0.PRDATA_reg[5] , \COREAPBLSRAM_0.PRDATA_reg[6] , 
        \COREAPBLSRAM_0.PRDATA_reg[7] , \COREAPBLSRAM_0.PRDATA_reg[8] , 
        \COREAPBLSRAM_0.PRDATA_reg[9] , 
        \COREAPBLSRAM_0.PRDATA_reg[10] , 
        \COREAPBLSRAM_0.PRDATA_reg[11] , 
        \COREAPBLSRAM_0.PRDATA_reg[12] , 
        \COREAPBLSRAM_0.PRDATA_reg[13] , 
        \COREAPBLSRAM_0.PRDATA_reg[14] , 
        \COREAPBLSRAM_0.PRDATA_reg[15] , 
        \COREAPBLSRAM_0.PRDATA_reg[16] , 
        \COREAPBLSRAM_0.PRDATA_reg[17] , 
        \COREAPBLSRAM_0.PRDATA_reg[18] , 
        \COREAPBLSRAM_0.PRDATA_reg[19] , 
        \COREAPBLSRAM_0.PRDATA_reg[20] , 
        \COREAPBLSRAM_0.PRDATA_reg[21] , 
        \COREAPBLSRAM_0.PRDATA_reg[22] , 
        \COREAPBLSRAM_0.PRDATA_reg[23] , 
        \COREAPBLSRAM_0.PRDATA_reg[24] , 
        \COREAPBLSRAM_0.PRDATA_reg[25] , 
        \COREAPBLSRAM_0.PRDATA_reg[26] , 
        \COREAPBLSRAM_0.PRDATA_reg[27] , 
        \COREAPBLSRAM_0.PRDATA_reg[28] , 
        \COREAPBLSRAM_0.PRDATA_reg[29] , 
        \COREAPBLSRAM_0.PRDATA_reg[30] , 
        \COREAPBLSRAM_0.PRDATA_reg[31] , N_928, 
        \WRITE_GEN.mem_0__2_i_0_0_a2[0] , \PRDATA_0_iv_0_0_a2_1[3] , 
        \WRITE_GEN.mem_8__2_i_0_0_a2[2] , \GPIO_OUT_1_c[0] , 
        \GPIO_OUT_1_c[1] , \GPIO_OUT_1_c[2] , \GPIO_OUT_1_c[3] , 
        \GPIO_OUT_1_c[4] , \GPIO_OUT_1_c[5] , \GPIO_OUT_1_c[6] , 
        \GPIO_OUT_1_c[7] , MSS_RESET_N_M2F_c, 
        \CoreAPB3_0.u_mux_p_to_b3.PRDATA_0_iv_0_0_a2_2_4[3] , 
        N_676_i_0;
    
    CoreAPB3_Z1 CoreAPB3_0 (.PRDATA_0_iv_0_0_a2_1({
        \PRDATA_0_iv_0_0_a2_1[3] }), 
        .hello_regs_MSS_0_FIC_0_APB_MASTER_PADDR({
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PADDR[27] , 
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PADDR[26] , 
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PADDR[25] , 
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PADDR[24] , 
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PADDR[23] , 
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PADDR[22] , 
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PADDR[21] , 
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PADDR[20] , 
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PADDR[19] , 
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PADDR[18] , 
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PADDR[17] , 
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PADDR[16] , 
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PADDR[15] , 
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PADDR[14] , 
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PADDR[13] , 
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PADDR[12] , 
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PADDR[11] , 
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PADDR[10] , 
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PADDR[9] }), 
        .mem_8__2_i_0_0_a2({\WRITE_GEN.mem_8__2_i_0_0_a2[2] }), 
        .mem_0__2_i_0_0_a2({\WRITE_GEN.mem_0__2_i_0_0_a2[0] }), 
        .PRDATA_0_iv_0_0_a2_2_4({
        \CoreAPB3_0.u_mux_p_to_b3.PRDATA_0_iv_0_0_a2_2_4[3] }), 
        .CoreAPB3_0_APBmslave5_PRDATA({
        \CoreAPB3_0_APBmslave5_PRDATA[7] , 
        \CoreAPB3_0_APBmslave5_PRDATA[6] , 
        \CoreAPB3_0_APBmslave5_PRDATA[5] , 
        \CoreAPB3_0_APBmslave5_PRDATA[4] , 
        \CoreAPB3_0_APBmslave5_PRDATA[3] , 
        \CoreAPB3_0_APBmslave5_PRDATA[2] , 
        \CoreAPB3_0_APBmslave5_PRDATA[1] , 
        \CoreAPB3_0_APBmslave5_PRDATA[0] }), .PRDATA_reg({
        \COREAPBLSRAM_0.PRDATA_reg[31] , 
        \COREAPBLSRAM_0.PRDATA_reg[30] , 
        \COREAPBLSRAM_0.PRDATA_reg[29] , 
        \COREAPBLSRAM_0.PRDATA_reg[28] , 
        \COREAPBLSRAM_0.PRDATA_reg[27] , 
        \COREAPBLSRAM_0.PRDATA_reg[26] , 
        \COREAPBLSRAM_0.PRDATA_reg[25] , 
        \COREAPBLSRAM_0.PRDATA_reg[24] , 
        \COREAPBLSRAM_0.PRDATA_reg[23] , 
        \COREAPBLSRAM_0.PRDATA_reg[22] , 
        \COREAPBLSRAM_0.PRDATA_reg[21] , 
        \COREAPBLSRAM_0.PRDATA_reg[20] , 
        \COREAPBLSRAM_0.PRDATA_reg[19] , 
        \COREAPBLSRAM_0.PRDATA_reg[18] , 
        \COREAPBLSRAM_0.PRDATA_reg[17] , 
        \COREAPBLSRAM_0.PRDATA_reg[16] , 
        \COREAPBLSRAM_0.PRDATA_reg[15] , 
        \COREAPBLSRAM_0.PRDATA_reg[14] , 
        \COREAPBLSRAM_0.PRDATA_reg[13] , 
        \COREAPBLSRAM_0.PRDATA_reg[12] , 
        \COREAPBLSRAM_0.PRDATA_reg[11] , 
        \COREAPBLSRAM_0.PRDATA_reg[10] , 
        \COREAPBLSRAM_0.PRDATA_reg[9] , \COREAPBLSRAM_0.PRDATA_reg[8] , 
        \COREAPBLSRAM_0.PRDATA_reg[7] , \COREAPBLSRAM_0.PRDATA_reg[6] , 
        \COREAPBLSRAM_0.PRDATA_reg[5] , \COREAPBLSRAM_0.PRDATA_reg[4] , 
        \COREAPBLSRAM_0.PRDATA_reg[3] , \COREAPBLSRAM_0.PRDATA_reg[2] , 
        \COREAPBLSRAM_0.PRDATA_reg[1] , \COREAPBLSRAM_0.PRDATA_reg[0] })
        , .lsram_width32_PRDATA({
        \COREAPBLSRAM_0.lsram_width32_PRDATA[31] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[30] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[29] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[28] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[27] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[26] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[25] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[24] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[23] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[22] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[21] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[20] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[19] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[18] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[17] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[16] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[15] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[14] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[13] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[12] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[11] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[10] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[9] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[8] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[7] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[6] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[5] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[4] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[3] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[2] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[1] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[0] }), .GPIO_OUT_1_c({
        \GPIO_OUT_1_c[7] , \GPIO_OUT_1_c[6] , \GPIO_OUT_1_c[5] , 
        \GPIO_OUT_1_c[4] , \GPIO_OUT_1_c[3] , \GPIO_OUT_1_c[2] , 
        \GPIO_OUT_1_c[1] , \GPIO_OUT_1_c[0] }), 
        .hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA({
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[31] , 
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[30] , 
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[29] , 
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[28] , 
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[27] , 
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[26] , 
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[25] , 
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[24] , 
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[23] , 
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[22] , 
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[21] , 
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[20] , 
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[19] , 
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[18] , 
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[17] , 
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[16] , 
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[15] , 
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[14] , 
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[13] , 
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[12] , 
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[11] , 
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[10] , 
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[9] , 
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[8] , 
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[7] , 
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[6] , 
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[5] , 
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[4] , 
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[3] , 
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[2] , 
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[1] , 
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[0] }), 
        .CoreAPB3_0_APBmslave4_PWDATA({
        \CoreAPB3_0_APBmslave4_PWDATA[31] , 
        \CoreAPB3_0_APBmslave4_PWDATA[30] , 
        \CoreAPB3_0_APBmslave4_PWDATA[29] , 
        \CoreAPB3_0_APBmslave4_PWDATA[28] , 
        \CoreAPB3_0_APBmslave4_PWDATA[27] , 
        \CoreAPB3_0_APBmslave4_PWDATA[26] , 
        \CoreAPB3_0_APBmslave4_PWDATA[25] , 
        \CoreAPB3_0_APBmslave4_PWDATA[24] , 
        \CoreAPB3_0_APBmslave4_PWDATA[23] , 
        \CoreAPB3_0_APBmslave4_PWDATA[22] , 
        \CoreAPB3_0_APBmslave4_PWDATA[21] , 
        \CoreAPB3_0_APBmslave4_PWDATA[20] , 
        \CoreAPB3_0_APBmslave4_PWDATA[19] , 
        \CoreAPB3_0_APBmslave4_PWDATA[18] , 
        \CoreAPB3_0_APBmslave4_PWDATA[17] , 
        \CoreAPB3_0_APBmslave4_PWDATA[16] , 
        \CoreAPB3_0_APBmslave4_PWDATA[15] , 
        \CoreAPB3_0_APBmslave4_PWDATA[14] , 
        \CoreAPB3_0_APBmslave4_PWDATA[13] , 
        \CoreAPB3_0_APBmslave4_PWDATA[12] , 
        \CoreAPB3_0_APBmslave4_PWDATA[11] , 
        \CoreAPB3_0_APBmslave4_PWDATA[10] , 
        \CoreAPB3_0_APBmslave4_PWDATA[9] , 
        \CoreAPB3_0_APBmslave4_PWDATA[8] , 
        \CoreAPB3_0_APBmslave4_PWDATA[7] , 
        \CoreAPB3_0_APBmslave4_PWDATA[6] , 
        \CoreAPB3_0_APBmslave4_PWDATA[5] , 
        \CoreAPB3_0_APBmslave4_PWDATA[4] , 
        \CoreAPB3_0_APBmslave4_PWDATA[3] , 
        \CoreAPB3_0_APBmslave4_PWDATA[2] , 
        \CoreAPB3_0_APBmslave4_PWDATA[1] , 
        \CoreAPB3_0_APBmslave4_PWDATA[0] }), 
        .CoreAPB3_0_APBmslave4_PADDR_8(
        \CoreAPB3_0_APBmslave4_PADDR[8] ), 
        .CoreAPB3_0_APBmslave4_PADDR_7(
        \CoreAPB3_0_APBmslave4_PADDR[7] ), 
        .CoreAPB3_0_APBmslave4_PADDR_0(
        \CoreAPB3_0_APBmslave4_PADDR[0] ), 
        .CoreAPB3_0_APBmslave4_PADDR_6(
        \CoreAPB3_0_APBmslave4_PADDR[6] ), 
        .CoreAPB3_0_APBmslave4_PADDR_1(
        \CoreAPB3_0_APBmslave4_PADDR[1] ), 
        .hello_regs_MSS_0_FIC_0_APB_MASTER_PSELx(
        hello_regs_MSS_0_FIC_0_APB_MASTER_PSELx), .N_928(N_928), 
        .CoreAPB3_0_APBmslave4_PWRITE(CoreAPB3_0_APBmslave4_PWRITE), 
        .CoreAPB3_0_APBmslave4_PENABLE(CoreAPB3_0_APBmslave4_PENABLE), 
        .PRDATA4(\COREAPBLSRAM_0.PRDATA4 ), 
        .CoreAPB3_0_APBmslave4_PREADY(CoreAPB3_0_APBmslave4_PREADY), 
        .N_676_i_0(N_676_i_0), .MSS_RESET_N_M2F_c(MSS_RESET_N_M2F_c), 
        .FCCC_0_GL1(FCCC_0_GL1));
    OUTBUF \GPIO_OUT_1_obuf[7]  (.D(\GPIO_OUT_1_c[7] ), .PAD(
        GPIO_OUT_1[7]));
    OUTBUF \GPIO_OUT_1_obuf[1]  (.D(\GPIO_OUT_1_c[1] ), .PAD(
        GPIO_OUT_1[1]));
    GND GND (.Y(GND_net_1));
    hello_regs_OSC_0_OSC OSC_0 (
        .OSC_0_RCOSC_25_50MHZ_CCC_OUT_RCOSC_25_50MHZ_CCC(
        OSC_0_RCOSC_25_50MHZ_CCC_OUT_RCOSC_25_50MHZ_CCC));
    OUTBUF MSS_RESET_N_M2F_obuf (.D(MSS_RESET_N_M2F_c), .PAD(
        MSS_RESET_N_M2F));
    OUTBUF \GPIO_OUT_1_obuf[3]  (.D(\GPIO_OUT_1_c[3] ), .PAD(
        GPIO_OUT_1[3]));
    OUTBUF \GPIO_OUT_1_obuf[4]  (.D(\GPIO_OUT_1_c[4] ), .PAD(
        GPIO_OUT_1[4]));
    hello_regs_MSS hello_regs_MSS_0 (.CoreAPB3_0_APBmslave4_PADDR({
        \CoreAPB3_0_APBmslave4_PADDR[8] , 
        \CoreAPB3_0_APBmslave4_PADDR[7] , 
        \CoreAPB3_0_APBmslave4_PADDR[6] , 
        \CoreAPB3_0_APBmslave4_PADDR[5] , 
        \CoreAPB3_0_APBmslave4_PADDR[4] , 
        \CoreAPB3_0_APBmslave4_PADDR[3] , 
        \CoreAPB3_0_APBmslave4_PADDR[2] , 
        \CoreAPB3_0_APBmslave4_PADDR[1] , 
        \CoreAPB3_0_APBmslave4_PADDR[0] }), 
        .hello_regs_MSS_0_FIC_0_APB_MASTER_PADDR({
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PADDR[27] , 
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PADDR[26] , 
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PADDR[25] , 
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PADDR[24] , 
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PADDR[23] , 
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PADDR[22] , 
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PADDR[21] , 
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PADDR[20] , 
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PADDR[19] , 
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PADDR[18] , 
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PADDR[17] , 
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PADDR[16] , 
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PADDR[15] , 
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PADDR[14] , 
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PADDR[13] , 
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PADDR[12] , 
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PADDR[11] , 
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PADDR[10] , 
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PADDR[9] }), 
        .CoreAPB3_0_APBmslave4_PWDATA({
        \CoreAPB3_0_APBmslave4_PWDATA[31] , 
        \CoreAPB3_0_APBmslave4_PWDATA[30] , 
        \CoreAPB3_0_APBmslave4_PWDATA[29] , 
        \CoreAPB3_0_APBmslave4_PWDATA[28] , 
        \CoreAPB3_0_APBmslave4_PWDATA[27] , 
        \CoreAPB3_0_APBmslave4_PWDATA[26] , 
        \CoreAPB3_0_APBmslave4_PWDATA[25] , 
        \CoreAPB3_0_APBmslave4_PWDATA[24] , 
        \CoreAPB3_0_APBmslave4_PWDATA[23] , 
        \CoreAPB3_0_APBmslave4_PWDATA[22] , 
        \CoreAPB3_0_APBmslave4_PWDATA[21] , 
        \CoreAPB3_0_APBmslave4_PWDATA[20] , 
        \CoreAPB3_0_APBmslave4_PWDATA[19] , 
        \CoreAPB3_0_APBmslave4_PWDATA[18] , 
        \CoreAPB3_0_APBmslave4_PWDATA[17] , 
        \CoreAPB3_0_APBmslave4_PWDATA[16] , 
        \CoreAPB3_0_APBmslave4_PWDATA[15] , 
        \CoreAPB3_0_APBmslave4_PWDATA[14] , 
        \CoreAPB3_0_APBmslave4_PWDATA[13] , 
        \CoreAPB3_0_APBmslave4_PWDATA[12] , 
        \CoreAPB3_0_APBmslave4_PWDATA[11] , 
        \CoreAPB3_0_APBmslave4_PWDATA[10] , 
        \CoreAPB3_0_APBmslave4_PWDATA[9] , 
        \CoreAPB3_0_APBmslave4_PWDATA[8] , 
        \CoreAPB3_0_APBmslave4_PWDATA[7] , 
        \CoreAPB3_0_APBmslave4_PWDATA[6] , 
        \CoreAPB3_0_APBmslave4_PWDATA[5] , 
        \CoreAPB3_0_APBmslave4_PWDATA[4] , 
        \CoreAPB3_0_APBmslave4_PWDATA[3] , 
        \CoreAPB3_0_APBmslave4_PWDATA[2] , 
        \CoreAPB3_0_APBmslave4_PWDATA[1] , 
        \CoreAPB3_0_APBmslave4_PWDATA[0] }), 
        .hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA({
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[31] , 
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[30] , 
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[29] , 
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[28] , 
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[27] , 
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[26] , 
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[25] , 
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[24] , 
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[23] , 
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[22] , 
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[21] , 
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[20] , 
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[19] , 
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[18] , 
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[17] , 
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[16] , 
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[15] , 
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[14] , 
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[13] , 
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[12] , 
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[11] , 
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[10] , 
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[9] , 
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[8] , 
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[7] , 
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[6] , 
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[5] , 
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[4] , 
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[3] , 
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[2] , 
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[1] , 
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PRDATA[0] }), 
        .MSS_RESET_N_M2F_c(MSS_RESET_N_M2F_c), .MMUART_0_TXD(
        MMUART_0_TXD), .MMUART_0_RXD(MMUART_0_RXD), 
        .CoreAPB3_0_APBmslave4_PENABLE(CoreAPB3_0_APBmslave4_PENABLE), 
        .hello_regs_MSS_0_FIC_0_APB_MASTER_PSELx(
        hello_regs_MSS_0_FIC_0_APB_MASTER_PSELx), 
        .CoreAPB3_0_APBmslave4_PWRITE(CoreAPB3_0_APBmslave4_PWRITE), 
        .N_676_i_0(N_676_i_0), .FCCC_0_LOCK(FCCC_0_LOCK), .FCCC_0_GL1(
        FCCC_0_GL1));
    hello_regs_FCCC_0_FCCC FCCC_0 (.FCCC_0_GL1(FCCC_0_GL1), 
        .FCCC_0_LOCK(FCCC_0_LOCK), 
        .OSC_0_RCOSC_25_50MHZ_CCC_OUT_RCOSC_25_50MHZ_CCC(
        OSC_0_RCOSC_25_50MHZ_CCC_OUT_RCOSC_25_50MHZ_CCC));
    reg_apb_wrp reg_apb_wrp_0 (.PRDATA_0_iv_0_0_a2_1({
        \PRDATA_0_iv_0_0_a2_1[3] }), .CoreAPB3_0_APBmslave5_PRDATA({
        \CoreAPB3_0_APBmslave5_PRDATA[7] , 
        \CoreAPB3_0_APBmslave5_PRDATA[6] , 
        \CoreAPB3_0_APBmslave5_PRDATA[5] , 
        \CoreAPB3_0_APBmslave5_PRDATA[4] , 
        \CoreAPB3_0_APBmslave5_PRDATA[3] , 
        \CoreAPB3_0_APBmslave5_PRDATA[2] , 
        \CoreAPB3_0_APBmslave5_PRDATA[1] , 
        \CoreAPB3_0_APBmslave5_PRDATA[0] }), 
        .CoreAPB3_0_APBmslave4_PWDATA({
        \CoreAPB3_0_APBmslave4_PWDATA[7] , 
        \CoreAPB3_0_APBmslave4_PWDATA[6] , 
        \CoreAPB3_0_APBmslave4_PWDATA[5] , 
        \CoreAPB3_0_APBmslave4_PWDATA[4] , 
        \CoreAPB3_0_APBmslave4_PWDATA[3] , 
        \CoreAPB3_0_APBmslave4_PWDATA[2] , 
        \CoreAPB3_0_APBmslave4_PWDATA[1] , 
        \CoreAPB3_0_APBmslave4_PWDATA[0] }), 
        .CoreAPB3_0_APBmslave4_PADDR({\CoreAPB3_0_APBmslave4_PADDR[5] , 
        \CoreAPB3_0_APBmslave4_PADDR[4] , 
        \CoreAPB3_0_APBmslave4_PADDR[3] , 
        \CoreAPB3_0_APBmslave4_PADDR[2] }), .mem_8__2_i_0_0_a2({
        \WRITE_GEN.mem_8__2_i_0_0_a2[2] }), .mem_0__2_i_0_0_a2({
        \WRITE_GEN.mem_0__2_i_0_0_a2[0] }), 
        .CoreAPB3_0_APBmslave4_PWRITE(CoreAPB3_0_APBmslave4_PWRITE), 
        .MSS_RESET_N_M2F_c(MSS_RESET_N_M2F_c), .FCCC_0_GL1(FCCC_0_GL1), 
        .CoreAPB3_0_APBmslave4_PENABLE(CoreAPB3_0_APBmslave4_PENABLE));
    VCC VCC (.Y(VCC_net_1));
    OUTBUF \GPIO_OUT_1_obuf[0]  (.D(\GPIO_OUT_1_c[0] ), .PAD(
        GPIO_OUT_1[0]));
    OUTBUF \GPIO_OUT_1_obuf[5]  (.D(\GPIO_OUT_1_c[5] ), .PAD(
        GPIO_OUT_1[5]));
    OUTBUF \GPIO_OUT_1_obuf[2]  (.D(\GPIO_OUT_1_c[2] ), .PAD(
        GPIO_OUT_1[2]));
    CoreGPIO_Z3 CoreGPIO_0 (.GPIO_OUT_1_c({\GPIO_OUT_1_c[7] , 
        \GPIO_OUT_1_c[6] , \GPIO_OUT_1_c[5] , \GPIO_OUT_1_c[4] , 
        \GPIO_OUT_1_c[3] , \GPIO_OUT_1_c[2] , \GPIO_OUT_1_c[1] , 
        \GPIO_OUT_1_c[0] }), .CoreAPB3_0_APBmslave4_PWDATA({
        \CoreAPB3_0_APBmslave4_PWDATA[7] , 
        \CoreAPB3_0_APBmslave4_PWDATA[6] , 
        \CoreAPB3_0_APBmslave4_PWDATA[5] , 
        \CoreAPB3_0_APBmslave4_PWDATA[4] , 
        \CoreAPB3_0_APBmslave4_PWDATA[3] , 
        \CoreAPB3_0_APBmslave4_PWDATA[2] , 
        \CoreAPB3_0_APBmslave4_PWDATA[1] , 
        \CoreAPB3_0_APBmslave4_PWDATA[0] }), .mem_8__2_i_0_0_a2({
        \WRITE_GEN.mem_8__2_i_0_0_a2[2] }), .PRDATA_0_iv_0_0_a2_2_4({
        \CoreAPB3_0.u_mux_p_to_b3.PRDATA_0_iv_0_0_a2_2_4[3] }), 
        .MSS_RESET_N_M2F_c(MSS_RESET_N_M2F_c), .FCCC_0_GL1(FCCC_0_GL1), 
        .CoreAPB3_0_APBmslave4_PWRITE(CoreAPB3_0_APBmslave4_PWRITE), 
        .CoreAPB3_0_APBmslave4_PENABLE(CoreAPB3_0_APBmslave4_PENABLE));
    OUTBUF \GPIO_OUT_1_obuf[6]  (.D(\GPIO_OUT_1_c[6] ), .PAD(
        GPIO_OUT_1[6]));
    hello_regs_COREAPBLSRAM_0_COREAPBLSRAM_Z2 COREAPBLSRAM_0 (
        .PRDATA_reg({\COREAPBLSRAM_0.PRDATA_reg[31] , 
        \COREAPBLSRAM_0.PRDATA_reg[30] , 
        \COREAPBLSRAM_0.PRDATA_reg[29] , 
        \COREAPBLSRAM_0.PRDATA_reg[28] , 
        \COREAPBLSRAM_0.PRDATA_reg[27] , 
        \COREAPBLSRAM_0.PRDATA_reg[26] , 
        \COREAPBLSRAM_0.PRDATA_reg[25] , 
        \COREAPBLSRAM_0.PRDATA_reg[24] , 
        \COREAPBLSRAM_0.PRDATA_reg[23] , 
        \COREAPBLSRAM_0.PRDATA_reg[22] , 
        \COREAPBLSRAM_0.PRDATA_reg[21] , 
        \COREAPBLSRAM_0.PRDATA_reg[20] , 
        \COREAPBLSRAM_0.PRDATA_reg[19] , 
        \COREAPBLSRAM_0.PRDATA_reg[18] , 
        \COREAPBLSRAM_0.PRDATA_reg[17] , 
        \COREAPBLSRAM_0.PRDATA_reg[16] , 
        \COREAPBLSRAM_0.PRDATA_reg[15] , 
        \COREAPBLSRAM_0.PRDATA_reg[14] , 
        \COREAPBLSRAM_0.PRDATA_reg[13] , 
        \COREAPBLSRAM_0.PRDATA_reg[12] , 
        \COREAPBLSRAM_0.PRDATA_reg[11] , 
        \COREAPBLSRAM_0.PRDATA_reg[10] , 
        \COREAPBLSRAM_0.PRDATA_reg[9] , \COREAPBLSRAM_0.PRDATA_reg[8] , 
        \COREAPBLSRAM_0.PRDATA_reg[7] , \COREAPBLSRAM_0.PRDATA_reg[6] , 
        \COREAPBLSRAM_0.PRDATA_reg[5] , \COREAPBLSRAM_0.PRDATA_reg[4] , 
        \COREAPBLSRAM_0.PRDATA_reg[3] , \COREAPBLSRAM_0.PRDATA_reg[2] , 
        \COREAPBLSRAM_0.PRDATA_reg[1] , \COREAPBLSRAM_0.PRDATA_reg[0] })
        , .lsram_width32_PRDATA({
        \COREAPBLSRAM_0.lsram_width32_PRDATA[31] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[30] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[29] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[28] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[27] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[26] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[25] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[24] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[23] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[22] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[21] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[20] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[19] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[18] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[17] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[16] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[15] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[14] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[13] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[12] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[11] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[10] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[9] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[8] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[7] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[6] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[5] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[4] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[3] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[2] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[1] , 
        \COREAPBLSRAM_0.lsram_width32_PRDATA[0] }), 
        .hello_regs_MSS_0_FIC_0_APB_MASTER_PADDR({
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PADDR[27] , 
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PADDR[26] , 
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PADDR[25] , 
        \hello_regs_MSS_0_FIC_0_APB_MASTER_PADDR[24] }), 
        .CoreAPB3_0_APBmslave4_PADDR({\CoreAPB3_0_APBmslave4_PADDR[8] , 
        \CoreAPB3_0_APBmslave4_PADDR[7] , 
        \CoreAPB3_0_APBmslave4_PADDR[6] , 
        \CoreAPB3_0_APBmslave4_PADDR[5] , 
        \CoreAPB3_0_APBmslave4_PADDR[4] , 
        \CoreAPB3_0_APBmslave4_PADDR[3] , 
        \CoreAPB3_0_APBmslave4_PADDR[2] , 
        \CoreAPB3_0_APBmslave4_PADDR[1] , 
        \CoreAPB3_0_APBmslave4_PADDR[0] }), 
        .CoreAPB3_0_APBmslave4_PWDATA({
        \CoreAPB3_0_APBmslave4_PWDATA[31] , 
        \CoreAPB3_0_APBmslave4_PWDATA[30] , 
        \CoreAPB3_0_APBmslave4_PWDATA[29] , 
        \CoreAPB3_0_APBmslave4_PWDATA[28] , 
        \CoreAPB3_0_APBmslave4_PWDATA[27] , 
        \CoreAPB3_0_APBmslave4_PWDATA[26] , 
        \CoreAPB3_0_APBmslave4_PWDATA[25] , 
        \CoreAPB3_0_APBmslave4_PWDATA[24] , 
        \CoreAPB3_0_APBmslave4_PWDATA[23] , 
        \CoreAPB3_0_APBmslave4_PWDATA[22] , 
        \CoreAPB3_0_APBmslave4_PWDATA[21] , 
        \CoreAPB3_0_APBmslave4_PWDATA[20] , 
        \CoreAPB3_0_APBmslave4_PWDATA[19] , 
        \CoreAPB3_0_APBmslave4_PWDATA[18] , 
        \CoreAPB3_0_APBmslave4_PWDATA[17] , 
        \CoreAPB3_0_APBmslave4_PWDATA[16] , 
        \CoreAPB3_0_APBmslave4_PWDATA[15] , 
        \CoreAPB3_0_APBmslave4_PWDATA[14] , 
        \CoreAPB3_0_APBmslave4_PWDATA[13] , 
        \CoreAPB3_0_APBmslave4_PWDATA[12] , 
        \CoreAPB3_0_APBmslave4_PWDATA[11] , 
        \CoreAPB3_0_APBmslave4_PWDATA[10] , 
        \CoreAPB3_0_APBmslave4_PWDATA[9] , 
        \CoreAPB3_0_APBmslave4_PWDATA[8] , 
        \CoreAPB3_0_APBmslave4_PWDATA[7] , 
        \CoreAPB3_0_APBmslave4_PWDATA[6] , 
        \CoreAPB3_0_APBmslave4_PWDATA[5] , 
        \CoreAPB3_0_APBmslave4_PWDATA[4] , 
        \CoreAPB3_0_APBmslave4_PWDATA[3] , 
        \CoreAPB3_0_APBmslave4_PWDATA[2] , 
        \CoreAPB3_0_APBmslave4_PWDATA[1] , 
        \CoreAPB3_0_APBmslave4_PWDATA[0] }), .MSS_RESET_N_M2F_c(
        MSS_RESET_N_M2F_c), .FCCC_0_GL1(FCCC_0_GL1), .PRDATA4(
        \COREAPBLSRAM_0.PRDATA4 ), .CoreAPB3_0_APBmslave4_PREADY(
        CoreAPB3_0_APBmslave4_PREADY), .CoreAPB3_0_APBmslave4_PWRITE(
        CoreAPB3_0_APBmslave4_PWRITE), .CoreAPB3_0_APBmslave4_PENABLE(
        CoreAPB3_0_APBmslave4_PENABLE), .N_928(N_928), 
        .hello_regs_MSS_0_FIC_0_APB_MASTER_PSELx(
        hello_regs_MSS_0_FIC_0_APB_MASTER_PSELx));
    
endmodule
